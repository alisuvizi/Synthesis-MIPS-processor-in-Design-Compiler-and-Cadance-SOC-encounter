module instruction_mem (
	clk, 
	pc, 
	instruction);
   input clk;
   input [7:0] pc;
   output [15:0] instruction;

   assign instruction[0] = 1'b0 ;
   assign instruction[1] = 1'b0 ;
   assign instruction[2] = 1'b0 ;
   assign instruction[3] = 1'b0 ;
   assign instruction[4] = 1'b0 ;
   assign instruction[5] = 1'b0 ;
   assign instruction[6] = 1'b0 ;
   assign instruction[7] = 1'b0 ;
   assign instruction[8] = 1'b0 ;
   assign instruction[9] = 1'b0 ;
   assign instruction[10] = 1'b0 ;
   assign instruction[11] = 1'b0 ;
   assign instruction[12] = 1'b0 ;
   assign instruction[13] = 1'b0 ;
   assign instruction[14] = 1'b0 ;
   assign instruction[15] = 1'b0 ;
endmodule

module IF_stage_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   ADDFX2 U1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.CI(n1), 
	.B(B[1]), 
	.A(A[1]));
   ADDFX2 U1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(B[5]), 
	.A(A[5]));
   ADDFX2 U1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(B[4]), 
	.A(A[4]));
   ADDFX2 U1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(B[3]), 
	.A(A[3]));
   ADDFX2 U1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(B[2]), 
	.A(A[2]));
   ADDFX2 U1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(B[6]), 
	.A(A[6]));
   XOR3X2 U1_7 (.Y(SUM[7]), 
	.C(carry[7]), 
	.B(B[7]), 
	.A(A[7]));
   XOR2X1 U1 (.Y(SUM[0]), 
	.B(A[0]), 
	.A(B[0]));
   AND2X2 U2 (.Y(n1), 
	.B(A[0]), 
	.A(B[0]));
endmodule

module IF_stage (
	clk, 
	rst, 
	instruction_fetch_en, 
	branch_offset_imm, 
	branch_taken, 
	pc, 
	instruction);
   input clk;
   input rst;
   input instruction_fetch_en;
   input [5:0] branch_offset_imm;
   input branch_taken;
   output [7:0] pc;
   output [15:0] instruction;

   // Internal wires
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire \U3/U1/Z_0 ;
   wire \U3/U1/Z_1 ;
   wire \U3/U1/Z_2 ;
   wire \U3/U1/Z_3 ;
   wire \U3/U1/Z_4 ;
   wire \U3/U1/Z_7 ;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;

   assign instruction[15] = 1'b0 ;
   assign instruction[14] = 1'b0 ;
   assign instruction[13] = 1'b0 ;
   assign instruction[12] = 1'b0 ;
   assign instruction[11] = 1'b0 ;
   assign instruction[10] = 1'b0 ;
   assign instruction[9] = 1'b0 ;
   assign instruction[8] = 1'b0 ;
   assign instruction[7] = 1'b0 ;
   assign instruction[6] = 1'b0 ;
   assign instruction[5] = 1'b0 ;
   assign instruction[4] = 1'b0 ;
   assign instruction[3] = 1'b0 ;
   assign instruction[2] = 1'b0 ;
   assign instruction[1] = 1'b0 ;
   assign instruction[0] = 1'b0 ;

   instruction_mem imem (.clk(clk), 
	.pc({ pc[7],
		pc[6],
		pc[5],
		pc[4],
		pc[3],
		pc[2],
		pc[1],
		pc[0] }), 
	.instruction ());
   IF_stage_DW01_add_0 r56 (.A({ pc[7],
		pc[6],
		pc[5],
		pc[4],
		pc[3],
		pc[2],
		pc[1],
		pc[0] }), 
	.B({ \U3/U1/Z_7 ,
		\U3/U1/Z_7 ,
		\U3/U1/Z_7 ,
		\U3/U1/Z_4 ,
		\U3/U1/Z_3 ,
		\U3/U1/Z_2 ,
		\U3/U1/Z_1 ,
		\U3/U1/Z_0  }), 
	.CI(1'b0), 
	.SUM({ N29,
		N28,
		N27,
		N26,
		N25,
		N24,
		N23,
		N22 }));
   DFFRHQX1 \pc_reg[1]  (.RN(n19), 
	.Q(pc[1]), 
	.D(n17), 
	.CK(clk));
   DFFRHQX1 \pc_reg[2]  (.RN(n19), 
	.Q(pc[2]), 
	.D(n16), 
	.CK(clk));
   DFFRHQX1 \pc_reg[3]  (.RN(n19), 
	.Q(pc[3]), 
	.D(n15), 
	.CK(clk));
   DFFRHQX1 \pc_reg[4]  (.RN(n19), 
	.Q(pc[4]), 
	.D(n14), 
	.CK(clk));
   DFFRHQX1 \pc_reg[5]  (.RN(n19), 
	.Q(pc[5]), 
	.D(n13), 
	.CK(clk));
   DFFRHQX1 \pc_reg[6]  (.RN(n19), 
	.Q(pc[6]), 
	.D(n12), 
	.CK(clk));
   DFFRHQX1 \pc_reg[7]  (.RN(n19), 
	.Q(pc[7]), 
	.D(n11), 
	.CK(clk));
   DFFRHQX1 \pc_reg[0]  (.RN(n19), 
	.Q(pc[0]), 
	.D(n18), 
	.CK(clk));
   MX2X1 U4 (.Y(n11), 
	.S0(instruction_fetch_en), 
	.B(N29), 
	.A(pc[7]));
   MX2X1 U5 (.Y(n12), 
	.S0(instruction_fetch_en), 
	.B(N28), 
	.A(pc[6]));
   MX2X1 U6 (.Y(n13), 
	.S0(instruction_fetch_en), 
	.B(N27), 
	.A(pc[5]));
   MX2X1 U7 (.Y(n14), 
	.S0(instruction_fetch_en), 
	.B(N26), 
	.A(pc[4]));
   MX2X1 U8 (.Y(n15), 
	.S0(instruction_fetch_en), 
	.B(N25), 
	.A(pc[3]));
   MX2X1 U9 (.Y(n16), 
	.S0(instruction_fetch_en), 
	.B(N24), 
	.A(pc[2]));
   MX2X1 U10 (.Y(n17), 
	.S0(instruction_fetch_en), 
	.B(N23), 
	.A(pc[1]));
   MX2X1 U11 (.Y(n18), 
	.S0(instruction_fetch_en), 
	.B(N22), 
	.A(pc[0]));
   INVX1 U12 (.Y(n19), 
	.A(rst));
   AND2X1 U13 (.Y(\U3/U1/Z_7 ), 
	.B(branch_offset_imm[5]), 
	.A(branch_taken));
   AND2X1 U14 (.Y(\U3/U1/Z_4 ), 
	.B(branch_taken), 
	.A(branch_offset_imm[4]));
   AND2X1 U15 (.Y(\U3/U1/Z_3 ), 
	.B(branch_taken), 
	.A(branch_offset_imm[3]));
   AND2X1 U16 (.Y(\U3/U1/Z_2 ), 
	.B(branch_taken), 
	.A(branch_offset_imm[2]));
   AND2X1 U17 (.Y(\U3/U1/Z_1 ), 
	.B(branch_taken), 
	.A(branch_offset_imm[1]));
   NAND2BX1 U18 (.Y(\U3/U1/Z_0 ), 
	.B(branch_taken), 
	.AN(branch_offset_imm[0]));
endmodule

module ID_stage (
	clk, 
	rst, 
	instruction_decode_en, 
	pipeline_reg_out, 
	instruction, 
	branch_offset_imm, 
	branch_taken, 
	reg_read_addr_1, 
	reg_read_addr_2, 
	reg_read_data_1, 
	reg_read_data_2, 
	decoding_op_src1, 
	decoding_op_src2);
   input clk;
   input rst;
   input instruction_decode_en;
   output [56:0] pipeline_reg_out;
   input [15:0] instruction;
   output [5:0] branch_offset_imm;
   output branch_taken;
   output [2:0] reg_read_addr_1;
   output [2:0] reg_read_addr_2;
   input [15:0] reg_read_data_1;
   input [15:0] reg_read_data_2;
   output [2:0] decoding_op_src1;
   output [2:0] decoding_op_src2;

   // Internal wires
   wire write_back_en;
   wire n78;
   wire n80;
   wire n54;
   wire n55;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n79;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n135;
   wire n136;
   wire [15:9] instruction_reg;
   wire [2:0] ex_alu_cmd;
   wire [15:0] ex_alu_src2;

   assign decoding_op_src1[2] = reg_read_addr_1[2] ;
   assign decoding_op_src1[1] = reg_read_addr_1[1] ;
   assign decoding_op_src1[0] = reg_read_addr_1[0] ;

   DFFRHQXL \instruction_reg_reg[2]  (.RN(n136), 
	.Q(branch_offset_imm[2]), 
	.D(n125), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[1]  (.RN(n136), 
	.Q(branch_offset_imm[1]), 
	.D(n126), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[0]  (.RN(n136), 
	.Q(branch_offset_imm[0]), 
	.D(n127), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[11]  (.RN(n136), 
	.Q(instruction_reg[11]), 
	.D(n116), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[10]  (.RN(n136), 
	.Q(instruction_reg[10]), 
	.D(n117), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[9]  (.RN(n136), 
	.Q(instruction_reg[9]), 
	.D(n118), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[4]  (.RN(n136), 
	.Q(branch_offset_imm[4]), 
	.D(n123), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[3]  (.RN(n136), 
	.Q(branch_offset_imm[3]), 
	.D(n124), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[5]  (.RN(n136), 
	.Q(branch_offset_imm[5]), 
	.D(n122), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[3]  (.RN(n136), 
	.Q(pipeline_reg_out[3]), 
	.D(n130), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[2]  (.RN(n136), 
	.Q(pipeline_reg_out[2]), 
	.D(n129), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[1]  (.RN(n136), 
	.Q(pipeline_reg_out[1]), 
	.D(n131), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[56]  (.RN(n136), 
	.Q(pipeline_reg_out[56]), 
	.D(ex_alu_cmd[2]), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[15]  (.RN(n136), 
	.Q(instruction_reg[15]), 
	.D(n80), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[12]  (.RN(n136), 
	.Q(instruction_reg[12]), 
	.D(n54), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[13]  (.RN(n136), 
	.Q(instruction_reg[13]), 
	.D(n55), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[14]  (.RN(n136), 
	.Q(instruction_reg[14]), 
	.D(n78), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[55]  (.RN(n136), 
	.Q(pipeline_reg_out[55]), 
	.D(ex_alu_cmd[1]), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[7]  (.RN(n136), 
	.Q(reg_read_addr_1[1]), 
	.D(n120), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[6]  (.RN(n136), 
	.Q(reg_read_addr_1[0]), 
	.D(n121), 
	.CK(clk));
   DFFRHQXL \instruction_reg_reg[8]  (.RN(n136), 
	.Q(reg_read_addr_1[2]), 
	.D(n119), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[38]  (.RN(n136), 
	.Q(pipeline_reg_out[38]), 
	.D(reg_read_data_1[0]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[33]  (.RN(n136), 
	.Q(pipeline_reg_out[33]), 
	.D(ex_alu_src2[11]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[35]  (.RN(n136), 
	.Q(pipeline_reg_out[35]), 
	.D(ex_alu_src2[13]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[36]  (.RN(n136), 
	.Q(pipeline_reg_out[36]), 
	.D(ex_alu_src2[14]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[29]  (.RN(n136), 
	.Q(pipeline_reg_out[29]), 
	.D(ex_alu_src2[7]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[32]  (.RN(n136), 
	.Q(pipeline_reg_out[32]), 
	.D(ex_alu_src2[10]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[26]  (.RN(n136), 
	.Q(pipeline_reg_out[26]), 
	.D(n111), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[27]  (.RN(n136), 
	.Q(pipeline_reg_out[27]), 
	.D(ex_alu_src2[5]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[52]  (.RN(n136), 
	.Q(pipeline_reg_out[52]), 
	.D(reg_read_data_1[14]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[28]  (.RN(n136), 
	.Q(pipeline_reg_out[28]), 
	.D(ex_alu_src2[6]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[34]  (.RN(n136), 
	.Q(pipeline_reg_out[34]), 
	.D(ex_alu_src2[12]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[51]  (.RN(n136), 
	.Q(pipeline_reg_out[51]), 
	.D(reg_read_data_1[13]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[39]  (.RN(n136), 
	.Q(pipeline_reg_out[39]), 
	.D(reg_read_data_1[1]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[53]  (.RN(n136), 
	.Q(pipeline_reg_out[53]), 
	.D(reg_read_data_1[15]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[30]  (.RN(n136), 
	.Q(pipeline_reg_out[30]), 
	.D(ex_alu_src2[8]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[31]  (.RN(n136), 
	.Q(pipeline_reg_out[31]), 
	.D(ex_alu_src2[9]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[25]  (.RN(n136), 
	.Q(pipeline_reg_out[25]), 
	.D(n112), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[41]  (.RN(n136), 
	.Q(pipeline_reg_out[41]), 
	.D(reg_read_data_1[3]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[42]  (.RN(n136), 
	.Q(pipeline_reg_out[42]), 
	.D(reg_read_data_1[4]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[50]  (.RN(n136), 
	.Q(pipeline_reg_out[50]), 
	.D(reg_read_data_1[12]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[45]  (.RN(n136), 
	.Q(pipeline_reg_out[45]), 
	.D(reg_read_data_1[7]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[49]  (.RN(n136), 
	.Q(pipeline_reg_out[49]), 
	.D(reg_read_data_1[11]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[48]  (.RN(n136), 
	.Q(pipeline_reg_out[48]), 
	.D(reg_read_data_1[10]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[46]  (.RN(n136), 
	.Q(pipeline_reg_out[46]), 
	.D(reg_read_data_1[8]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[47]  (.RN(n136), 
	.Q(pipeline_reg_out[47]), 
	.D(reg_read_data_1[9]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[44]  (.RN(n136), 
	.Q(pipeline_reg_out[44]), 
	.D(reg_read_data_1[6]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[40]  (.RN(n136), 
	.Q(pipeline_reg_out[40]), 
	.D(reg_read_data_1[2]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[37]  (.RN(n136), 
	.Q(pipeline_reg_out[37]), 
	.D(ex_alu_src2[15]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[43]  (.RN(n136), 
	.Q(pipeline_reg_out[43]), 
	.D(reg_read_data_1[5]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[22]  (.RN(n136), 
	.Q(pipeline_reg_out[22]), 
	.D(n115), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[24]  (.RN(n136), 
	.Q(pipeline_reg_out[24]), 
	.D(n113), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[23]  (.RN(n136), 
	.Q(pipeline_reg_out[23]), 
	.D(n114), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[21]  (.RN(n136), 
	.Q(pipeline_reg_out[21]), 
	.D(n135), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[20]  (.RN(n136), 
	.Q(pipeline_reg_out[20]), 
	.D(reg_read_data_2[15]), 
	.CK(clk));
   DFFRHQXL \pipeline_reg_out_reg[19]  (.RN(n136), 
	.Q(pipeline_reg_out[19]), 
	.D(reg_read_data_2[14]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[18]  (.RN(n136), 
	.Q(pipeline_reg_out[18]), 
	.D(reg_read_data_2[13]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[17]  (.RN(n136), 
	.Q(pipeline_reg_out[17]), 
	.D(reg_read_data_2[12]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[16]  (.RN(n136), 
	.Q(pipeline_reg_out[16]), 
	.D(reg_read_data_2[11]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[15]  (.RN(n136), 
	.Q(pipeline_reg_out[15]), 
	.D(reg_read_data_2[10]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[14]  (.RN(n136), 
	.Q(pipeline_reg_out[14]), 
	.D(reg_read_data_2[9]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[13]  (.RN(n136), 
	.Q(pipeline_reg_out[13]), 
	.D(reg_read_data_2[8]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[12]  (.RN(n136), 
	.Q(pipeline_reg_out[12]), 
	.D(reg_read_data_2[7]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[11]  (.RN(n136), 
	.Q(pipeline_reg_out[11]), 
	.D(reg_read_data_2[6]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[10]  (.RN(n136), 
	.Q(pipeline_reg_out[10]), 
	.D(reg_read_data_2[5]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[9]  (.RN(n136), 
	.Q(pipeline_reg_out[9]), 
	.D(reg_read_data_2[4]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[8]  (.RN(n136), 
	.Q(pipeline_reg_out[8]), 
	.D(reg_read_data_2[3]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[7]  (.RN(n136), 
	.Q(pipeline_reg_out[7]), 
	.D(reg_read_data_2[2]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[6]  (.RN(n136), 
	.Q(pipeline_reg_out[6]), 
	.D(reg_read_data_2[1]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[5]  (.RN(n136), 
	.Q(pipeline_reg_out[5]), 
	.D(reg_read_data_2[0]), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[4]  (.RN(n136), 
	.Q(pipeline_reg_out[4]), 
	.D(write_back_en), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[0]  (.RN(n136), 
	.Q(pipeline_reg_out[0]), 
	.D(n128), 
	.CK(clk));
   DFFRHQX1 \pipeline_reg_out_reg[54]  (.RN(n136), 
	.Q(pipeline_reg_out[54]), 
	.D(ex_alu_cmd[0]), 
	.CK(clk));
   NOR4X1 U3 (.Y(write_back_en), 
	.D(n69), 
	.C(n68), 
	.B(n67), 
	.A(rst));
   AND3X1 U4 (.Y(n69), 
	.C(n72), 
	.B(n71), 
	.A(n70));
   MX2X1 U5 (.Y(n111), 
	.S0(n73), 
	.B(reg_read_data_2[4]), 
	.A(branch_offset_imm[4]));
   MX2X1 U6 (.Y(n112), 
	.S0(n73), 
	.B(reg_read_data_2[3]), 
	.A(branch_offset_imm[3]));
   MX2X1 U7 (.Y(n113), 
	.S0(n73), 
	.B(reg_read_data_2[2]), 
	.A(branch_offset_imm[2]));
   MX2X1 U8 (.Y(n114), 
	.S0(n73), 
	.B(reg_read_data_2[1]), 
	.A(branch_offset_imm[1]));
   MX2X1 U9 (.Y(n115), 
	.S0(n73), 
	.B(reg_read_data_2[0]), 
	.A(branch_offset_imm[0]));
   MX2X1 U10 (.Y(n116), 
	.S0(instruction_decode_en), 
	.B(instruction[11]), 
	.A(instruction_reg[11]));
   MX2X1 U11 (.Y(n117), 
	.S0(instruction_decode_en), 
	.B(instruction[10]), 
	.A(instruction_reg[10]));
   MX2X1 U12 (.Y(n118), 
	.S0(instruction_decode_en), 
	.B(instruction[9]), 
	.A(instruction_reg[9]));
   MX2X1 U13 (.Y(n119), 
	.S0(instruction_decode_en), 
	.B(instruction[8]), 
	.A(reg_read_addr_1[2]));
   MX2X1 U14 (.Y(n120), 
	.S0(instruction_decode_en), 
	.B(instruction[7]), 
	.A(reg_read_addr_1[1]));
   MX2X1 U15 (.Y(n121), 
	.S0(instruction_decode_en), 
	.B(instruction[6]), 
	.A(reg_read_addr_1[0]));
   MX2X1 U16 (.Y(n122), 
	.S0(instruction_decode_en), 
	.B(instruction[5]), 
	.A(branch_offset_imm[5]));
   MX2X1 U17 (.Y(n123), 
	.S0(instruction_decode_en), 
	.B(instruction[4]), 
	.A(branch_offset_imm[4]));
   MX2X1 U18 (.Y(n124), 
	.S0(instruction_decode_en), 
	.B(instruction[3]), 
	.A(branch_offset_imm[3]));
   MX2X1 U19 (.Y(n125), 
	.S0(instruction_decode_en), 
	.B(instruction[2]), 
	.A(branch_offset_imm[2]));
   MX2X1 U20 (.Y(n126), 
	.S0(instruction_decode_en), 
	.B(instruction[1]), 
	.A(branch_offset_imm[1]));
   MX2X1 U21 (.Y(n127), 
	.S0(instruction_decode_en), 
	.B(instruction[0]), 
	.A(branch_offset_imm[0]));
   INVX1 U22 (.Y(n128), 
	.A(n74));
   INVX1 U23 (.Y(reg_read_addr_2[2]), 
	.A(n75));
   INVX1 U24 (.Y(reg_read_addr_2[1]), 
	.A(n76));
   INVX1 U25 (.Y(reg_read_addr_2[0]), 
	.A(n77));
   MX2X1 U26 (.Y(n80), 
	.S0(instruction_decode_en), 
	.B(instruction[15]), 
	.A(instruction_reg[15]));
   MX2X1 U27 (.Y(n78), 
	.S0(instruction_decode_en), 
	.B(instruction[14]), 
	.A(instruction_reg[14]));
   MX2X1 U28 (.Y(n55), 
	.S0(instruction_decode_en), 
	.B(instruction[13]), 
	.A(instruction_reg[13]));
   MX2X1 U29 (.Y(n54), 
	.S0(instruction_decode_en), 
	.B(instruction[12]), 
	.A(instruction_reg[12]));
   OAI2BB1X1 U30 (.Y(ex_alu_src2[9]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[9]));
   OAI2BB1X1 U31 (.Y(ex_alu_src2[8]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[8]));
   OAI2BB1X1 U32 (.Y(ex_alu_src2[7]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[7]));
   OAI2BB1X1 U33 (.Y(ex_alu_src2[6]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[6]));
   OAI2BB1X1 U34 (.Y(ex_alu_src2[5]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[5]));
   OAI2BB1X1 U35 (.Y(ex_alu_src2[15]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[15]));
   OAI2BB1X1 U36 (.Y(ex_alu_src2[14]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[14]));
   OAI2BB1X1 U37 (.Y(ex_alu_src2[13]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[13]));
   OAI2BB1X1 U38 (.Y(ex_alu_src2[12]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[12]));
   OAI2BB1X1 U39 (.Y(ex_alu_src2[11]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[11]));
   OAI2BB1X1 U40 (.Y(ex_alu_src2[10]), 
	.B0(n79), 
	.A1N(n73), 
	.A0N(reg_read_data_2[10]));
   NAND2X1 U41 (.Y(n79), 
	.B(n81), 
	.A(branch_offset_imm[5]));
   INVX1 U42 (.Y(n73), 
	.A(n81));
   OAI21XL U43 (.Y(n81), 
	.B0(n74), 
	.A1(n82), 
	.A0(rst));
   NAND3X1 U44 (.Y(n74), 
	.C(n84), 
	.B(n136), 
	.A(n83));
   AOI211X1 U45 (.Y(n82), 
	.C0(n85), 
	.B0(n68), 
	.A1(n70), 
	.A0(n67));
   AND3X1 U46 (.Y(n85), 
	.C(n88), 
	.B(n87), 
	.A(n86));
   NOR2BX1 U47 (.Y(n68), 
	.B(n83), 
	.AN(n84));
   NOR3X1 U48 (.Y(n84), 
	.C(n90), 
	.B(n89), 
	.A(n71));
   NOR2X1 U49 (.Y(n67), 
	.B(n72), 
	.A(n71));
   OAI31X1 U50 (.Y(ex_alu_cmd[2]), 
	.B0(n92), 
	.A2(n72), 
	.A1(n70), 
	.A0(n91));
   OAI21XL U51 (.Y(ex_alu_cmd[1]), 
	.B0(n92), 
	.A1(n91), 
	.A0(n93));
   AOI22X1 U52 (.Y(n93), 
	.B1(n94), 
	.B0(n88), 
	.A1(n89), 
	.A0(n70));
   OAI31X1 U53 (.Y(ex_alu_cmd[0]), 
	.B0(n92), 
	.A2(n86), 
	.A1(n88), 
	.A0(n91));
   NAND4X1 U54 (.Y(n92), 
	.D(n136), 
	.C(n72), 
	.B(n87), 
	.A(n70));
   INVX1 U55 (.Y(n87), 
	.A(n71));
   NOR2X1 U56 (.Y(n70), 
	.B(n88), 
	.A(n94));
   NOR2X1 U57 (.Y(n86), 
	.B(n89), 
	.A(n94));
   INVX1 U58 (.Y(n89), 
	.A(n72));
   NAND2X1 U59 (.Y(n72), 
	.B(instruction_decode_en), 
	.A(instruction_reg[14]));
   INVX1 U60 (.Y(n94), 
	.A(n90));
   NAND2X1 U61 (.Y(n90), 
	.B(instruction_decode_en), 
	.A(instruction_reg[13]));
   INVX1 U62 (.Y(n88), 
	.A(n83));
   NAND2X1 U63 (.Y(n83), 
	.B(instruction_decode_en), 
	.A(instruction_reg[12]));
   NAND2X1 U64 (.Y(n91), 
	.B(n136), 
	.A(n71));
   INVX1 U65 (.Y(n136), 
	.A(rst));
   NAND2X1 U66 (.Y(n71), 
	.B(instruction_decode_en), 
	.A(instruction_reg[15]));
   NOR2X1 U67 (.Y(decoding_op_src2[2]), 
	.B(n95), 
	.A(n75));
   MXI2X1 U68 (.Y(n75), 
	.S0(n135), 
	.B(instruction_reg[11]), 
	.A(branch_offset_imm[5]));
   NOR2X1 U69 (.Y(decoding_op_src2[1]), 
	.B(n95), 
	.A(n76));
   MXI2X1 U70 (.Y(n76), 
	.S0(n135), 
	.B(instruction_reg[10]), 
	.A(branch_offset_imm[4]));
   NOR2X1 U71 (.Y(decoding_op_src2[0]), 
	.B(n95), 
	.A(n77));
   MX2X1 U72 (.Y(n95), 
	.S0(instruction_reg[15]), 
	.B(n97), 
	.A(n96));
   MXI2X1 U73 (.Y(n97), 
	.S0(n100), 
	.B(n99), 
	.A(n98));
   XNOR2X1 U74 (.Y(n99), 
	.B(instruction_reg[13]), 
	.A(instruction_reg[12]));
   NOR2X1 U75 (.Y(n96), 
	.B(n98), 
	.A(instruction_reg[14]));
   INVX1 U76 (.Y(n98), 
	.A(n101));
   MXI2X1 U77 (.Y(n77), 
	.S0(n135), 
	.B(instruction_reg[9]), 
	.A(branch_offset_imm[3]));
   AND4X1 U78 (.Y(n135), 
	.D(instruction_reg[15]), 
	.C(instruction_reg[12]), 
	.B(instruction_reg[13]), 
	.A(n100));
   INVX1 U79 (.Y(n100), 
	.A(instruction_reg[14]));
   NOR2X1 U80 (.Y(branch_taken), 
	.B(n103), 
	.A(n102));
   NAND4X1 U81 (.Y(n103), 
	.D(n105), 
	.C(n104), 
	.B(instruction_reg[14]), 
	.A(n101));
   NOR4BX1 U82 (.Y(n105), 
	.D(reg_read_data_1[0]), 
	.C(n129), 
	.B(reg_read_data_1[10]), 
	.AN(n106));
   AND2X1 U83 (.Y(n129), 
	.B(instruction_decode_en), 
	.A(instruction_reg[10]));
   NOR3X1 U84 (.Y(n106), 
	.C(reg_read_data_1[12]), 
	.B(reg_read_data_1[13]), 
	.A(reg_read_data_1[11]));
   NOR3BX1 U85 (.Y(n104), 
	.C(n131), 
	.B(n130), 
	.AN(instruction_reg[15]));
   AND2X1 U86 (.Y(n131), 
	.B(instruction_decode_en), 
	.A(instruction_reg[9]));
   AND2X1 U87 (.Y(n130), 
	.B(instruction_decode_en), 
	.A(instruction_reg[11]));
   NOR2X1 U88 (.Y(n101), 
	.B(instruction_reg[13]), 
	.A(instruction_reg[12]));
   NAND4X1 U89 (.Y(n102), 
	.D(n110), 
	.C(n109), 
	.B(n108), 
	.A(n107));
   NOR3X1 U90 (.Y(n110), 
	.C(reg_read_data_1[8]), 
	.B(reg_read_data_1[9]), 
	.A(reg_read_data_1[7]));
   NOR3X1 U91 (.Y(n109), 
	.C(reg_read_data_1[5]), 
	.B(reg_read_data_1[6]), 
	.A(reg_read_data_1[4]));
   NOR3X1 U92 (.Y(n108), 
	.C(reg_read_data_1[2]), 
	.B(reg_read_data_1[3]), 
	.A(reg_read_data_1[1]));
   NOR2X1 U93 (.Y(n107), 
	.B(reg_read_data_1[14]), 
	.A(reg_read_data_1[15]));
endmodule

module alu_DW01_addsub_0 (
	A, 
	B, 
	CI, 
	ADD_SUB, 
	SUM, 
	CO);
   input [15:0] A;
   input [15:0] B;
   input CI;
   input ADD_SUB;
   output [15:0] SUM;
   output CO;

   // Internal wires
   wire [16:0] carry;
   wire [15:0] B_AS;

   assign carry[0] = ADD_SUB ;

   ADDFX2 U1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(B_AS[5]), 
	.A(A[5]));
   ADDFX2 U1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.CI(carry[8]), 
	.B(B_AS[8]), 
	.A(A[8]));
   ADDFX2 U1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(B_AS[7]), 
	.A(A[7]));
   ADDFX2 U1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(B_AS[4]), 
	.A(A[4]));
   ADDFX2 U1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(B_AS[6]), 
	.A(A[6]));
   ADDFX2 U1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(B_AS[3]), 
	.A(A[3]));
   ADDFX2 U1_13 (.S(SUM[13]), 
	.CO(carry[14]), 
	.CI(carry[13]), 
	.B(B_AS[13]), 
	.A(A[13]));
   ADDFX2 U1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(B_AS[2]), 
	.A(A[2]));
   ADDFX2 U1_12 (.S(SUM[12]), 
	.CO(carry[13]), 
	.CI(carry[12]), 
	.B(B_AS[12]), 
	.A(A[12]));
   ADDFX2 U1_11 (.S(SUM[11]), 
	.CO(carry[12]), 
	.CI(carry[11]), 
	.B(B_AS[11]), 
	.A(A[11]));
   ADDFX2 U1_10 (.S(SUM[10]), 
	.CO(carry[11]), 
	.CI(carry[10]), 
	.B(B_AS[10]), 
	.A(A[10]));
   ADDFX2 U1_9 (.S(SUM[9]), 
	.CO(carry[10]), 
	.CI(carry[9]), 
	.B(B_AS[9]), 
	.A(A[9]));
   ADDFX2 U1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(B_AS[1]), 
	.A(A[1]));
   ADDFX2 U1_0 (.S(SUM[0]), 
	.CO(carry[1]), 
	.CI(carry[0]), 
	.B(B_AS[0]), 
	.A(A[0]));
   ADDFX2 U1_14 (.S(SUM[14]), 
	.CO(carry[15]), 
	.CI(carry[14]), 
	.B(B_AS[14]), 
	.A(A[14]));
   XOR3X2 U1_15 (.Y(SUM[15]), 
	.C(carry[15]), 
	.B(B_AS[15]), 
	.A(A[15]));
   XOR2X1 U1 (.Y(B_AS[15]), 
	.B(carry[0]), 
	.A(B[15]));
   XOR2X1 U2 (.Y(B_AS[14]), 
	.B(carry[0]), 
	.A(B[14]));
   XOR2X1 U3 (.Y(B_AS[0]), 
	.B(carry[0]), 
	.A(B[0]));
   XOR2X1 U4 (.Y(B_AS[1]), 
	.B(carry[0]), 
	.A(B[1]));
   XOR2X1 U5 (.Y(B_AS[9]), 
	.B(carry[0]), 
	.A(B[9]));
   XOR2X1 U6 (.Y(B_AS[10]), 
	.B(carry[0]), 
	.A(B[10]));
   XOR2X1 U7 (.Y(B_AS[11]), 
	.B(carry[0]), 
	.A(B[11]));
   XOR2X1 U8 (.Y(B_AS[12]), 
	.B(carry[0]), 
	.A(B[12]));
   XOR2X1 U9 (.Y(B_AS[2]), 
	.B(carry[0]), 
	.A(B[2]));
   XOR2X1 U10 (.Y(B_AS[13]), 
	.B(carry[0]), 
	.A(B[13]));
   XOR2X1 U11 (.Y(B_AS[3]), 
	.B(carry[0]), 
	.A(B[3]));
   XOR2X1 U12 (.Y(B_AS[6]), 
	.B(carry[0]), 
	.A(B[6]));
   XOR2X1 U13 (.Y(B_AS[4]), 
	.B(carry[0]), 
	.A(B[4]));
   XOR2X1 U14 (.Y(B_AS[7]), 
	.B(carry[0]), 
	.A(B[7]));
   XOR2X1 U15 (.Y(B_AS[8]), 
	.B(carry[0]), 
	.A(B[8]));
   XOR2X1 U16 (.Y(B_AS[5]), 
	.B(carry[0]), 
	.A(B[5]));
endmodule

module alu_DW_rash_0 (
	A, 
	DATA_TC, 
	SH, 
	SH_TC, 
	B);
   input [15:0] A;
   input DATA_TC;
   input [15:0] SH;
   input SH_TC;
   output [15:0] B;

   // Internal wires
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;

   OAI222XL U3 (.Y(B[4]), 
	.C1(n71), 
	.C0(n36), 
	.B1(n30), 
	.B0(n27), 
	.A1(n25), 
	.A0(n26));
   OAI221XL U4 (.Y(B[2]), 
	.C0(n46), 
	.B1(n30), 
	.B0(n32), 
	.A1(n45), 
	.A0(n33));
   AOI2BB2X1 U5 (.Y(n46), 
	.B1(n48), 
	.B0(n47), 
	.A1N(n34), 
	.A0N(n25));
   OAI221XL U6 (.Y(n48), 
	.C0(n51), 
	.B1(n89), 
	.B0(n44), 
	.A1(n87), 
	.A0(n50));
   NOR2X1 U7 (.Y(B[11]), 
	.B(n57), 
	.A(n37));
   NOR2X1 U8 (.Y(B[12]), 
	.B(n71), 
	.A(n27));
   NOR2X1 U9 (.Y(B[13]), 
	.B(n71), 
	.A(n24));
   NOR2X1 U10 (.Y(B[14]), 
	.B(n71), 
	.A(n33));
   OAI22X1 U11 (.Y(B[8]), 
	.B1(n25), 
	.B0(n27), 
	.A1(n71), 
	.A0(n26));
   OAI221XL U12 (.Y(B[0]), 
	.C0(n60), 
	.B1(n30), 
	.B0(n26), 
	.A1(n45), 
	.A0(n27));
   AOI2BB2X1 U13 (.Y(n60), 
	.B1(n61), 
	.B0(n47), 
	.A1N(n36), 
	.A0N(n25));
   OR2X2 U14 (.Y(n25), 
	.B(n86), 
	.A(n57));
   OAI22X1 U15 (.Y(B[10]), 
	.B1(n25), 
	.B0(n33), 
	.A1(n71), 
	.A0(n32));
   OAI22X1 U16 (.Y(B[9]), 
	.B1(n25), 
	.B0(n24), 
	.A1(n71), 
	.A0(n23));
   INVX1 U17 (.Y(n71), 
	.A(n47));
   NAND2X1 U18 (.Y(n30), 
	.B(n86), 
	.A(n72));
   NOR2X1 U19 (.Y(B[15]), 
	.B(n29), 
	.A(n71));
   MX2X1 U20 (.Y(n37), 
	.S0(n86), 
	.B(n28), 
	.A(n29));
   INVX1 U21 (.Y(n84), 
	.A(n50));
   INVX1 U22 (.Y(n73), 
	.A(n44));
   INVX1 U23 (.Y(n72), 
	.A(n38));
   OAI222XL U24 (.Y(B[5]), 
	.C1(n71), 
	.C0(n35), 
	.B1(n30), 
	.B0(n24), 
	.A1(n25), 
	.A0(n23));
   OAI222XL U25 (.Y(B[6]), 
	.C1(n71), 
	.C0(n34), 
	.B1(n30), 
	.B0(n33), 
	.A1(n25), 
	.A0(n32));
   OAI222XL U26 (.Y(B[7]), 
	.C1(n71), 
	.C0(n31), 
	.B1(n30), 
	.B0(n29), 
	.A1(n25), 
	.A0(n28));
   NOR2X1 U27 (.Y(n42), 
	.B(SH[1]), 
	.A(SH[0]));
   NOR2X1 U28 (.Y(n41), 
	.B(SH[1]), 
	.A(n83));
   OAI222XL U29 (.Y(B[3]), 
	.C1(n25), 
	.C0(n31), 
	.B1(n71), 
	.B0(n39), 
	.A1(n38), 
	.A0(n37));
   AOI221X1 U30 (.Y(n39), 
	.C0(n43), 
	.B1(n42), 
	.B0(A[3]), 
	.A1(n41), 
	.A0(A[4]));
   OAI2BB2X1 U31 (.Y(n43), 
	.B1(n87), 
	.B0(n44), 
	.A1N(A[6]), 
	.A0N(n84));
   NOR2X1 U32 (.Y(n47), 
	.B(SH[2]), 
	.A(n57));
   AOI22X1 U33 (.Y(n33), 
	.B1(n41), 
	.B0(A[15]), 
	.A1(n42), 
	.A0(A[14]));
   NAND3BX1 U34 (.Y(n57), 
	.C(n64), 
	.B(n85), 
	.AN(SH[3]));
   AOI22X1 U35 (.Y(n51), 
	.B1(n42), 
	.B0(A[2]), 
	.A1(n41), 
	.A0(A[3]));
   NAND2X1 U36 (.Y(n44), 
	.B(SH[1]), 
	.A(n83));
   NAND2X1 U37 (.Y(n29), 
	.B(A[15]), 
	.A(n42));
   NAND3X1 U38 (.Y(n38), 
	.C(n64), 
	.B(n85), 
	.A(SH[3]));
   NOR3X1 U39 (.Y(n69), 
	.C(SH[8]), 
	.B(SH[9]), 
	.A(SH[7]));
   NAND2X1 U40 (.Y(n50), 
	.B(SH[1]), 
	.A(SH[0]));
   AOI221X1 U41 (.Y(n27), 
	.C0(n82), 
	.B1(A[14]), 
	.B0(n73), 
	.A1(n84), 
	.A0(A[15]));
   INVX1 U42 (.Y(n82), 
	.A(n70));
   AOI22X1 U43 (.Y(n70), 
	.B1(n42), 
	.B0(A[12]), 
	.A1(n41), 
	.A0(A[13]));
   AOI222X1 U44 (.Y(n24), 
	.C1(A[13]), 
	.C0(n42), 
	.B1(A[15]), 
	.B0(n73), 
	.A1(A[14]), 
	.A0(n41));
   AND4X2 U45 (.Y(n64), 
	.D(n69), 
	.C(n68), 
	.B(n67), 
	.A(n66));
   NOR2X1 U46 (.Y(n66), 
	.B(SH[10]), 
	.A(SH[11]));
   NOR3X1 U47 (.Y(n67), 
	.C(SH[13]), 
	.B(SH[14]), 
	.A(SH[12]));
   NOR3X1 U48 (.Y(n68), 
	.C(SH[5]), 
	.B(SH[6]), 
	.A(SH[4]));
   INVX1 U49 (.Y(n86), 
	.A(SH[2]));
   INVX1 U50 (.Y(n83), 
	.A(SH[0]));
   INVX1 U51 (.Y(n85), 
	.A(SH[15]));
   NAND2X1 U52 (.Y(n45), 
	.B(SH[2]), 
	.A(n72));
   AOI221X1 U53 (.Y(n26), 
	.C0(n81), 
	.B1(A[10]), 
	.B0(n73), 
	.A1(A[11]), 
	.A0(n84));
   INVX1 U54 (.Y(n81), 
	.A(n65));
   AOI22X1 U55 (.Y(n65), 
	.B1(n42), 
	.B0(A[8]), 
	.A1(n41), 
	.A0(A[9]));
   AOI221X1 U56 (.Y(n32), 
	.C0(n79), 
	.B1(A[12]), 
	.B0(n73), 
	.A1(n84), 
	.A0(A[13]));
   INVX1 U57 (.Y(n79), 
	.A(n59));
   AOI22X1 U58 (.Y(n59), 
	.B1(n42), 
	.B0(A[10]), 
	.A1(n41), 
	.A0(A[11]));
   AOI221X1 U59 (.Y(n23), 
	.C0(n77), 
	.B1(A[11]), 
	.B0(n73), 
	.A1(A[12]), 
	.A0(n84));
   INVX1 U60 (.Y(n77), 
	.A(n56));
   AOI22X1 U61 (.Y(n56), 
	.B1(n42), 
	.B0(A[9]), 
	.A1(n41), 
	.A0(A[10]));
   INVX1 U62 (.Y(n87), 
	.A(A[5]));
   OAI221XL U63 (.Y(n61), 
	.C0(n63), 
	.B1(n88), 
	.B0(n44), 
	.A1(n90), 
	.A0(n50));
   INVX1 U64 (.Y(n88), 
	.A(A[2]));
   AOI22X1 U65 (.Y(n63), 
	.B1(n42), 
	.B0(A[0]), 
	.A1(n41), 
	.A0(A[1]));
   INVX1 U66 (.Y(n89), 
	.A(A[4]));
   INVX1 U67 (.Y(n90), 
	.A(A[3]));
   AOI221X1 U68 (.Y(n35), 
	.C0(n76), 
	.B1(A[7]), 
	.B0(n73), 
	.A1(A[8]), 
	.A0(n84));
   INVX1 U69 (.Y(n76), 
	.A(n54));
   AOI22X1 U70 (.Y(n54), 
	.B1(n42), 
	.B0(A[5]), 
	.A1(n41), 
	.A0(A[6]));
   AOI221X1 U71 (.Y(n36), 
	.C0(n80), 
	.B1(A[6]), 
	.B0(n73), 
	.A1(A[7]), 
	.A0(n84));
   INVX1 U72 (.Y(n80), 
	.A(n62));
   AOI22X1 U73 (.Y(n62), 
	.B1(n42), 
	.B0(A[4]), 
	.A1(n41), 
	.A0(A[5]));
   AOI221X1 U74 (.Y(n34), 
	.C0(n75), 
	.B1(A[8]), 
	.B0(n73), 
	.A1(A[9]), 
	.A0(n84));
   INVX1 U75 (.Y(n75), 
	.A(n49));
   AOI22X1 U76 (.Y(n49), 
	.B1(n42), 
	.B0(A[6]), 
	.A1(n41), 
	.A0(A[7]));
   AOI221X1 U77 (.Y(n28), 
	.C0(n78), 
	.B1(A[13]), 
	.B0(n73), 
	.A1(n84), 
	.A0(A[14]));
   INVX1 U78 (.Y(n78), 
	.A(n58));
   AOI22X1 U79 (.Y(n58), 
	.B1(n42), 
	.B0(A[11]), 
	.A1(n41), 
	.A0(A[12]));
   AOI221X1 U80 (.Y(n31), 
	.C0(n74), 
	.B1(A[9]), 
	.B0(n73), 
	.A1(A[10]), 
	.A0(n84));
   INVX1 U81 (.Y(n74), 
	.A(n40));
   AOI22X1 U82 (.Y(n40), 
	.B1(n42), 
	.B0(A[7]), 
	.A1(n41), 
	.A0(A[8]));
   OAI221XL U83 (.Y(B[1]), 
	.C0(n52), 
	.B1(n30), 
	.B0(n23), 
	.A1(n45), 
	.A0(n24));
   AOI2BB2X1 U84 (.Y(n52), 
	.B1(n53), 
	.B0(n47), 
	.A1N(n35), 
	.A0N(n25));
   OAI221XL U85 (.Y(n53), 
	.C0(n55), 
	.B1(n90), 
	.B0(n44), 
	.A1(n89), 
	.A0(n50));
   AOI22X1 U86 (.Y(n55), 
	.B1(n42), 
	.B0(A[1]), 
	.A1(n41), 
	.A0(A[2]));
endmodule

module alu_DW01_ash_0 (
	A, 
	DATA_TC, 
	SH, 
	SH_TC, 
	B);
   input [15:0] A;
   input DATA_TC;
   input [15:0] SH;
   input SH_TC;
   output [15:0] B;

   // Internal wires
   wire \ML_int[1][15] ;
   wire \ML_int[1][14] ;
   wire \ML_int[1][13] ;
   wire \ML_int[1][12] ;
   wire \ML_int[1][11] ;
   wire \ML_int[1][10] ;
   wire \ML_int[1][9] ;
   wire \ML_int[1][8] ;
   wire \ML_int[1][7] ;
   wire \ML_int[1][6] ;
   wire \ML_int[1][5] ;
   wire \ML_int[1][4] ;
   wire \ML_int[1][3] ;
   wire \ML_int[1][2] ;
   wire \ML_int[1][1] ;
   wire \ML_int[1][0] ;
   wire \ML_int[2][15] ;
   wire \ML_int[2][14] ;
   wire \ML_int[2][13] ;
   wire \ML_int[2][12] ;
   wire \ML_int[2][11] ;
   wire \ML_int[2][10] ;
   wire \ML_int[2][9] ;
   wire \ML_int[2][8] ;
   wire \ML_int[2][7] ;
   wire \ML_int[2][6] ;
   wire \ML_int[2][5] ;
   wire \ML_int[2][4] ;
   wire \ML_int[2][3] ;
   wire \ML_int[2][2] ;
   wire \ML_int[2][1] ;
   wire \ML_int[2][0] ;
   wire \ML_int[3][15] ;
   wire \ML_int[3][14] ;
   wire \ML_int[3][13] ;
   wire \ML_int[3][12] ;
   wire \ML_int[3][8] ;
   wire \ML_int[3][7] ;
   wire \ML_int[3][6] ;
   wire \ML_int[3][5] ;
   wire \ML_int[3][4] ;
   wire \ML_int[4][15] ;
   wire \ML_int[4][14] ;
   wire \ML_int[4][13] ;
   wire \ML_int[4][12] ;
   wire \ML_int[4][11] ;
   wire \ML_int[4][10] ;
   wire \ML_int[4][9] ;
   wire \ML_int[4][8] ;
   wire \ML_int[6][15] ;
   wire \ML_int[6][14] ;
   wire \ML_int[6][13] ;
   wire \ML_int[6][12] ;
   wire \ML_int[6][11] ;
   wire \ML_int[6][10] ;
   wire \ML_int[6][9] ;
   wire \ML_int[6][8] ;
   wire \ML_int[6][7] ;
   wire \ML_int[6][6] ;
   wire \ML_int[6][5] ;
   wire \ML_int[6][4] ;
   wire \ML_int[6][3] ;
   wire \ML_int[6][2] ;
   wire \ML_int[6][1] ;
   wire \ML_int[6][0] ;
   wire n3;
   wire n4;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire [4:0] SHMAG;

   assign B[15] = \ML_int[6][15]  ;
   assign B[14] = \ML_int[6][14]  ;
   assign B[13] = \ML_int[6][13]  ;
   assign B[12] = \ML_int[6][12]  ;
   assign B[11] = \ML_int[6][11]  ;
   assign B[10] = \ML_int[6][10]  ;
   assign B[9] = \ML_int[6][9]  ;
   assign B[8] = \ML_int[6][8]  ;
   assign B[7] = \ML_int[6][7]  ;
   assign B[6] = \ML_int[6][6]  ;
   assign B[5] = \ML_int[6][5]  ;
   assign B[4] = \ML_int[6][4]  ;
   assign B[3] = \ML_int[6][3]  ;
   assign B[2] = \ML_int[6][2]  ;
   assign B[1] = \ML_int[6][1]  ;
   assign B[0] = \ML_int[6][0]  ;

   MX2X1 M1_0_15 (.Y(\ML_int[1][15] ), 
	.S0(n35), 
	.B(A[14]), 
	.A(A[15]));
   MX2X1 M1_1_15 (.Y(\ML_int[2][15] ), 
	.S0(n34), 
	.B(\ML_int[1][13] ), 
	.A(\ML_int[1][15] ));
   MX2X1 M1_2_15 (.Y(\ML_int[3][15] ), 
	.S0(n32), 
	.B(\ML_int[2][11] ), 
	.A(\ML_int[2][15] ));
   MX2X1 M1_3_15 (.Y(\ML_int[4][15] ), 
	.S0(n31), 
	.B(\ML_int[3][7] ), 
	.A(\ML_int[3][15] ));
   MX2X1 M1_0_14 (.Y(\ML_int[1][14] ), 
	.S0(n35), 
	.B(A[13]), 
	.A(A[14]));
   MX2X1 M1_0_1 (.Y(\ML_int[1][1] ), 
	.S0(n35), 
	.B(A[0]), 
	.A(A[1]));
   MX2X1 M1_0_2 (.Y(\ML_int[1][2] ), 
	.S0(n35), 
	.B(A[1]), 
	.A(A[2]));
   MX2X1 M1_0_4 (.Y(\ML_int[1][4] ), 
	.S0(n35), 
	.B(A[3]), 
	.A(A[4]));
   MX2X1 M1_0_5 (.Y(\ML_int[1][5] ), 
	.S0(n35), 
	.B(A[4]), 
	.A(A[5]));
   MX2X1 M1_0_13 (.Y(\ML_int[1][13] ), 
	.S0(n35), 
	.B(A[12]), 
	.A(A[13]));
   MX2X1 M1_0_11 (.Y(\ML_int[1][11] ), 
	.S0(n35), 
	.B(A[10]), 
	.A(A[11]));
   MX2X1 M1_0_9 (.Y(\ML_int[1][9] ), 
	.S0(n35), 
	.B(A[8]), 
	.A(A[9]));
   MX2X1 M1_0_12 (.Y(\ML_int[1][12] ), 
	.S0(n35), 
	.B(A[11]), 
	.A(A[12]));
   MX2X1 M1_0_8 (.Y(\ML_int[1][8] ), 
	.S0(n35), 
	.B(A[7]), 
	.A(A[8]));
   MX2X1 M1_0_10 (.Y(\ML_int[1][10] ), 
	.S0(n35), 
	.B(A[9]), 
	.A(A[10]));
   MX2X1 M1_0_7 (.Y(\ML_int[1][7] ), 
	.S0(n35), 
	.B(A[6]), 
	.A(A[7]));
   MX2X1 M1_0_3 (.Y(\ML_int[1][3] ), 
	.S0(n35), 
	.B(A[2]), 
	.A(A[3]));
   MX2X1 M1_0_6 (.Y(\ML_int[1][6] ), 
	.S0(n35), 
	.B(A[5]), 
	.A(A[6]));
   MX2X1 M1_1_14 (.Y(\ML_int[2][14] ), 
	.S0(n34), 
	.B(\ML_int[1][12] ), 
	.A(\ML_int[1][14] ));
   MX2X1 M1_2_14 (.Y(\ML_int[3][14] ), 
	.S0(n32), 
	.B(\ML_int[2][10] ), 
	.A(\ML_int[2][14] ));
   MX2X1 M1_3_14 (.Y(\ML_int[4][14] ), 
	.S0(n31), 
	.B(\ML_int[3][6] ), 
	.A(\ML_int[3][14] ));
   MX2X1 M1_1_13 (.Y(\ML_int[2][13] ), 
	.S0(n34), 
	.B(\ML_int[1][11] ), 
	.A(\ML_int[1][13] ));
   MX2X1 M1_2_13 (.Y(\ML_int[3][13] ), 
	.S0(n32), 
	.B(\ML_int[2][9] ), 
	.A(\ML_int[2][13] ));
   MX2X1 M1_3_13 (.Y(\ML_int[4][13] ), 
	.S0(n31), 
	.B(\ML_int[3][5] ), 
	.A(\ML_int[3][13] ));
   MX2X1 M1_1_12 (.Y(\ML_int[2][12] ), 
	.S0(n34), 
	.B(\ML_int[1][10] ), 
	.A(\ML_int[1][12] ));
   MX2X1 M1_2_12 (.Y(\ML_int[3][12] ), 
	.S0(n32), 
	.B(\ML_int[2][8] ), 
	.A(\ML_int[2][12] ));
   MX2X1 M1_3_12 (.Y(\ML_int[4][12] ), 
	.S0(n31), 
	.B(\ML_int[3][4] ), 
	.A(\ML_int[3][12] ));
   MX2X1 M1_1_11 (.Y(\ML_int[2][11] ), 
	.S0(n34), 
	.B(\ML_int[1][9] ), 
	.A(\ML_int[1][11] ));
   MX2X1 M1_1_7 (.Y(\ML_int[2][7] ), 
	.S0(n34), 
	.B(\ML_int[1][5] ), 
	.A(\ML_int[1][7] ));
   MX2X1 M1_1_8 (.Y(\ML_int[2][8] ), 
	.S0(n34), 
	.B(\ML_int[1][6] ), 
	.A(\ML_int[1][8] ));
   MX2X1 M1_1_4 (.Y(\ML_int[2][4] ), 
	.S0(n34), 
	.B(\ML_int[1][2] ), 
	.A(\ML_int[1][4] ));
   MX2X1 M1_1_10 (.Y(\ML_int[2][10] ), 
	.S0(n34), 
	.B(\ML_int[1][8] ), 
	.A(\ML_int[1][10] ));
   MX2X1 M1_1_9 (.Y(\ML_int[2][9] ), 
	.S0(n34), 
	.B(\ML_int[1][7] ), 
	.A(\ML_int[1][9] ));
   MX2X1 M1_1_6 (.Y(\ML_int[2][6] ), 
	.S0(n34), 
	.B(\ML_int[1][4] ), 
	.A(\ML_int[1][6] ));
   MX2X1 M1_1_5 (.Y(\ML_int[2][5] ), 
	.S0(n34), 
	.B(\ML_int[1][3] ), 
	.A(\ML_int[1][5] ));
   MX2X1 M1_1_2 (.Y(\ML_int[2][2] ), 
	.S0(n34), 
	.B(\ML_int[1][0] ), 
	.A(\ML_int[1][2] ));
   MX2X1 M1_1_3 (.Y(\ML_int[2][3] ), 
	.S0(n34), 
	.B(\ML_int[1][1] ), 
	.A(\ML_int[1][3] ));
   MX2X1 M1_3_8 (.Y(\ML_int[4][8] ), 
	.S0(n31), 
	.B(n33), 
	.A(\ML_int[3][8] ));
   MX2X1 M1_2_8 (.Y(\ML_int[3][8] ), 
	.S0(n32), 
	.B(\ML_int[2][4] ), 
	.A(\ML_int[2][8] ));
   MX2X1 M1_2_7 (.Y(\ML_int[3][7] ), 
	.S0(n32), 
	.B(\ML_int[2][3] ), 
	.A(\ML_int[2][7] ));
   MX2X1 M1_2_6 (.Y(\ML_int[3][6] ), 
	.S0(n32), 
	.B(\ML_int[2][2] ), 
	.A(\ML_int[2][6] ));
   MX2X1 M1_2_4 (.Y(\ML_int[3][4] ), 
	.S0(n32), 
	.B(\ML_int[2][0] ), 
	.A(\ML_int[2][4] ));
   MX2X1 M1_2_5 (.Y(\ML_int[3][5] ), 
	.S0(n32), 
	.B(\ML_int[2][1] ), 
	.A(\ML_int[2][5] ));
   AND2X2 U3 (.Y(\ML_int[6][11] ), 
	.B(n14), 
	.A(\ML_int[4][11] ));
   NOR2X1 U4 (.Y(\ML_int[6][1] ), 
	.B(n18), 
	.A(n15));
   NOR2X1 U5 (.Y(\ML_int[6][2] ), 
	.B(n17), 
	.A(n15));
   NOR2X1 U6 (.Y(\ML_int[6][3] ), 
	.B(n16), 
	.A(n15));
   NOR2BX1 U7 (.Y(\ML_int[6][4] ), 
	.B(n15), 
	.AN(\ML_int[3][4] ));
   NOR2BX1 U8 (.Y(\ML_int[6][7] ), 
	.B(n15), 
	.AN(\ML_int[3][7] ));
   NOR2BX1 U9 (.Y(\ML_int[6][6] ), 
	.B(n15), 
	.AN(\ML_int[3][6] ));
   NOR2BX1 U10 (.Y(\ML_int[6][5] ), 
	.B(n15), 
	.AN(\ML_int[3][5] ));
   INVX1 U11 (.Y(n33), 
	.A(n19));
   NAND2X1 U12 (.Y(n15), 
	.B(SHMAG[3]), 
	.A(n14));
   AND2X2 U13 (.Y(\ML_int[6][8] ), 
	.B(n14), 
	.A(\ML_int[4][8] ));
   NOR2X1 U14 (.Y(\ML_int[6][0] ), 
	.B(n19), 
	.A(n15));
   INVX1 U15 (.Y(n32), 
	.A(SHMAG[2]));
   INVX1 U16 (.Y(n35), 
	.A(SHMAG[0]));
   INVX1 U17 (.Y(n34), 
	.A(SHMAG[1]));
   NAND2X1 U18 (.Y(n16), 
	.B(SHMAG[2]), 
	.A(\ML_int[2][3] ));
   NAND2X1 U19 (.Y(n19), 
	.B(SHMAG[2]), 
	.A(\ML_int[2][0] ));
   INVX1 U20 (.Y(n31), 
	.A(SHMAG[3]));
   NAND2X1 U21 (.Y(n18), 
	.B(SHMAG[2]), 
	.A(\ML_int[2][1] ));
   NAND2X1 U22 (.Y(n17), 
	.B(SHMAG[2]), 
	.A(\ML_int[2][2] ));
   AND2X2 U23 (.Y(\ML_int[2][1] ), 
	.B(SHMAG[1]), 
	.A(\ML_int[1][1] ));
   AND2X2 U24 (.Y(\ML_int[2][0] ), 
	.B(SHMAG[1]), 
	.A(\ML_int[1][0] ));
   MXI2X1 U25 (.Y(\ML_int[4][11] ), 
	.S0(n31), 
	.B(n16), 
	.A(n30));
   MXI2X1 U26 (.Y(n30), 
	.S0(n32), 
	.B(\ML_int[2][7] ), 
	.A(\ML_int[2][11] ));
   AND2X2 U27 (.Y(\ML_int[6][12] ), 
	.B(n14), 
	.A(\ML_int[4][12] ));
   AND2X2 U28 (.Y(\ML_int[6][13] ), 
	.B(n14), 
	.A(\ML_int[4][13] ));
   AND2X2 U29 (.Y(\ML_int[6][14] ), 
	.B(n14), 
	.A(\ML_int[4][14] ));
   AND2X2 U30 (.Y(\ML_int[6][9] ), 
	.B(n14), 
	.A(\ML_int[4][9] ));
   MXI2X1 U31 (.Y(\ML_int[4][9] ), 
	.S0(n31), 
	.B(n18), 
	.A(n3));
   MXI2X1 U32 (.Y(n3), 
	.S0(n32), 
	.B(\ML_int[2][5] ), 
	.A(\ML_int[2][9] ));
   AND2X2 U33 (.Y(\ML_int[6][10] ), 
	.B(n14), 
	.A(\ML_int[4][10] ));
   MXI2X1 U34 (.Y(\ML_int[4][10] ), 
	.S0(n31), 
	.B(n17), 
	.A(n4));
   MXI2X1 U35 (.Y(n4), 
	.S0(n32), 
	.B(\ML_int[2][6] ), 
	.A(\ML_int[2][10] ));
   AOI21X1 U36 (.Y(SHMAG[2]), 
	.B0(n21), 
	.A1(n20), 
	.A0(SH[2]));
   AOI2BB1X1 U37 (.Y(n21), 
	.B0(SH[15]), 
	.A1N(n23), 
	.A0N(n22));
   OR4X2 U38 (.Y(n23), 
	.D(SH[12]), 
	.C(SH[11]), 
	.B(SH[10]), 
	.A(n24));
   NAND4X1 U39 (.Y(n22), 
	.D(n36), 
	.C(n25), 
	.B(n38), 
	.A(n37));
   OR2X2 U40 (.Y(n24), 
	.B(SH[13]), 
	.A(SH[14]));
   NOR2BX1 U41 (.Y(n14), 
	.B(SH[15]), 
	.AN(SHMAG[4]));
   AOI21X1 U42 (.Y(SHMAG[4]), 
	.B0(n21), 
	.A1(n20), 
	.A0(SH[4]));
   NAND2X1 U43 (.Y(n20), 
	.B(n26), 
	.A(SH[15]));
   NAND4BXL U44 (.Y(n26), 
	.D(n28), 
	.C(SH[8]), 
	.B(SH[9]), 
	.AN(n27));
   NAND3BX1 U45 (.Y(n27), 
	.C(SH[14]), 
	.B(SH[13]), 
	.AN(n29));
   NOR3X1 U46 (.Y(n28), 
	.C(n38), 
	.B(n37), 
	.A(n36));
   AOI21X1 U47 (.Y(SHMAG[3]), 
	.B0(n21), 
	.A1(n20), 
	.A0(SH[3]));
   AOI21X1 U48 (.Y(SHMAG[1]), 
	.B0(n21), 
	.A1(n20), 
	.A0(SH[1]));
   AOI21X1 U49 (.Y(SHMAG[0]), 
	.B0(n21), 
	.A1(n20), 
	.A0(SH[0]));
   NOR2X1 U50 (.Y(n25), 
	.B(SH[8]), 
	.A(SH[9]));
   AND2X2 U51 (.Y(\ML_int[6][15] ), 
	.B(n14), 
	.A(\ML_int[4][15] ));
   NAND3X1 U52 (.Y(n29), 
	.C(SH[12]), 
	.B(SH[10]), 
	.A(SH[11]));
   INVX1 U53 (.Y(n36), 
	.A(SH[7]));
   INVX1 U54 (.Y(n38), 
	.A(SH[6]));
   INVX1 U55 (.Y(n37), 
	.A(SH[5]));
   AND2X2 U56 (.Y(\ML_int[1][0] ), 
	.B(SHMAG[0]), 
	.A(A[0]));
endmodule

module alu (
	a, 
	b, 
	cmd, 
	r);
   input [15:0] a;
   input [15:0] b;
   input [2:0] cmd;
   output [15:0] r;

   // Internal wires
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N147;
   wire N148;
   wire N149;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire \U2/U2/Z_0 ;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;

   assign \U2/U2/Z_0  = cmd[0] ;

   alu_DW01_addsub_0 r71 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.B({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.CI(1'b0), 
	.ADD_SUB(\U2/U2/Z_0 ), 
	.SUM({ N66,
		N65,
		N64,
		N63,
		N62,
		N61,
		N60,
		N59,
		N58,
		N57,
		N56,
		N55,
		N54,
		N53,
		N52,
		N51 }));
   alu_DW_rash_0 srl_40 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.DATA_TC(1'b0), 
	.SH({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.SH_TC(1'b0), 
	.B({ N162,
		N161,
		N160,
		N159,
		N158,
		N157,
		N156,
		N155,
		N154,
		N153,
		N152,
		N151,
		N150,
		N149,
		N148,
		N147 }));
   alu_DW01_ash_0 sll_36 (.A({ a[15],
		a[14],
		a[13],
		a[12],
		a[11],
		a[10],
		a[9],
		a[8],
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }), 
	.DATA_TC(1'b0), 
	.SH({ b[15],
		b[14],
		b[13],
		b[12],
		b[11],
		b[10],
		b[9],
		b[8],
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }), 
	.SH_TC(1'b0), 
	.B({ N130,
		N129,
		N128,
		N127,
		N126,
		N125,
		N124,
		N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115 }));
   NAND4X1 U2 (.Y(r[9]), 
	.D(n228), 
	.C(n227), 
	.B(n226), 
	.A(n225));
   AOI211X1 U4 (.Y(n228), 
	.C0(n231), 
	.B0(n230), 
	.A1(n229), 
	.A0(a[9]));
   OAI21XL U7 (.Y(n229), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[9]));
   AOI22X1 U8 (.Y(n227), 
	.B1(n236), 
	.B0(n235), 
	.A1(n234), 
	.A0(b[9]));
   NAND2X1 U9 (.Y(n234), 
	.B(n233), 
	.A(n237));
   MXI2X1 U10 (.Y(n237), 
	.S0(a[9]), 
	.B(n239), 
	.A(n238));
   AOI222X1 U11 (.Y(n226), 
	.C1(n244), 
	.C0(n243), 
	.B1(n242), 
	.B0(n241), 
	.A1(n240), 
	.A0(N60));
   AOI22X1 U12 (.Y(n225), 
	.B1(n246), 
	.B0(N124), 
	.A1(n245), 
	.A0(N156));
   NAND4X1 U13 (.Y(r[8]), 
	.D(n250), 
	.C(n249), 
	.B(n248), 
	.A(n247));
   AOI211X1 U14 (.Y(n250), 
	.C0(n243), 
	.B0(n231), 
	.A1(n251), 
	.A0(a[8]));
   OAI21XL U15 (.Y(n251), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[8]));
   AOI22X1 U16 (.Y(n249), 
	.B1(n253), 
	.B0(n241), 
	.A1(n252), 
	.A0(b[8]));
   NAND2X1 U17 (.Y(n252), 
	.B(n233), 
	.A(n254));
   MXI2X1 U18 (.Y(n254), 
	.S0(a[8]), 
	.B(n239), 
	.A(n238));
   AOI22X1 U19 (.Y(n248), 
	.B1(n240), 
	.B0(N59), 
	.A1(n255), 
	.A0(n235));
   AOI22X1 U20 (.Y(n247), 
	.B1(n246), 
	.B0(N123), 
	.A1(n245), 
	.A0(N155));
   NAND3X1 U21 (.Y(r[7]), 
	.C(n258), 
	.B(n257), 
	.A(n256));
   AOI211X1 U22 (.Y(n258), 
	.C0(n261), 
	.B0(n260), 
	.A1(n259), 
	.A0(a[7]));
   AOI21X1 U23 (.Y(n261), 
	.B0(n263), 
	.A1(n233), 
	.A0(n262));
   INVX1 U24 (.Y(n263), 
	.A(b[7]));
   MXI2X1 U25 (.Y(n262), 
	.S0(a[7]), 
	.B(n239), 
	.A(n238));
   NAND3X1 U26 (.Y(n260), 
	.C(n266), 
	.B(n265), 
	.A(n264));
   NAND4X1 U27 (.Y(n266), 
	.D(b[3]), 
	.C(n269), 
	.B(n268), 
	.A(n267));
   NOR2X1 U28 (.Y(n269), 
	.B(n271), 
	.A(n270));
   OAI21XL U29 (.Y(n259), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[7]));
   AOI222X1 U30 (.Y(n257), 
	.C1(n273), 
	.C0(n241), 
	.B1(n272), 
	.B0(n235), 
	.A1(n240), 
	.A0(N58));
   AOI22X1 U31 (.Y(n256), 
	.B1(n246), 
	.B0(N122), 
	.A1(n245), 
	.A0(N154));
   NAND4X1 U32 (.Y(r[6]), 
	.D(n277), 
	.C(n276), 
	.B(n275), 
	.A(n274));
   AOI211X1 U33 (.Y(n277), 
	.C0(n243), 
	.B0(n279), 
	.A1(n278), 
	.A0(a[6]));
   OAI21XL U34 (.Y(n278), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[6]));
   AOI222X1 U35 (.Y(n276), 
	.C1(n284), 
	.C0(n283), 
	.B1(n282), 
	.B0(n281), 
	.A1(n280), 
	.A0(b[6]));
   NAND2X1 U36 (.Y(n280), 
	.B(n233), 
	.A(n285));
   MXI2X1 U37 (.Y(n285), 
	.S0(a[6]), 
	.B(n239), 
	.A(n238));
   AOI222X1 U38 (.Y(n275), 
	.C1(n287), 
	.C0(n241), 
	.B1(n286), 
	.B0(n235), 
	.A1(n240), 
	.A0(N57));
   AOI22X1 U39 (.Y(n274), 
	.B1(n246), 
	.B0(N121), 
	.A1(n245), 
	.A0(N153));
   NAND4X1 U40 (.Y(r[5]), 
	.D(n291), 
	.C(n290), 
	.B(n289), 
	.A(n288));
   AOI211X1 U41 (.Y(n291), 
	.C0(n243), 
	.B0(n279), 
	.A1(n292), 
	.A0(a[5]));
   OAI21XL U42 (.Y(n292), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[5]));
   AOI222X1 U43 (.Y(n290), 
	.C1(n242), 
	.C0(n283), 
	.B1(n244), 
	.B0(n281), 
	.A1(n293), 
	.A0(b[5]));
   INVX1 U44 (.Y(n281), 
	.A(n294));
   NAND2X1 U45 (.Y(n293), 
	.B(n233), 
	.A(n295));
   MXI2X1 U46 (.Y(n295), 
	.S0(a[5]), 
	.B(n239), 
	.A(n238));
   AOI222X1 U47 (.Y(n289), 
	.C1(n296), 
	.C0(n235), 
	.B1(n236), 
	.B0(n241), 
	.A1(n240), 
	.A0(N56));
   AOI22X1 U48 (.Y(n288), 
	.B1(n246), 
	.B0(N120), 
	.A1(n245), 
	.A0(N152));
   NAND4X1 U49 (.Y(r[4]), 
	.D(n300), 
	.C(n299), 
	.B(n298), 
	.A(n297));
   AOI221X1 U50 (.Y(n300), 
	.C0(n279), 
	.B1(n301), 
	.B0(a[4]), 
	.A1(n253), 
	.A0(n283));
   OAI21XL U51 (.Y(n301), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[4]));
   AOI22X1 U52 (.Y(n299), 
	.B1(n255), 
	.B0(n241), 
	.A1(n302), 
	.A0(b[4]));
   NAND2X1 U53 (.Y(n302), 
	.B(n233), 
	.A(n303));
   MXI2X1 U54 (.Y(n303), 
	.S0(a[4]), 
	.B(n239), 
	.A(n238));
   AOI222X1 U55 (.Y(n298), 
	.C1(n240), 
	.C0(N55), 
	.B1(n304), 
	.B0(n235), 
	.A1(n245), 
	.A0(N151));
   AOI21X1 U56 (.Y(n297), 
	.B0(n305), 
	.A1(n246), 
	.A0(N119));
   NAND4X1 U57 (.Y(r[3]), 
	.D(n309), 
	.C(n308), 
	.B(n307), 
	.A(n306));
   AOI211X1 U58 (.Y(n309), 
	.C0(n311), 
	.B0(n279), 
	.A1(n310), 
	.A0(a[3]));
   NOR3X1 U59 (.Y(n311), 
	.C(n314), 
	.B(n313), 
	.A(n312));
   NOR2X1 U60 (.Y(n279), 
	.B(n315), 
	.A(n265));
   OAI21XL U61 (.Y(n310), 
	.B0(n316), 
	.A1(n232), 
	.A0(b[3]));
   AOI221X1 U62 (.Y(n308), 
	.C0(n318), 
	.B1(n317), 
	.B0(n235), 
	.A1(n273), 
	.A0(n283));
   AOI21X1 U63 (.Y(n318), 
	.B0(n320), 
	.A1(n233), 
	.A0(n319));
   MXI2X1 U64 (.Y(n319), 
	.S0(a[3]), 
	.B(n239), 
	.A(n238));
   OAI222XL U65 (.Y(n317), 
	.C1(n325), 
	.C0(n244), 
	.B1(n324), 
	.B0(n323), 
	.A1(n322), 
	.A0(n321));
   AOI222X1 U66 (.Y(n307), 
	.C1(n240), 
	.C0(N54), 
	.B1(n272), 
	.B0(n241), 
	.A1(n245), 
	.A0(N150));
   OAI221XL U67 (.Y(n272), 
	.C0(n328), 
	.B1(n244), 
	.B0(n327), 
	.A1(n321), 
	.A0(n326));
   AOI22X1 U68 (.Y(n328), 
	.B1(n329), 
	.B0(a[8]), 
	.A1(n267), 
	.A0(a[7]));
   AOI21X1 U69 (.Y(n306), 
	.B0(n305), 
	.A1(n246), 
	.A0(N118));
   NAND4X1 U70 (.Y(r[2]), 
	.D(n333), 
	.C(n332), 
	.B(n331), 
	.A(n330));
   AOI21X1 U71 (.Y(n333), 
	.B0(n334), 
	.A1(n287), 
	.A0(n283));
   INVX1 U72 (.Y(n334), 
	.A(n335));
   AOI32X1 U73 (.Y(n335), 
	.B1(a[2]), 
	.B0(n338), 
	.A2(n337), 
	.A1(n282), 
	.A0(n336));
   OAI21XL U74 (.Y(n338), 
	.B0(n316), 
	.A1(b[2]), 
	.A0(n232));
   NOR2X1 U75 (.Y(n283), 
	.B(n314), 
	.A(n339));
   AOI22X1 U76 (.Y(n332), 
	.B1(n341), 
	.B0(b[2]), 
	.A1(n340), 
	.A0(n235));
   NAND3X1 U77 (.Y(n341), 
	.C(n343), 
	.B(n233), 
	.A(n342));
   MXI2X1 U78 (.Y(n343), 
	.S0(a[2]), 
	.B(n239), 
	.A(n238));
   NAND3X1 U79 (.Y(n342), 
	.C(n344), 
	.B(n284), 
	.A(n336));
   OAI222XL U80 (.Y(n340), 
	.C1(n322), 
	.C0(n244), 
	.B1(n345), 
	.B0(n323), 
	.A1(n324), 
	.A0(n321));
   INVX1 U81 (.Y(n322), 
	.A(a[5]));
   AOI222X1 U82 (.Y(n331), 
	.C1(n240), 
	.C0(N53), 
	.B1(n286), 
	.B0(n241), 
	.A1(n245), 
	.A0(N149));
   OAI221XL U83 (.Y(n286), 
	.C0(n347), 
	.B1(n244), 
	.B0(n326), 
	.A1(n346), 
	.A0(n321));
   AOI22X1 U84 (.Y(n347), 
	.B1(n329), 
	.B0(a[7]), 
	.A1(n267), 
	.A0(a[6]));
   INVX1 U85 (.Y(n326), 
	.A(a[9]));
   AOI21X1 U86 (.Y(n330), 
	.B0(n305), 
	.A1(n246), 
	.A0(N117));
   NAND4X1 U87 (.Y(r[1]), 
	.D(n351), 
	.C(n350), 
	.B(n349), 
	.A(n348));
   AOI222X1 U88 (.Y(n351), 
	.C1(n354), 
	.C0(n336), 
	.B1(n353), 
	.B0(a[1]), 
	.A1(n352), 
	.A0(n235));
   OAI221XL U89 (.Y(n354), 
	.C0(n357), 
	.B1(n313), 
	.B0(n356), 
	.A1(n339), 
	.A0(n355));
   NAND3X1 U90 (.Y(n357), 
	.C(n358), 
	.B(n242), 
	.A(b[3]));
   INVX1 U91 (.Y(n313), 
	.A(n337));
   INVX1 U92 (.Y(n356), 
	.A(n244));
   INVX1 U93 (.Y(n355), 
	.A(n236));
   OAI221XL U94 (.Y(n236), 
	.C0(n361), 
	.B1(n360), 
	.B0(n244), 
	.A1(n359), 
	.A0(n321));
   AOI22X1 U95 (.Y(n361), 
	.B1(n329), 
	.B0(a[10]), 
	.A1(a[9]), 
	.A0(n267));
   OAI21XL U96 (.Y(n353), 
	.B0(n316), 
	.A1(n232), 
	.A0(b[1]));
   AOI21X1 U97 (.Y(n316), 
	.B0(n362), 
	.A1(n235), 
	.A0(n267));
   OAI222XL U98 (.Y(n352), 
	.C1(n324), 
	.C0(n244), 
	.B1(n363), 
	.B0(n323), 
	.A1(n345), 
	.A0(n321));
   INVX1 U99 (.Y(n324), 
	.A(a[4]));
   AOI22X1 U100 (.Y(n350), 
	.B1(n296), 
	.B0(n241), 
	.A1(n364), 
	.A0(b[1]));
   OAI221XL U101 (.Y(n296), 
	.C0(n366), 
	.B1(n346), 
	.B0(n244), 
	.A1(n365), 
	.A0(n321));
   AOI22X1 U102 (.Y(n366), 
	.B1(n329), 
	.B0(a[6]), 
	.A1(n267), 
	.A0(a[5]));
   INVX1 U103 (.Y(n346), 
	.A(a[8]));
   NAND2X1 U104 (.Y(n364), 
	.B(n233), 
	.A(n367));
   MXI2X1 U105 (.Y(n367), 
	.S0(a[1]), 
	.B(n239), 
	.A(n238));
   AOI22X1 U106 (.Y(n349), 
	.B1(n245), 
	.B0(N148), 
	.A1(n240), 
	.A0(N52));
   AOI21X1 U107 (.Y(n348), 
	.B0(n305), 
	.A1(n246), 
	.A0(N116));
   NAND2X1 U108 (.Y(n305), 
	.B(n294), 
	.A(n264));
   NAND2X1 U109 (.Y(n294), 
	.B(n337), 
	.A(n268));
   NAND2X1 U110 (.Y(r[15]), 
	.B(n369), 
	.A(n368));
   AOI222X1 U111 (.Y(n369), 
	.C1(n371), 
	.C0(a[15]), 
	.B1(n370), 
	.B0(b[15]), 
	.A1(n240), 
	.A0(N66));
   OR3XL U112 (.Y(n371), 
	.C(n373), 
	.B(n372), 
	.A(n362));
   MXI2X1 U113 (.Y(n373), 
	.S0(b[15]), 
	.B(n374), 
	.A(n232));
   NOR3X1 U114 (.Y(n372), 
	.C(n270), 
	.B(n375), 
	.A(n314));
   AOI31X1 U115 (.Y(n375), 
	.B0(n376), 
	.A2(n267), 
	.A1(n320), 
	.A0(n315));
   INVX1 U116 (.Y(n362), 
	.A(n233));
   OAI21XL U117 (.Y(n370), 
	.B0(n233), 
	.A1(n232), 
	.A0(a[15]));
   AOI22X1 U118 (.Y(n368), 
	.B1(n246), 
	.B0(N130), 
	.A1(n245), 
	.A0(N162));
   NAND4X1 U119 (.Y(r[14]), 
	.D(n380), 
	.C(n379), 
	.B(n378), 
	.A(n377));
   AOI22X1 U120 (.Y(n380), 
	.B1(n382), 
	.B0(b[14]), 
	.A1(n381), 
	.A0(a[14]));
   NAND2X1 U121 (.Y(n382), 
	.B(n233), 
	.A(n383));
   MXI2X1 U122 (.Y(n383), 
	.S0(a[14]), 
	.B(n239), 
	.A(n238));
   OAI21XL U123 (.Y(n381), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[14]));
   AOI22X1 U124 (.Y(n379), 
	.B1(n284), 
	.B0(n235), 
	.A1(n282), 
	.A0(n230));
   AOI22X1 U125 (.Y(n378), 
	.B1(n245), 
	.B0(N161), 
	.A1(n240), 
	.A0(N65));
   AOI21X1 U126 (.Y(n377), 
	.B0(n384), 
	.A1(n246), 
	.A0(N129));
   NAND4X1 U127 (.Y(r[13]), 
	.D(n388), 
	.C(n387), 
	.B(n386), 
	.A(n385));
   AOI22X1 U128 (.Y(n388), 
	.B1(n390), 
	.B0(b[13]), 
	.A1(n389), 
	.A0(a[13]));
   NAND2X1 U129 (.Y(n390), 
	.B(n233), 
	.A(n391));
   MXI2X1 U130 (.Y(n391), 
	.S0(a[13]), 
	.B(n239), 
	.A(n238));
   OAI21XL U131 (.Y(n389), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[13]));
   AOI22X1 U132 (.Y(n387), 
	.B1(n244), 
	.B0(n230), 
	.A1(n242), 
	.A0(n235));
   OAI222XL U133 (.Y(n242), 
	.C1(n282), 
	.C0(n271), 
	.B1(n393), 
	.B0(n312), 
	.A1(n392), 
	.A0(n323));
   AOI22X1 U134 (.Y(n386), 
	.B1(n245), 
	.B0(N160), 
	.A1(n240), 
	.A0(N64));
   AOI21X1 U135 (.Y(n385), 
	.B0(n384), 
	.A1(n246), 
	.A0(N128));
   NAND4X1 U136 (.Y(r[12]), 
	.D(n397), 
	.C(n396), 
	.B(n395), 
	.A(n394));
   AOI21X1 U137 (.Y(n397), 
	.B0(n230), 
	.A1(n398), 
	.A0(a[12]));
   OAI21XL U138 (.Y(n398), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[12]));
   AOI22X1 U139 (.Y(n396), 
	.B1(n253), 
	.B0(n235), 
	.A1(n399), 
	.A0(b[12]));
   NAND2X1 U140 (.Y(n399), 
	.B(n233), 
	.A(n400));
   MXI2X1 U141 (.Y(n400), 
	.S0(a[12]), 
	.B(n239), 
	.A(n238));
   AOI22X1 U142 (.Y(n395), 
	.B1(n245), 
	.B0(N159), 
	.A1(n240), 
	.A0(N63));
   AOI21X1 U143 (.Y(n394), 
	.B0(n384), 
	.A1(n246), 
	.A0(N127));
   NAND4X1 U144 (.Y(r[11]), 
	.D(n404), 
	.C(n403), 
	.B(n402), 
	.A(n401));
   AOI211X1 U145 (.Y(n404), 
	.C0(n230), 
	.B0(n406), 
	.A1(n405), 
	.A0(a[11]));
   AOI21X1 U146 (.Y(n406), 
	.B0(n408), 
	.A1(n233), 
	.A0(n407));
   MXI2X1 U147 (.Y(n407), 
	.S0(a[11]), 
	.B(n239), 
	.A(n238));
   OAI21XL U148 (.Y(n405), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[11]));
   AOI22X1 U149 (.Y(n403), 
	.B1(n243), 
	.B0(n267), 
	.A1(n273), 
	.A0(n235));
   OAI221XL U150 (.Y(n273), 
	.C0(n409), 
	.B1(n392), 
	.B0(n244), 
	.A1(n393), 
	.A0(n321));
   AOI22X1 U151 (.Y(n409), 
	.B1(n329), 
	.B0(a[12]), 
	.A1(n267), 
	.A0(a[11]));
   AOI22X1 U152 (.Y(n402), 
	.B1(n245), 
	.B0(N158), 
	.A1(n240), 
	.A0(N62));
   AOI21X1 U153 (.Y(n401), 
	.B0(n384), 
	.A1(n246), 
	.A0(N126));
   OAI31X1 U154 (.Y(n384), 
	.B0(n265), 
	.A2(n314), 
	.A1(n271), 
	.A0(n410));
   NAND4X1 U155 (.Y(r[10]), 
	.D(n414), 
	.C(n413), 
	.B(n412), 
	.A(n411));
   AOI211X1 U156 (.Y(n414), 
	.C0(n231), 
	.B0(n230), 
	.A1(n415), 
	.A0(a[10]));
   INVX1 U157 (.Y(n231), 
	.A(n265));
   NAND3X1 U158 (.Y(n265), 
	.C(n344), 
	.B(a[15]), 
	.A(n336));
   NOR2X1 U159 (.Y(n230), 
	.B(b[2]), 
	.A(n264));
   OAI21XL U160 (.Y(n415), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[10]));
   AOI22X1 U161 (.Y(n413), 
	.B1(n284), 
	.B0(n241), 
	.A1(n416), 
	.A0(b[10]));
   MXI2X1 U162 (.Y(n284), 
	.S0(n312), 
	.B(n271), 
	.A(n392));
   NAND2X1 U163 (.Y(n416), 
	.B(n233), 
	.A(n417));
   MXI2X1 U164 (.Y(n417), 
	.S0(a[10]), 
	.B(n239), 
	.A(n238));
   AOI222X1 U165 (.Y(n412), 
	.C1(n287), 
	.C0(n235), 
	.B1(n282), 
	.B0(n243), 
	.A1(n240), 
	.A0(N61));
   OAI221XL U166 (.Y(n287), 
	.C0(n418), 
	.B1(n393), 
	.B0(n244), 
	.A1(n360), 
	.A0(n321));
   AOI22X1 U167 (.Y(n418), 
	.B1(n329), 
	.B0(a[11]), 
	.A1(n267), 
	.A0(a[10]));
   INVX1 U168 (.Y(n393), 
	.A(a[13]));
   INVX1 U169 (.Y(n360), 
	.A(a[12]));
   INVX1 U170 (.Y(n243), 
	.A(n264));
   NAND3X1 U171 (.Y(n264), 
	.C(n336), 
	.B(n320), 
	.A(n337));
   AOI22X1 U172 (.Y(n411), 
	.B1(n246), 
	.B0(N125), 
	.A1(n245), 
	.A0(N157));
   NAND4X1 U173 (.Y(r[0]), 
	.D(n422), 
	.C(n421), 
	.B(n420), 
	.A(n419));
   AOI22X1 U174 (.Y(n422), 
	.B1(n424), 
	.B0(n336), 
	.A1(n423), 
	.A0(a[0]));
   OAI21XL U175 (.Y(n424), 
	.B0(n426), 
	.A1(n339), 
	.A0(n425));
   AOI31X1 U176 (.Y(n426), 
	.B0(n337), 
	.A2(n358), 
	.A1(n253), 
	.A0(b[3]));
   NOR3X1 U177 (.Y(n337), 
	.C(n376), 
	.B(n270), 
	.A(n271));
   INVX1 U178 (.Y(n376), 
	.A(b[4]));
   INVX1 U179 (.Y(n358), 
	.A(n410));
   OAI221XL U180 (.Y(n253), 
	.C0(n427), 
	.B1(n244), 
	.B0(n271), 
	.A1(n392), 
	.A0(n321));
   AOI22X1 U181 (.Y(n427), 
	.B1(n329), 
	.B0(a[13]), 
	.A1(n267), 
	.A0(a[12]));
   INVX1 U182 (.Y(n271), 
	.A(a[15]));
   INVX1 U183 (.Y(n392), 
	.A(a[14]));
   NAND2X1 U184 (.Y(n339), 
	.B(n315), 
	.A(n344));
   INVX1 U185 (.Y(n315), 
	.A(b[2]));
   NOR2BX1 U186 (.Y(n344), 
	.B(n320), 
	.AN(n428));
   INVX1 U187 (.Y(n425), 
	.A(n255));
   OAI221XL U188 (.Y(n255), 
	.C0(n429), 
	.B1(n244), 
	.B0(n359), 
	.A1(n321), 
	.A0(n327));
   AOI22X1 U189 (.Y(n429), 
	.B1(a[9]), 
	.B0(n329), 
	.A1(n267), 
	.A0(a[8]));
   INVX1 U190 (.Y(n359), 
	.A(a[11]));
   INVX1 U191 (.Y(n327), 
	.A(a[10]));
   INVX1 U192 (.Y(n336), 
	.A(n314));
   OAI21XL U193 (.Y(n423), 
	.B0(n233), 
	.A1(n232), 
	.A0(b[0]));
   AOI22X1 U194 (.Y(n421), 
	.B1(n304), 
	.B0(n241), 
	.A1(n430), 
	.A0(b[0]));
   OAI221XL U195 (.Y(n304), 
	.C0(n431), 
	.B1(n365), 
	.B0(n244), 
	.A1(n325), 
	.A0(n321));
   AOI22X1 U196 (.Y(n431), 
	.B1(n329), 
	.B0(a[5]), 
	.A1(n267), 
	.A0(a[4]));
   INVX1 U197 (.Y(n365), 
	.A(a[7]));
   INVX1 U198 (.Y(n325), 
	.A(a[6]));
   NOR3X1 U199 (.Y(n241), 
	.C(n410), 
	.B(b[3]), 
	.A(n314));
   NAND2X1 U200 (.Y(n410), 
	.B(n428), 
	.A(b[2]));
   NAND2X1 U201 (.Y(n430), 
	.B(n233), 
	.A(n432));
   NAND2X1 U202 (.Y(n233), 
	.B(n239), 
	.A(\U2/U2/Z_0 ));
   MXI2X1 U203 (.Y(n432), 
	.S0(a[0]), 
	.B(n239), 
	.A(n238));
   INVX1 U204 (.Y(n239), 
	.A(n374));
   NAND2X1 U205 (.Y(n374), 
	.B(n433), 
	.A(cmd[1]));
   INVX1 U206 (.Y(n238), 
	.A(n232));
   NAND3X1 U207 (.Y(n232), 
	.C(cmd[2]), 
	.B(n435), 
	.A(n434));
   AOI22X1 U208 (.Y(n420), 
	.B1(n240), 
	.B0(N51), 
	.A1(n436), 
	.A0(n235));
   NOR2X1 U209 (.Y(n240), 
	.B(cmd[2]), 
	.A(cmd[1]));
   OAI221XL U210 (.Y(n436), 
	.C0(n437), 
	.B1(n345), 
	.B0(n244), 
	.A1(n363), 
	.A0(n321));
   AOI22X1 U211 (.Y(n437), 
	.B1(n329), 
	.B0(a[1]), 
	.A1(n267), 
	.A0(a[0]));
   INVX1 U212 (.Y(n329), 
	.A(n323));
   NAND2X1 U213 (.Y(n323), 
	.B(n282), 
	.A(b[0]));
   INVX1 U214 (.Y(n267), 
	.A(n312));
   NAND2X1 U215 (.Y(n312), 
	.B(n438), 
	.A(n282));
   INVX1 U216 (.Y(n282), 
	.A(b[1]));
   INVX1 U217 (.Y(n345), 
	.A(a[3]));
   NAND2X1 U218 (.Y(n244), 
	.B(b[0]), 
	.A(b[1]));
   INVX1 U219 (.Y(n363), 
	.A(a[2]));
   NAND2X1 U220 (.Y(n321), 
	.B(n438), 
	.A(b[1]));
   INVX1 U221 (.Y(n438), 
	.A(b[0]));
   AND3X1 U222 (.Y(n235), 
	.C(n268), 
	.B(n320), 
	.A(n428));
   NOR2X1 U223 (.Y(n268), 
	.B(b[2]), 
	.A(n314));
   NAND3X1 U224 (.Y(n314), 
	.C(cmd[2]), 
	.B(n434), 
	.A(cmd[1]));
   INVX1 U225 (.Y(n320), 
	.A(b[3]));
   NOR2X1 U226 (.Y(n428), 
	.B(b[4]), 
	.A(n270));
   NAND4BXL U227 (.Y(n270), 
	.D(n440), 
	.C(n439), 
	.B(n408), 
	.AN(b[10]));
   NOR4X1 U228 (.Y(n440), 
	.D(b[5]), 
	.C(b[6]), 
	.B(b[15]), 
	.A(n441));
   OR3XL U229 (.Y(n441), 
	.C(b[7]), 
	.B(b[9]), 
	.A(b[8]));
   NOR3X1 U230 (.Y(n439), 
	.C(b[13]), 
	.B(b[14]), 
	.A(b[12]));
   INVX1 U231 (.Y(n408), 
	.A(b[11]));
   AOI22X1 U232 (.Y(n419), 
	.B1(n246), 
	.B0(N115), 
	.A1(n245), 
	.A0(N147));
   NOR3X1 U233 (.Y(n246), 
	.C(n434), 
	.B(cmd[1]), 
	.A(n433));
   NOR3X1 U234 (.Y(n245), 
	.C(n434), 
	.B(n435), 
	.A(n433));
   INVX1 U235 (.Y(n434), 
	.A(\U2/U2/Z_0 ));
   INVX1 U236 (.Y(n435), 
	.A(cmd[1]));
   INVX1 U237 (.Y(n433), 
	.A(cmd[2]));
endmodule

module EX_stage (
	clk, 
	rst, 
	pipeline_reg_in, 
	pipeline_reg_out, 
	ex_op_dest);
   input clk;
   input rst;
   input [56:0] pipeline_reg_in;
   output [37:0] pipeline_reg_out;
   output [2:0] ex_op_dest;

   // Internal wires
   wire pipeline_reg_in_0;
   wire \pipeline_reg_in[3] ;
   wire \pipeline_reg_in[2] ;
   wire \pipeline_reg_in[1] ;
   wire n77;
   wire [15:0] ex_alu_result;

   assign pipeline_reg_in_0 = pipeline_reg_in[0] ;
   assign ex_op_dest[2] = \pipeline_reg_in[3]  ;
   assign \pipeline_reg_in[3]  = pipeline_reg_in[3] ;
   assign ex_op_dest[1] = \pipeline_reg_in[2]  ;
   assign \pipeline_reg_in[2]  = pipeline_reg_in[2] ;
   assign ex_op_dest[0] = \pipeline_reg_in[1]  ;
   assign \pipeline_reg_in[1]  = pipeline_reg_in[1] ;

   DFFTRX4 \pipeline_reg_out_reg[21]  (.RN(n77), 
	.Q(pipeline_reg_out[21]), 
	.D(pipeline_reg_in[21]), 
	.CK(clk));
   alu alu_inst (.a({ pipeline_reg_in[53],
		pipeline_reg_in[52],
		pipeline_reg_in[51],
		pipeline_reg_in[50],
		pipeline_reg_in[49],
		pipeline_reg_in[48],
		pipeline_reg_in[47],
		pipeline_reg_in[46],
		pipeline_reg_in[45],
		pipeline_reg_in[44],
		pipeline_reg_in[43],
		pipeline_reg_in[42],
		pipeline_reg_in[41],
		pipeline_reg_in[40],
		pipeline_reg_in[39],
		pipeline_reg_in[38] }), 
	.b({ pipeline_reg_in[37],
		pipeline_reg_in[36],
		pipeline_reg_in[35],
		pipeline_reg_in[34],
		pipeline_reg_in[33],
		pipeline_reg_in[32],
		pipeline_reg_in[31],
		pipeline_reg_in[30],
		pipeline_reg_in[29],
		pipeline_reg_in[28],
		pipeline_reg_in[27],
		pipeline_reg_in[26],
		pipeline_reg_in[25],
		pipeline_reg_in[24],
		pipeline_reg_in[23],
		pipeline_reg_in[22] }), 
	.cmd({ pipeline_reg_in[56],
		pipeline_reg_in[55],
		pipeline_reg_in[54] }), 
	.r({ ex_alu_result[15],
		ex_alu_result[14],
		ex_alu_result[13],
		ex_alu_result[12],
		ex_alu_result[11],
		ex_alu_result[10],
		ex_alu_result[9],
		ex_alu_result[8],
		ex_alu_result[7],
		ex_alu_result[6],
		ex_alu_result[5],
		ex_alu_result[4],
		ex_alu_result[3],
		ex_alu_result[2],
		ex_alu_result[1],
		ex_alu_result[0] }));
   DFFTRX1 \pipeline_reg_out_reg[6]  (.RN(n77), 
	.Q(pipeline_reg_out[6]), 
	.D(pipeline_reg_in[6]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[20]  (.RN(n77), 
	.Q(pipeline_reg_out[20]), 
	.D(pipeline_reg_in[20]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[19]  (.RN(n77), 
	.Q(pipeline_reg_out[19]), 
	.D(pipeline_reg_in[19]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[18]  (.RN(n77), 
	.Q(pipeline_reg_out[18]), 
	.D(pipeline_reg_in[18]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[17]  (.RN(n77), 
	.Q(pipeline_reg_out[17]), 
	.D(pipeline_reg_in[17]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[16]  (.RN(n77), 
	.Q(pipeline_reg_out[16]), 
	.D(pipeline_reg_in[16]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[15]  (.RN(n77), 
	.Q(pipeline_reg_out[15]), 
	.D(pipeline_reg_in[15]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[14]  (.RN(n77), 
	.Q(pipeline_reg_out[14]), 
	.D(pipeline_reg_in[14]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[13]  (.RN(n77), 
	.Q(pipeline_reg_out[13]), 
	.D(pipeline_reg_in[13]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[12]  (.RN(n77), 
	.Q(pipeline_reg_out[12]), 
	.D(pipeline_reg_in[12]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[11]  (.RN(n77), 
	.Q(pipeline_reg_out[11]), 
	.D(pipeline_reg_in[11]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[10]  (.RN(n77), 
	.Q(pipeline_reg_out[10]), 
	.D(pipeline_reg_in[10]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[9]  (.RN(n77), 
	.Q(pipeline_reg_out[9]), 
	.D(pipeline_reg_in[9]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[8]  (.RN(n77), 
	.Q(pipeline_reg_out[8]), 
	.D(pipeline_reg_in[8]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[7]  (.RN(n77), 
	.Q(pipeline_reg_out[7]), 
	.D(pipeline_reg_in[7]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[5]  (.RN(n77), 
	.Q(pipeline_reg_out[5]), 
	.D(pipeline_reg_in[5]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[26]  (.RN(n77), 
	.Q(pipeline_reg_out[26]), 
	.D(ex_alu_result[4]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[25]  (.RN(n77), 
	.Q(pipeline_reg_out[25]), 
	.D(ex_alu_result[3]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[23]  (.RN(n77), 
	.Q(pipeline_reg_out[23]), 
	.D(ex_alu_result[1]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[29]  (.RN(n77), 
	.Q(pipeline_reg_out[29]), 
	.D(ex_alu_result[7]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[3]  (.RN(n77), 
	.Q(pipeline_reg_out[3]), 
	.D(\pipeline_reg_in[3] ), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[2]  (.RN(n77), 
	.Q(pipeline_reg_out[2]), 
	.D(\pipeline_reg_in[2] ), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[1]  (.RN(n77), 
	.Q(pipeline_reg_out[1]), 
	.D(\pipeline_reg_in[1] ), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[27]  (.RN(n77), 
	.Q(pipeline_reg_out[27]), 
	.D(ex_alu_result[5]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[24]  (.RN(n77), 
	.Q(pipeline_reg_out[24]), 
	.D(ex_alu_result[2]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[28]  (.RN(n77), 
	.Q(pipeline_reg_out[28]), 
	.D(ex_alu_result[6]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[22]  (.RN(n77), 
	.Q(pipeline_reg_out[22]), 
	.D(ex_alu_result[0]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[37]  (.RN(n77), 
	.Q(pipeline_reg_out[37]), 
	.D(ex_alu_result[15]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[36]  (.RN(n77), 
	.Q(pipeline_reg_out[36]), 
	.D(ex_alu_result[14]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[35]  (.RN(n77), 
	.Q(pipeline_reg_out[35]), 
	.D(ex_alu_result[13]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[34]  (.RN(n77), 
	.Q(pipeline_reg_out[34]), 
	.D(ex_alu_result[12]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[33]  (.RN(n77), 
	.Q(pipeline_reg_out[33]), 
	.D(ex_alu_result[11]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[32]  (.RN(n77), 
	.Q(pipeline_reg_out[32]), 
	.D(ex_alu_result[10]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[31]  (.RN(n77), 
	.Q(pipeline_reg_out[31]), 
	.D(ex_alu_result[9]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[30]  (.RN(n77), 
	.Q(pipeline_reg_out[30]), 
	.D(ex_alu_result[8]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[4]  (.RN(n77), 
	.Q(pipeline_reg_out[4]), 
	.D(pipeline_reg_in[4]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[0]  (.RN(n77), 
	.Q(pipeline_reg_out[0]), 
	.D(pipeline_reg_in_0), 
	.CK(clk));
   INVX1 U3 (.Y(n77), 
	.A(rst));
endmodule

module data_mem (
	clk, 
	mem_access_addr, 
	mem_write_data, 
	mem_write_en, 
	mem_read_data);
   input clk;
   input [15:0] mem_access_addr;
   input [15:0] mem_write_data;
   input mem_write_en;
   output [15:0] mem_read_data;

   // Internal wires
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire \ram[255][15] ;
   wire \ram[255][14] ;
   wire \ram[255][13] ;
   wire \ram[255][12] ;
   wire \ram[255][11] ;
   wire \ram[255][10] ;
   wire \ram[255][9] ;
   wire \ram[255][8] ;
   wire \ram[255][7] ;
   wire \ram[255][6] ;
   wire \ram[255][5] ;
   wire \ram[255][4] ;
   wire \ram[255][3] ;
   wire \ram[255][2] ;
   wire \ram[255][1] ;
   wire \ram[255][0] ;
   wire \ram[254][15] ;
   wire \ram[254][14] ;
   wire \ram[254][13] ;
   wire \ram[254][12] ;
   wire \ram[254][11] ;
   wire \ram[254][10] ;
   wire \ram[254][9] ;
   wire \ram[254][8] ;
   wire \ram[254][7] ;
   wire \ram[254][6] ;
   wire \ram[254][5] ;
   wire \ram[254][4] ;
   wire \ram[254][3] ;
   wire \ram[254][2] ;
   wire \ram[254][1] ;
   wire \ram[254][0] ;
   wire \ram[253][15] ;
   wire \ram[253][14] ;
   wire \ram[253][13] ;
   wire \ram[253][12] ;
   wire \ram[253][11] ;
   wire \ram[253][10] ;
   wire \ram[253][9] ;
   wire \ram[253][8] ;
   wire \ram[253][7] ;
   wire \ram[253][6] ;
   wire \ram[253][5] ;
   wire \ram[253][4] ;
   wire \ram[253][3] ;
   wire \ram[253][2] ;
   wire \ram[253][1] ;
   wire \ram[253][0] ;
   wire \ram[252][15] ;
   wire \ram[252][14] ;
   wire \ram[252][13] ;
   wire \ram[252][12] ;
   wire \ram[252][11] ;
   wire \ram[252][10] ;
   wire \ram[252][9] ;
   wire \ram[252][8] ;
   wire \ram[252][7] ;
   wire \ram[252][6] ;
   wire \ram[252][5] ;
   wire \ram[252][4] ;
   wire \ram[252][3] ;
   wire \ram[252][2] ;
   wire \ram[252][1] ;
   wire \ram[252][0] ;
   wire \ram[251][15] ;
   wire \ram[251][14] ;
   wire \ram[251][13] ;
   wire \ram[251][12] ;
   wire \ram[251][11] ;
   wire \ram[251][10] ;
   wire \ram[251][9] ;
   wire \ram[251][8] ;
   wire \ram[251][7] ;
   wire \ram[251][6] ;
   wire \ram[251][5] ;
   wire \ram[251][4] ;
   wire \ram[251][3] ;
   wire \ram[251][2] ;
   wire \ram[251][1] ;
   wire \ram[251][0] ;
   wire \ram[250][15] ;
   wire \ram[250][14] ;
   wire \ram[250][13] ;
   wire \ram[250][12] ;
   wire \ram[250][11] ;
   wire \ram[250][10] ;
   wire \ram[250][9] ;
   wire \ram[250][8] ;
   wire \ram[250][7] ;
   wire \ram[250][6] ;
   wire \ram[250][5] ;
   wire \ram[250][4] ;
   wire \ram[250][3] ;
   wire \ram[250][2] ;
   wire \ram[250][1] ;
   wire \ram[250][0] ;
   wire \ram[249][15] ;
   wire \ram[249][14] ;
   wire \ram[249][13] ;
   wire \ram[249][12] ;
   wire \ram[249][11] ;
   wire \ram[249][10] ;
   wire \ram[249][9] ;
   wire \ram[249][8] ;
   wire \ram[249][7] ;
   wire \ram[249][6] ;
   wire \ram[249][5] ;
   wire \ram[249][4] ;
   wire \ram[249][3] ;
   wire \ram[249][2] ;
   wire \ram[249][1] ;
   wire \ram[249][0] ;
   wire \ram[248][15] ;
   wire \ram[248][14] ;
   wire \ram[248][13] ;
   wire \ram[248][12] ;
   wire \ram[248][11] ;
   wire \ram[248][10] ;
   wire \ram[248][9] ;
   wire \ram[248][8] ;
   wire \ram[248][7] ;
   wire \ram[248][6] ;
   wire \ram[248][5] ;
   wire \ram[248][4] ;
   wire \ram[248][3] ;
   wire \ram[248][2] ;
   wire \ram[248][1] ;
   wire \ram[248][0] ;
   wire \ram[247][15] ;
   wire \ram[247][14] ;
   wire \ram[247][13] ;
   wire \ram[247][12] ;
   wire \ram[247][11] ;
   wire \ram[247][10] ;
   wire \ram[247][9] ;
   wire \ram[247][8] ;
   wire \ram[247][7] ;
   wire \ram[247][6] ;
   wire \ram[247][5] ;
   wire \ram[247][4] ;
   wire \ram[247][3] ;
   wire \ram[247][2] ;
   wire \ram[247][1] ;
   wire \ram[247][0] ;
   wire \ram[246][15] ;
   wire \ram[246][14] ;
   wire \ram[246][13] ;
   wire \ram[246][12] ;
   wire \ram[246][11] ;
   wire \ram[246][10] ;
   wire \ram[246][9] ;
   wire \ram[246][8] ;
   wire \ram[246][7] ;
   wire \ram[246][6] ;
   wire \ram[246][5] ;
   wire \ram[246][4] ;
   wire \ram[246][3] ;
   wire \ram[246][2] ;
   wire \ram[246][1] ;
   wire \ram[246][0] ;
   wire \ram[245][15] ;
   wire \ram[245][14] ;
   wire \ram[245][13] ;
   wire \ram[245][12] ;
   wire \ram[245][11] ;
   wire \ram[245][10] ;
   wire \ram[245][9] ;
   wire \ram[245][8] ;
   wire \ram[245][7] ;
   wire \ram[245][6] ;
   wire \ram[245][5] ;
   wire \ram[245][4] ;
   wire \ram[245][3] ;
   wire \ram[245][2] ;
   wire \ram[245][1] ;
   wire \ram[245][0] ;
   wire \ram[244][15] ;
   wire \ram[244][14] ;
   wire \ram[244][13] ;
   wire \ram[244][12] ;
   wire \ram[244][11] ;
   wire \ram[244][10] ;
   wire \ram[244][9] ;
   wire \ram[244][8] ;
   wire \ram[244][7] ;
   wire \ram[244][6] ;
   wire \ram[244][5] ;
   wire \ram[244][4] ;
   wire \ram[244][3] ;
   wire \ram[244][2] ;
   wire \ram[244][1] ;
   wire \ram[244][0] ;
   wire \ram[243][15] ;
   wire \ram[243][14] ;
   wire \ram[243][13] ;
   wire \ram[243][12] ;
   wire \ram[243][11] ;
   wire \ram[243][10] ;
   wire \ram[243][9] ;
   wire \ram[243][8] ;
   wire \ram[243][7] ;
   wire \ram[243][6] ;
   wire \ram[243][5] ;
   wire \ram[243][4] ;
   wire \ram[243][3] ;
   wire \ram[243][2] ;
   wire \ram[243][1] ;
   wire \ram[243][0] ;
   wire \ram[242][15] ;
   wire \ram[242][14] ;
   wire \ram[242][13] ;
   wire \ram[242][12] ;
   wire \ram[242][11] ;
   wire \ram[242][10] ;
   wire \ram[242][9] ;
   wire \ram[242][8] ;
   wire \ram[242][7] ;
   wire \ram[242][6] ;
   wire \ram[242][5] ;
   wire \ram[242][4] ;
   wire \ram[242][3] ;
   wire \ram[242][2] ;
   wire \ram[242][1] ;
   wire \ram[242][0] ;
   wire \ram[241][15] ;
   wire \ram[241][14] ;
   wire \ram[241][13] ;
   wire \ram[241][12] ;
   wire \ram[241][11] ;
   wire \ram[241][10] ;
   wire \ram[241][9] ;
   wire \ram[241][8] ;
   wire \ram[241][7] ;
   wire \ram[241][6] ;
   wire \ram[241][5] ;
   wire \ram[241][4] ;
   wire \ram[241][3] ;
   wire \ram[241][2] ;
   wire \ram[241][1] ;
   wire \ram[241][0] ;
   wire \ram[240][15] ;
   wire \ram[240][14] ;
   wire \ram[240][13] ;
   wire \ram[240][12] ;
   wire \ram[240][11] ;
   wire \ram[240][10] ;
   wire \ram[240][9] ;
   wire \ram[240][8] ;
   wire \ram[240][7] ;
   wire \ram[240][6] ;
   wire \ram[240][5] ;
   wire \ram[240][4] ;
   wire \ram[240][3] ;
   wire \ram[240][2] ;
   wire \ram[240][1] ;
   wire \ram[240][0] ;
   wire \ram[239][15] ;
   wire \ram[239][14] ;
   wire \ram[239][13] ;
   wire \ram[239][12] ;
   wire \ram[239][11] ;
   wire \ram[239][10] ;
   wire \ram[239][9] ;
   wire \ram[239][8] ;
   wire \ram[239][7] ;
   wire \ram[239][6] ;
   wire \ram[239][5] ;
   wire \ram[239][4] ;
   wire \ram[239][3] ;
   wire \ram[239][2] ;
   wire \ram[239][1] ;
   wire \ram[239][0] ;
   wire \ram[238][15] ;
   wire \ram[238][14] ;
   wire \ram[238][13] ;
   wire \ram[238][12] ;
   wire \ram[238][11] ;
   wire \ram[238][10] ;
   wire \ram[238][9] ;
   wire \ram[238][8] ;
   wire \ram[238][7] ;
   wire \ram[238][6] ;
   wire \ram[238][5] ;
   wire \ram[238][4] ;
   wire \ram[238][3] ;
   wire \ram[238][2] ;
   wire \ram[238][1] ;
   wire \ram[238][0] ;
   wire \ram[237][15] ;
   wire \ram[237][14] ;
   wire \ram[237][13] ;
   wire \ram[237][12] ;
   wire \ram[237][11] ;
   wire \ram[237][10] ;
   wire \ram[237][9] ;
   wire \ram[237][8] ;
   wire \ram[237][7] ;
   wire \ram[237][6] ;
   wire \ram[237][5] ;
   wire \ram[237][4] ;
   wire \ram[237][3] ;
   wire \ram[237][2] ;
   wire \ram[237][1] ;
   wire \ram[237][0] ;
   wire \ram[236][15] ;
   wire \ram[236][14] ;
   wire \ram[236][13] ;
   wire \ram[236][12] ;
   wire \ram[236][11] ;
   wire \ram[236][10] ;
   wire \ram[236][9] ;
   wire \ram[236][8] ;
   wire \ram[236][7] ;
   wire \ram[236][6] ;
   wire \ram[236][5] ;
   wire \ram[236][4] ;
   wire \ram[236][3] ;
   wire \ram[236][2] ;
   wire \ram[236][1] ;
   wire \ram[236][0] ;
   wire \ram[235][15] ;
   wire \ram[235][14] ;
   wire \ram[235][13] ;
   wire \ram[235][12] ;
   wire \ram[235][11] ;
   wire \ram[235][10] ;
   wire \ram[235][9] ;
   wire \ram[235][8] ;
   wire \ram[235][7] ;
   wire \ram[235][6] ;
   wire \ram[235][5] ;
   wire \ram[235][4] ;
   wire \ram[235][3] ;
   wire \ram[235][2] ;
   wire \ram[235][1] ;
   wire \ram[235][0] ;
   wire \ram[234][15] ;
   wire \ram[234][14] ;
   wire \ram[234][13] ;
   wire \ram[234][12] ;
   wire \ram[234][11] ;
   wire \ram[234][10] ;
   wire \ram[234][9] ;
   wire \ram[234][8] ;
   wire \ram[234][7] ;
   wire \ram[234][6] ;
   wire \ram[234][5] ;
   wire \ram[234][4] ;
   wire \ram[234][3] ;
   wire \ram[234][2] ;
   wire \ram[234][1] ;
   wire \ram[234][0] ;
   wire \ram[233][15] ;
   wire \ram[233][14] ;
   wire \ram[233][13] ;
   wire \ram[233][12] ;
   wire \ram[233][11] ;
   wire \ram[233][10] ;
   wire \ram[233][9] ;
   wire \ram[233][8] ;
   wire \ram[233][7] ;
   wire \ram[233][6] ;
   wire \ram[233][5] ;
   wire \ram[233][4] ;
   wire \ram[233][3] ;
   wire \ram[233][2] ;
   wire \ram[233][1] ;
   wire \ram[233][0] ;
   wire \ram[232][15] ;
   wire \ram[232][14] ;
   wire \ram[232][13] ;
   wire \ram[232][12] ;
   wire \ram[232][11] ;
   wire \ram[232][10] ;
   wire \ram[232][9] ;
   wire \ram[232][8] ;
   wire \ram[232][7] ;
   wire \ram[232][6] ;
   wire \ram[232][5] ;
   wire \ram[232][4] ;
   wire \ram[232][3] ;
   wire \ram[232][2] ;
   wire \ram[232][1] ;
   wire \ram[232][0] ;
   wire \ram[231][15] ;
   wire \ram[231][14] ;
   wire \ram[231][13] ;
   wire \ram[231][12] ;
   wire \ram[231][11] ;
   wire \ram[231][10] ;
   wire \ram[231][9] ;
   wire \ram[231][8] ;
   wire \ram[231][7] ;
   wire \ram[231][6] ;
   wire \ram[231][5] ;
   wire \ram[231][4] ;
   wire \ram[231][3] ;
   wire \ram[231][2] ;
   wire \ram[231][1] ;
   wire \ram[231][0] ;
   wire \ram[230][15] ;
   wire \ram[230][14] ;
   wire \ram[230][13] ;
   wire \ram[230][12] ;
   wire \ram[230][11] ;
   wire \ram[230][10] ;
   wire \ram[230][9] ;
   wire \ram[230][8] ;
   wire \ram[230][7] ;
   wire \ram[230][6] ;
   wire \ram[230][5] ;
   wire \ram[230][4] ;
   wire \ram[230][3] ;
   wire \ram[230][2] ;
   wire \ram[230][1] ;
   wire \ram[230][0] ;
   wire \ram[229][15] ;
   wire \ram[229][14] ;
   wire \ram[229][13] ;
   wire \ram[229][12] ;
   wire \ram[229][11] ;
   wire \ram[229][10] ;
   wire \ram[229][9] ;
   wire \ram[229][8] ;
   wire \ram[229][7] ;
   wire \ram[229][6] ;
   wire \ram[229][5] ;
   wire \ram[229][4] ;
   wire \ram[229][3] ;
   wire \ram[229][2] ;
   wire \ram[229][1] ;
   wire \ram[229][0] ;
   wire \ram[228][15] ;
   wire \ram[228][14] ;
   wire \ram[228][13] ;
   wire \ram[228][12] ;
   wire \ram[228][11] ;
   wire \ram[228][10] ;
   wire \ram[228][9] ;
   wire \ram[228][8] ;
   wire \ram[228][7] ;
   wire \ram[228][6] ;
   wire \ram[228][5] ;
   wire \ram[228][4] ;
   wire \ram[228][3] ;
   wire \ram[228][2] ;
   wire \ram[228][1] ;
   wire \ram[228][0] ;
   wire \ram[227][15] ;
   wire \ram[227][14] ;
   wire \ram[227][13] ;
   wire \ram[227][12] ;
   wire \ram[227][11] ;
   wire \ram[227][10] ;
   wire \ram[227][9] ;
   wire \ram[227][8] ;
   wire \ram[227][7] ;
   wire \ram[227][6] ;
   wire \ram[227][5] ;
   wire \ram[227][4] ;
   wire \ram[227][3] ;
   wire \ram[227][2] ;
   wire \ram[227][1] ;
   wire \ram[227][0] ;
   wire \ram[226][15] ;
   wire \ram[226][14] ;
   wire \ram[226][13] ;
   wire \ram[226][12] ;
   wire \ram[226][11] ;
   wire \ram[226][10] ;
   wire \ram[226][9] ;
   wire \ram[226][8] ;
   wire \ram[226][7] ;
   wire \ram[226][6] ;
   wire \ram[226][5] ;
   wire \ram[226][4] ;
   wire \ram[226][3] ;
   wire \ram[226][2] ;
   wire \ram[226][1] ;
   wire \ram[226][0] ;
   wire \ram[225][15] ;
   wire \ram[225][14] ;
   wire \ram[225][13] ;
   wire \ram[225][12] ;
   wire \ram[225][11] ;
   wire \ram[225][10] ;
   wire \ram[225][9] ;
   wire \ram[225][8] ;
   wire \ram[225][7] ;
   wire \ram[225][6] ;
   wire \ram[225][5] ;
   wire \ram[225][4] ;
   wire \ram[225][3] ;
   wire \ram[225][2] ;
   wire \ram[225][1] ;
   wire \ram[225][0] ;
   wire \ram[224][15] ;
   wire \ram[224][14] ;
   wire \ram[224][13] ;
   wire \ram[224][12] ;
   wire \ram[224][11] ;
   wire \ram[224][10] ;
   wire \ram[224][9] ;
   wire \ram[224][8] ;
   wire \ram[224][7] ;
   wire \ram[224][6] ;
   wire \ram[224][5] ;
   wire \ram[224][4] ;
   wire \ram[224][3] ;
   wire \ram[224][2] ;
   wire \ram[224][1] ;
   wire \ram[224][0] ;
   wire \ram[223][15] ;
   wire \ram[223][14] ;
   wire \ram[223][13] ;
   wire \ram[223][12] ;
   wire \ram[223][11] ;
   wire \ram[223][10] ;
   wire \ram[223][9] ;
   wire \ram[223][8] ;
   wire \ram[223][7] ;
   wire \ram[223][6] ;
   wire \ram[223][5] ;
   wire \ram[223][4] ;
   wire \ram[223][3] ;
   wire \ram[223][2] ;
   wire \ram[223][1] ;
   wire \ram[223][0] ;
   wire \ram[222][15] ;
   wire \ram[222][14] ;
   wire \ram[222][13] ;
   wire \ram[222][12] ;
   wire \ram[222][11] ;
   wire \ram[222][10] ;
   wire \ram[222][9] ;
   wire \ram[222][8] ;
   wire \ram[222][7] ;
   wire \ram[222][6] ;
   wire \ram[222][5] ;
   wire \ram[222][4] ;
   wire \ram[222][3] ;
   wire \ram[222][2] ;
   wire \ram[222][1] ;
   wire \ram[222][0] ;
   wire \ram[221][15] ;
   wire \ram[221][14] ;
   wire \ram[221][13] ;
   wire \ram[221][12] ;
   wire \ram[221][11] ;
   wire \ram[221][10] ;
   wire \ram[221][9] ;
   wire \ram[221][8] ;
   wire \ram[221][7] ;
   wire \ram[221][6] ;
   wire \ram[221][5] ;
   wire \ram[221][4] ;
   wire \ram[221][3] ;
   wire \ram[221][2] ;
   wire \ram[221][1] ;
   wire \ram[221][0] ;
   wire \ram[220][15] ;
   wire \ram[220][14] ;
   wire \ram[220][13] ;
   wire \ram[220][12] ;
   wire \ram[220][11] ;
   wire \ram[220][10] ;
   wire \ram[220][9] ;
   wire \ram[220][8] ;
   wire \ram[220][7] ;
   wire \ram[220][6] ;
   wire \ram[220][5] ;
   wire \ram[220][4] ;
   wire \ram[220][3] ;
   wire \ram[220][2] ;
   wire \ram[220][1] ;
   wire \ram[220][0] ;
   wire \ram[219][15] ;
   wire \ram[219][14] ;
   wire \ram[219][13] ;
   wire \ram[219][12] ;
   wire \ram[219][11] ;
   wire \ram[219][10] ;
   wire \ram[219][9] ;
   wire \ram[219][8] ;
   wire \ram[219][7] ;
   wire \ram[219][6] ;
   wire \ram[219][5] ;
   wire \ram[219][4] ;
   wire \ram[219][3] ;
   wire \ram[219][2] ;
   wire \ram[219][1] ;
   wire \ram[219][0] ;
   wire \ram[218][15] ;
   wire \ram[218][14] ;
   wire \ram[218][13] ;
   wire \ram[218][12] ;
   wire \ram[218][11] ;
   wire \ram[218][10] ;
   wire \ram[218][9] ;
   wire \ram[218][8] ;
   wire \ram[218][7] ;
   wire \ram[218][6] ;
   wire \ram[218][5] ;
   wire \ram[218][4] ;
   wire \ram[218][3] ;
   wire \ram[218][2] ;
   wire \ram[218][1] ;
   wire \ram[218][0] ;
   wire \ram[217][15] ;
   wire \ram[217][14] ;
   wire \ram[217][13] ;
   wire \ram[217][12] ;
   wire \ram[217][11] ;
   wire \ram[217][10] ;
   wire \ram[217][9] ;
   wire \ram[217][8] ;
   wire \ram[217][7] ;
   wire \ram[217][6] ;
   wire \ram[217][5] ;
   wire \ram[217][4] ;
   wire \ram[217][3] ;
   wire \ram[217][2] ;
   wire \ram[217][1] ;
   wire \ram[217][0] ;
   wire \ram[216][15] ;
   wire \ram[216][14] ;
   wire \ram[216][13] ;
   wire \ram[216][12] ;
   wire \ram[216][11] ;
   wire \ram[216][10] ;
   wire \ram[216][9] ;
   wire \ram[216][8] ;
   wire \ram[216][7] ;
   wire \ram[216][6] ;
   wire \ram[216][5] ;
   wire \ram[216][4] ;
   wire \ram[216][3] ;
   wire \ram[216][2] ;
   wire \ram[216][1] ;
   wire \ram[216][0] ;
   wire \ram[215][15] ;
   wire \ram[215][14] ;
   wire \ram[215][13] ;
   wire \ram[215][12] ;
   wire \ram[215][11] ;
   wire \ram[215][10] ;
   wire \ram[215][9] ;
   wire \ram[215][8] ;
   wire \ram[215][7] ;
   wire \ram[215][6] ;
   wire \ram[215][5] ;
   wire \ram[215][4] ;
   wire \ram[215][3] ;
   wire \ram[215][2] ;
   wire \ram[215][1] ;
   wire \ram[215][0] ;
   wire \ram[214][15] ;
   wire \ram[214][14] ;
   wire \ram[214][13] ;
   wire \ram[214][12] ;
   wire \ram[214][11] ;
   wire \ram[214][10] ;
   wire \ram[214][9] ;
   wire \ram[214][8] ;
   wire \ram[214][7] ;
   wire \ram[214][6] ;
   wire \ram[214][5] ;
   wire \ram[214][4] ;
   wire \ram[214][3] ;
   wire \ram[214][2] ;
   wire \ram[214][1] ;
   wire \ram[214][0] ;
   wire \ram[213][15] ;
   wire \ram[213][14] ;
   wire \ram[213][13] ;
   wire \ram[213][12] ;
   wire \ram[213][11] ;
   wire \ram[213][10] ;
   wire \ram[213][9] ;
   wire \ram[213][8] ;
   wire \ram[213][7] ;
   wire \ram[213][6] ;
   wire \ram[213][5] ;
   wire \ram[213][4] ;
   wire \ram[213][3] ;
   wire \ram[213][2] ;
   wire \ram[213][1] ;
   wire \ram[213][0] ;
   wire \ram[212][15] ;
   wire \ram[212][14] ;
   wire \ram[212][13] ;
   wire \ram[212][12] ;
   wire \ram[212][11] ;
   wire \ram[212][10] ;
   wire \ram[212][9] ;
   wire \ram[212][8] ;
   wire \ram[212][7] ;
   wire \ram[212][6] ;
   wire \ram[212][5] ;
   wire \ram[212][4] ;
   wire \ram[212][3] ;
   wire \ram[212][2] ;
   wire \ram[212][1] ;
   wire \ram[212][0] ;
   wire \ram[211][15] ;
   wire \ram[211][14] ;
   wire \ram[211][13] ;
   wire \ram[211][12] ;
   wire \ram[211][11] ;
   wire \ram[211][10] ;
   wire \ram[211][9] ;
   wire \ram[211][8] ;
   wire \ram[211][7] ;
   wire \ram[211][6] ;
   wire \ram[211][5] ;
   wire \ram[211][4] ;
   wire \ram[211][3] ;
   wire \ram[211][2] ;
   wire \ram[211][1] ;
   wire \ram[211][0] ;
   wire \ram[210][15] ;
   wire \ram[210][14] ;
   wire \ram[210][13] ;
   wire \ram[210][12] ;
   wire \ram[210][11] ;
   wire \ram[210][10] ;
   wire \ram[210][9] ;
   wire \ram[210][8] ;
   wire \ram[210][7] ;
   wire \ram[210][6] ;
   wire \ram[210][5] ;
   wire \ram[210][4] ;
   wire \ram[210][3] ;
   wire \ram[210][2] ;
   wire \ram[210][1] ;
   wire \ram[210][0] ;
   wire \ram[209][15] ;
   wire \ram[209][14] ;
   wire \ram[209][13] ;
   wire \ram[209][12] ;
   wire \ram[209][11] ;
   wire \ram[209][10] ;
   wire \ram[209][9] ;
   wire \ram[209][8] ;
   wire \ram[209][7] ;
   wire \ram[209][6] ;
   wire \ram[209][5] ;
   wire \ram[209][4] ;
   wire \ram[209][3] ;
   wire \ram[209][2] ;
   wire \ram[209][1] ;
   wire \ram[209][0] ;
   wire \ram[208][15] ;
   wire \ram[208][14] ;
   wire \ram[208][13] ;
   wire \ram[208][12] ;
   wire \ram[208][11] ;
   wire \ram[208][10] ;
   wire \ram[208][9] ;
   wire \ram[208][8] ;
   wire \ram[208][7] ;
   wire \ram[208][6] ;
   wire \ram[208][5] ;
   wire \ram[208][4] ;
   wire \ram[208][3] ;
   wire \ram[208][2] ;
   wire \ram[208][1] ;
   wire \ram[208][0] ;
   wire \ram[207][15] ;
   wire \ram[207][14] ;
   wire \ram[207][13] ;
   wire \ram[207][12] ;
   wire \ram[207][11] ;
   wire \ram[207][10] ;
   wire \ram[207][9] ;
   wire \ram[207][8] ;
   wire \ram[207][7] ;
   wire \ram[207][6] ;
   wire \ram[207][5] ;
   wire \ram[207][4] ;
   wire \ram[207][3] ;
   wire \ram[207][2] ;
   wire \ram[207][1] ;
   wire \ram[207][0] ;
   wire \ram[206][15] ;
   wire \ram[206][14] ;
   wire \ram[206][13] ;
   wire \ram[206][12] ;
   wire \ram[206][11] ;
   wire \ram[206][10] ;
   wire \ram[206][9] ;
   wire \ram[206][8] ;
   wire \ram[206][7] ;
   wire \ram[206][6] ;
   wire \ram[206][5] ;
   wire \ram[206][4] ;
   wire \ram[206][3] ;
   wire \ram[206][2] ;
   wire \ram[206][1] ;
   wire \ram[206][0] ;
   wire \ram[205][15] ;
   wire \ram[205][14] ;
   wire \ram[205][13] ;
   wire \ram[205][12] ;
   wire \ram[205][11] ;
   wire \ram[205][10] ;
   wire \ram[205][9] ;
   wire \ram[205][8] ;
   wire \ram[205][7] ;
   wire \ram[205][6] ;
   wire \ram[205][5] ;
   wire \ram[205][4] ;
   wire \ram[205][3] ;
   wire \ram[205][2] ;
   wire \ram[205][1] ;
   wire \ram[205][0] ;
   wire \ram[204][15] ;
   wire \ram[204][14] ;
   wire \ram[204][13] ;
   wire \ram[204][12] ;
   wire \ram[204][11] ;
   wire \ram[204][10] ;
   wire \ram[204][9] ;
   wire \ram[204][8] ;
   wire \ram[204][7] ;
   wire \ram[204][6] ;
   wire \ram[204][5] ;
   wire \ram[204][4] ;
   wire \ram[204][3] ;
   wire \ram[204][2] ;
   wire \ram[204][1] ;
   wire \ram[204][0] ;
   wire \ram[203][15] ;
   wire \ram[203][14] ;
   wire \ram[203][13] ;
   wire \ram[203][12] ;
   wire \ram[203][11] ;
   wire \ram[203][10] ;
   wire \ram[203][9] ;
   wire \ram[203][8] ;
   wire \ram[203][7] ;
   wire \ram[203][6] ;
   wire \ram[203][5] ;
   wire \ram[203][4] ;
   wire \ram[203][3] ;
   wire \ram[203][2] ;
   wire \ram[203][1] ;
   wire \ram[203][0] ;
   wire \ram[202][15] ;
   wire \ram[202][14] ;
   wire \ram[202][13] ;
   wire \ram[202][12] ;
   wire \ram[202][11] ;
   wire \ram[202][10] ;
   wire \ram[202][9] ;
   wire \ram[202][8] ;
   wire \ram[202][7] ;
   wire \ram[202][6] ;
   wire \ram[202][5] ;
   wire \ram[202][4] ;
   wire \ram[202][3] ;
   wire \ram[202][2] ;
   wire \ram[202][1] ;
   wire \ram[202][0] ;
   wire \ram[201][15] ;
   wire \ram[201][14] ;
   wire \ram[201][13] ;
   wire \ram[201][12] ;
   wire \ram[201][11] ;
   wire \ram[201][10] ;
   wire \ram[201][9] ;
   wire \ram[201][8] ;
   wire \ram[201][7] ;
   wire \ram[201][6] ;
   wire \ram[201][5] ;
   wire \ram[201][4] ;
   wire \ram[201][3] ;
   wire \ram[201][2] ;
   wire \ram[201][1] ;
   wire \ram[201][0] ;
   wire \ram[200][15] ;
   wire \ram[200][14] ;
   wire \ram[200][13] ;
   wire \ram[200][12] ;
   wire \ram[200][11] ;
   wire \ram[200][10] ;
   wire \ram[200][9] ;
   wire \ram[200][8] ;
   wire \ram[200][7] ;
   wire \ram[200][6] ;
   wire \ram[200][5] ;
   wire \ram[200][4] ;
   wire \ram[200][3] ;
   wire \ram[200][2] ;
   wire \ram[200][1] ;
   wire \ram[200][0] ;
   wire \ram[199][15] ;
   wire \ram[199][14] ;
   wire \ram[199][13] ;
   wire \ram[199][12] ;
   wire \ram[199][11] ;
   wire \ram[199][10] ;
   wire \ram[199][9] ;
   wire \ram[199][8] ;
   wire \ram[199][7] ;
   wire \ram[199][6] ;
   wire \ram[199][5] ;
   wire \ram[199][4] ;
   wire \ram[199][3] ;
   wire \ram[199][2] ;
   wire \ram[199][1] ;
   wire \ram[199][0] ;
   wire \ram[198][15] ;
   wire \ram[198][14] ;
   wire \ram[198][13] ;
   wire \ram[198][12] ;
   wire \ram[198][11] ;
   wire \ram[198][10] ;
   wire \ram[198][9] ;
   wire \ram[198][8] ;
   wire \ram[198][7] ;
   wire \ram[198][6] ;
   wire \ram[198][5] ;
   wire \ram[198][4] ;
   wire \ram[198][3] ;
   wire \ram[198][2] ;
   wire \ram[198][1] ;
   wire \ram[198][0] ;
   wire \ram[197][15] ;
   wire \ram[197][14] ;
   wire \ram[197][13] ;
   wire \ram[197][12] ;
   wire \ram[197][11] ;
   wire \ram[197][10] ;
   wire \ram[197][9] ;
   wire \ram[197][8] ;
   wire \ram[197][7] ;
   wire \ram[197][6] ;
   wire \ram[197][5] ;
   wire \ram[197][4] ;
   wire \ram[197][3] ;
   wire \ram[197][2] ;
   wire \ram[197][1] ;
   wire \ram[197][0] ;
   wire \ram[196][15] ;
   wire \ram[196][14] ;
   wire \ram[196][13] ;
   wire \ram[196][12] ;
   wire \ram[196][11] ;
   wire \ram[196][10] ;
   wire \ram[196][9] ;
   wire \ram[196][8] ;
   wire \ram[196][7] ;
   wire \ram[196][6] ;
   wire \ram[196][5] ;
   wire \ram[196][4] ;
   wire \ram[196][3] ;
   wire \ram[196][2] ;
   wire \ram[196][1] ;
   wire \ram[196][0] ;
   wire \ram[195][15] ;
   wire \ram[195][14] ;
   wire \ram[195][13] ;
   wire \ram[195][12] ;
   wire \ram[195][11] ;
   wire \ram[195][10] ;
   wire \ram[195][9] ;
   wire \ram[195][8] ;
   wire \ram[195][7] ;
   wire \ram[195][6] ;
   wire \ram[195][5] ;
   wire \ram[195][4] ;
   wire \ram[195][3] ;
   wire \ram[195][2] ;
   wire \ram[195][1] ;
   wire \ram[195][0] ;
   wire \ram[194][15] ;
   wire \ram[194][14] ;
   wire \ram[194][13] ;
   wire \ram[194][12] ;
   wire \ram[194][11] ;
   wire \ram[194][10] ;
   wire \ram[194][9] ;
   wire \ram[194][8] ;
   wire \ram[194][7] ;
   wire \ram[194][6] ;
   wire \ram[194][5] ;
   wire \ram[194][4] ;
   wire \ram[194][3] ;
   wire \ram[194][2] ;
   wire \ram[194][1] ;
   wire \ram[194][0] ;
   wire \ram[193][15] ;
   wire \ram[193][14] ;
   wire \ram[193][13] ;
   wire \ram[193][12] ;
   wire \ram[193][11] ;
   wire \ram[193][10] ;
   wire \ram[193][9] ;
   wire \ram[193][8] ;
   wire \ram[193][7] ;
   wire \ram[193][6] ;
   wire \ram[193][5] ;
   wire \ram[193][4] ;
   wire \ram[193][3] ;
   wire \ram[193][2] ;
   wire \ram[193][1] ;
   wire \ram[193][0] ;
   wire \ram[192][15] ;
   wire \ram[192][14] ;
   wire \ram[192][13] ;
   wire \ram[192][12] ;
   wire \ram[192][11] ;
   wire \ram[192][10] ;
   wire \ram[192][9] ;
   wire \ram[192][8] ;
   wire \ram[192][7] ;
   wire \ram[192][6] ;
   wire \ram[192][5] ;
   wire \ram[192][4] ;
   wire \ram[192][3] ;
   wire \ram[192][2] ;
   wire \ram[192][1] ;
   wire \ram[192][0] ;
   wire \ram[191][15] ;
   wire \ram[191][14] ;
   wire \ram[191][13] ;
   wire \ram[191][12] ;
   wire \ram[191][11] ;
   wire \ram[191][10] ;
   wire \ram[191][9] ;
   wire \ram[191][8] ;
   wire \ram[191][7] ;
   wire \ram[191][6] ;
   wire \ram[191][5] ;
   wire \ram[191][4] ;
   wire \ram[191][3] ;
   wire \ram[191][2] ;
   wire \ram[191][1] ;
   wire \ram[191][0] ;
   wire \ram[190][15] ;
   wire \ram[190][14] ;
   wire \ram[190][13] ;
   wire \ram[190][12] ;
   wire \ram[190][11] ;
   wire \ram[190][10] ;
   wire \ram[190][9] ;
   wire \ram[190][8] ;
   wire \ram[190][7] ;
   wire \ram[190][6] ;
   wire \ram[190][5] ;
   wire \ram[190][4] ;
   wire \ram[190][3] ;
   wire \ram[190][2] ;
   wire \ram[190][1] ;
   wire \ram[190][0] ;
   wire \ram[189][15] ;
   wire \ram[189][14] ;
   wire \ram[189][13] ;
   wire \ram[189][12] ;
   wire \ram[189][11] ;
   wire \ram[189][10] ;
   wire \ram[189][9] ;
   wire \ram[189][8] ;
   wire \ram[189][7] ;
   wire \ram[189][6] ;
   wire \ram[189][5] ;
   wire \ram[189][4] ;
   wire \ram[189][3] ;
   wire \ram[189][2] ;
   wire \ram[189][1] ;
   wire \ram[189][0] ;
   wire \ram[188][15] ;
   wire \ram[188][14] ;
   wire \ram[188][13] ;
   wire \ram[188][12] ;
   wire \ram[188][11] ;
   wire \ram[188][10] ;
   wire \ram[188][9] ;
   wire \ram[188][8] ;
   wire \ram[188][7] ;
   wire \ram[188][6] ;
   wire \ram[188][5] ;
   wire \ram[188][4] ;
   wire \ram[188][3] ;
   wire \ram[188][2] ;
   wire \ram[188][1] ;
   wire \ram[188][0] ;
   wire \ram[187][15] ;
   wire \ram[187][14] ;
   wire \ram[187][13] ;
   wire \ram[187][12] ;
   wire \ram[187][11] ;
   wire \ram[187][10] ;
   wire \ram[187][9] ;
   wire \ram[187][8] ;
   wire \ram[187][7] ;
   wire \ram[187][6] ;
   wire \ram[187][5] ;
   wire \ram[187][4] ;
   wire \ram[187][3] ;
   wire \ram[187][2] ;
   wire \ram[187][1] ;
   wire \ram[187][0] ;
   wire \ram[186][15] ;
   wire \ram[186][14] ;
   wire \ram[186][13] ;
   wire \ram[186][12] ;
   wire \ram[186][11] ;
   wire \ram[186][10] ;
   wire \ram[186][9] ;
   wire \ram[186][8] ;
   wire \ram[186][7] ;
   wire \ram[186][6] ;
   wire \ram[186][5] ;
   wire \ram[186][4] ;
   wire \ram[186][3] ;
   wire \ram[186][2] ;
   wire \ram[186][1] ;
   wire \ram[186][0] ;
   wire \ram[185][15] ;
   wire \ram[185][14] ;
   wire \ram[185][13] ;
   wire \ram[185][12] ;
   wire \ram[185][11] ;
   wire \ram[185][10] ;
   wire \ram[185][9] ;
   wire \ram[185][8] ;
   wire \ram[185][7] ;
   wire \ram[185][6] ;
   wire \ram[185][5] ;
   wire \ram[185][4] ;
   wire \ram[185][3] ;
   wire \ram[185][2] ;
   wire \ram[185][1] ;
   wire \ram[185][0] ;
   wire \ram[184][15] ;
   wire \ram[184][14] ;
   wire \ram[184][13] ;
   wire \ram[184][12] ;
   wire \ram[184][11] ;
   wire \ram[184][10] ;
   wire \ram[184][9] ;
   wire \ram[184][8] ;
   wire \ram[184][7] ;
   wire \ram[184][6] ;
   wire \ram[184][5] ;
   wire \ram[184][4] ;
   wire \ram[184][3] ;
   wire \ram[184][2] ;
   wire \ram[184][1] ;
   wire \ram[184][0] ;
   wire \ram[183][15] ;
   wire \ram[183][14] ;
   wire \ram[183][13] ;
   wire \ram[183][12] ;
   wire \ram[183][11] ;
   wire \ram[183][10] ;
   wire \ram[183][9] ;
   wire \ram[183][8] ;
   wire \ram[183][7] ;
   wire \ram[183][6] ;
   wire \ram[183][5] ;
   wire \ram[183][4] ;
   wire \ram[183][3] ;
   wire \ram[183][2] ;
   wire \ram[183][1] ;
   wire \ram[183][0] ;
   wire \ram[182][15] ;
   wire \ram[182][14] ;
   wire \ram[182][13] ;
   wire \ram[182][12] ;
   wire \ram[182][11] ;
   wire \ram[182][10] ;
   wire \ram[182][9] ;
   wire \ram[182][8] ;
   wire \ram[182][7] ;
   wire \ram[182][6] ;
   wire \ram[182][5] ;
   wire \ram[182][4] ;
   wire \ram[182][3] ;
   wire \ram[182][2] ;
   wire \ram[182][1] ;
   wire \ram[182][0] ;
   wire \ram[181][15] ;
   wire \ram[181][14] ;
   wire \ram[181][13] ;
   wire \ram[181][12] ;
   wire \ram[181][11] ;
   wire \ram[181][10] ;
   wire \ram[181][9] ;
   wire \ram[181][8] ;
   wire \ram[181][7] ;
   wire \ram[181][6] ;
   wire \ram[181][5] ;
   wire \ram[181][4] ;
   wire \ram[181][3] ;
   wire \ram[181][2] ;
   wire \ram[181][1] ;
   wire \ram[181][0] ;
   wire \ram[180][15] ;
   wire \ram[180][14] ;
   wire \ram[180][13] ;
   wire \ram[180][12] ;
   wire \ram[180][11] ;
   wire \ram[180][10] ;
   wire \ram[180][9] ;
   wire \ram[180][8] ;
   wire \ram[180][7] ;
   wire \ram[180][6] ;
   wire \ram[180][5] ;
   wire \ram[180][4] ;
   wire \ram[180][3] ;
   wire \ram[180][2] ;
   wire \ram[180][1] ;
   wire \ram[180][0] ;
   wire \ram[179][15] ;
   wire \ram[179][14] ;
   wire \ram[179][13] ;
   wire \ram[179][12] ;
   wire \ram[179][11] ;
   wire \ram[179][10] ;
   wire \ram[179][9] ;
   wire \ram[179][8] ;
   wire \ram[179][7] ;
   wire \ram[179][6] ;
   wire \ram[179][5] ;
   wire \ram[179][4] ;
   wire \ram[179][3] ;
   wire \ram[179][2] ;
   wire \ram[179][1] ;
   wire \ram[179][0] ;
   wire \ram[178][15] ;
   wire \ram[178][14] ;
   wire \ram[178][13] ;
   wire \ram[178][12] ;
   wire \ram[178][11] ;
   wire \ram[178][10] ;
   wire \ram[178][9] ;
   wire \ram[178][8] ;
   wire \ram[178][7] ;
   wire \ram[178][6] ;
   wire \ram[178][5] ;
   wire \ram[178][4] ;
   wire \ram[178][3] ;
   wire \ram[178][2] ;
   wire \ram[178][1] ;
   wire \ram[178][0] ;
   wire \ram[177][15] ;
   wire \ram[177][14] ;
   wire \ram[177][13] ;
   wire \ram[177][12] ;
   wire \ram[177][11] ;
   wire \ram[177][10] ;
   wire \ram[177][9] ;
   wire \ram[177][8] ;
   wire \ram[177][7] ;
   wire \ram[177][6] ;
   wire \ram[177][5] ;
   wire \ram[177][4] ;
   wire \ram[177][3] ;
   wire \ram[177][2] ;
   wire \ram[177][1] ;
   wire \ram[177][0] ;
   wire \ram[176][15] ;
   wire \ram[176][14] ;
   wire \ram[176][13] ;
   wire \ram[176][12] ;
   wire \ram[176][11] ;
   wire \ram[176][10] ;
   wire \ram[176][9] ;
   wire \ram[176][8] ;
   wire \ram[176][7] ;
   wire \ram[176][6] ;
   wire \ram[176][5] ;
   wire \ram[176][4] ;
   wire \ram[176][3] ;
   wire \ram[176][2] ;
   wire \ram[176][1] ;
   wire \ram[176][0] ;
   wire \ram[175][15] ;
   wire \ram[175][14] ;
   wire \ram[175][13] ;
   wire \ram[175][12] ;
   wire \ram[175][11] ;
   wire \ram[175][10] ;
   wire \ram[175][9] ;
   wire \ram[175][8] ;
   wire \ram[175][7] ;
   wire \ram[175][6] ;
   wire \ram[175][5] ;
   wire \ram[175][4] ;
   wire \ram[175][3] ;
   wire \ram[175][2] ;
   wire \ram[175][1] ;
   wire \ram[175][0] ;
   wire \ram[174][15] ;
   wire \ram[174][14] ;
   wire \ram[174][13] ;
   wire \ram[174][12] ;
   wire \ram[174][11] ;
   wire \ram[174][10] ;
   wire \ram[174][9] ;
   wire \ram[174][8] ;
   wire \ram[174][7] ;
   wire \ram[174][6] ;
   wire \ram[174][5] ;
   wire \ram[174][4] ;
   wire \ram[174][3] ;
   wire \ram[174][2] ;
   wire \ram[174][1] ;
   wire \ram[174][0] ;
   wire \ram[173][15] ;
   wire \ram[173][14] ;
   wire \ram[173][13] ;
   wire \ram[173][12] ;
   wire \ram[173][11] ;
   wire \ram[173][10] ;
   wire \ram[173][9] ;
   wire \ram[173][8] ;
   wire \ram[173][7] ;
   wire \ram[173][6] ;
   wire \ram[173][5] ;
   wire \ram[173][4] ;
   wire \ram[173][3] ;
   wire \ram[173][2] ;
   wire \ram[173][1] ;
   wire \ram[173][0] ;
   wire \ram[172][15] ;
   wire \ram[172][14] ;
   wire \ram[172][13] ;
   wire \ram[172][12] ;
   wire \ram[172][11] ;
   wire \ram[172][10] ;
   wire \ram[172][9] ;
   wire \ram[172][8] ;
   wire \ram[172][7] ;
   wire \ram[172][6] ;
   wire \ram[172][5] ;
   wire \ram[172][4] ;
   wire \ram[172][3] ;
   wire \ram[172][2] ;
   wire \ram[172][1] ;
   wire \ram[172][0] ;
   wire \ram[171][15] ;
   wire \ram[171][14] ;
   wire \ram[171][13] ;
   wire \ram[171][12] ;
   wire \ram[171][11] ;
   wire \ram[171][10] ;
   wire \ram[171][9] ;
   wire \ram[171][8] ;
   wire \ram[171][7] ;
   wire \ram[171][6] ;
   wire \ram[171][5] ;
   wire \ram[171][4] ;
   wire \ram[171][3] ;
   wire \ram[171][2] ;
   wire \ram[171][1] ;
   wire \ram[171][0] ;
   wire \ram[170][15] ;
   wire \ram[170][14] ;
   wire \ram[170][13] ;
   wire \ram[170][12] ;
   wire \ram[170][11] ;
   wire \ram[170][10] ;
   wire \ram[170][9] ;
   wire \ram[170][8] ;
   wire \ram[170][7] ;
   wire \ram[170][6] ;
   wire \ram[170][5] ;
   wire \ram[170][4] ;
   wire \ram[170][3] ;
   wire \ram[170][2] ;
   wire \ram[170][1] ;
   wire \ram[170][0] ;
   wire \ram[169][15] ;
   wire \ram[169][14] ;
   wire \ram[169][13] ;
   wire \ram[169][12] ;
   wire \ram[169][11] ;
   wire \ram[169][10] ;
   wire \ram[169][9] ;
   wire \ram[169][8] ;
   wire \ram[169][7] ;
   wire \ram[169][6] ;
   wire \ram[169][5] ;
   wire \ram[169][4] ;
   wire \ram[169][3] ;
   wire \ram[169][2] ;
   wire \ram[169][1] ;
   wire \ram[169][0] ;
   wire \ram[168][15] ;
   wire \ram[168][14] ;
   wire \ram[168][13] ;
   wire \ram[168][12] ;
   wire \ram[168][11] ;
   wire \ram[168][10] ;
   wire \ram[168][9] ;
   wire \ram[168][8] ;
   wire \ram[168][7] ;
   wire \ram[168][6] ;
   wire \ram[168][5] ;
   wire \ram[168][4] ;
   wire \ram[168][3] ;
   wire \ram[168][2] ;
   wire \ram[168][1] ;
   wire \ram[168][0] ;
   wire \ram[167][15] ;
   wire \ram[167][14] ;
   wire \ram[167][13] ;
   wire \ram[167][12] ;
   wire \ram[167][11] ;
   wire \ram[167][10] ;
   wire \ram[167][9] ;
   wire \ram[167][8] ;
   wire \ram[167][7] ;
   wire \ram[167][6] ;
   wire \ram[167][5] ;
   wire \ram[167][4] ;
   wire \ram[167][3] ;
   wire \ram[167][2] ;
   wire \ram[167][1] ;
   wire \ram[167][0] ;
   wire \ram[166][15] ;
   wire \ram[166][14] ;
   wire \ram[166][13] ;
   wire \ram[166][12] ;
   wire \ram[166][11] ;
   wire \ram[166][10] ;
   wire \ram[166][9] ;
   wire \ram[166][8] ;
   wire \ram[166][7] ;
   wire \ram[166][6] ;
   wire \ram[166][5] ;
   wire \ram[166][4] ;
   wire \ram[166][3] ;
   wire \ram[166][2] ;
   wire \ram[166][1] ;
   wire \ram[166][0] ;
   wire \ram[165][15] ;
   wire \ram[165][14] ;
   wire \ram[165][13] ;
   wire \ram[165][12] ;
   wire \ram[165][11] ;
   wire \ram[165][10] ;
   wire \ram[165][9] ;
   wire \ram[165][8] ;
   wire \ram[165][7] ;
   wire \ram[165][6] ;
   wire \ram[165][5] ;
   wire \ram[165][4] ;
   wire \ram[165][3] ;
   wire \ram[165][2] ;
   wire \ram[165][1] ;
   wire \ram[165][0] ;
   wire \ram[164][15] ;
   wire \ram[164][14] ;
   wire \ram[164][13] ;
   wire \ram[164][12] ;
   wire \ram[164][11] ;
   wire \ram[164][10] ;
   wire \ram[164][9] ;
   wire \ram[164][8] ;
   wire \ram[164][7] ;
   wire \ram[164][6] ;
   wire \ram[164][5] ;
   wire \ram[164][4] ;
   wire \ram[164][3] ;
   wire \ram[164][2] ;
   wire \ram[164][1] ;
   wire \ram[164][0] ;
   wire \ram[163][15] ;
   wire \ram[163][14] ;
   wire \ram[163][13] ;
   wire \ram[163][12] ;
   wire \ram[163][11] ;
   wire \ram[163][10] ;
   wire \ram[163][9] ;
   wire \ram[163][8] ;
   wire \ram[163][7] ;
   wire \ram[163][6] ;
   wire \ram[163][5] ;
   wire \ram[163][4] ;
   wire \ram[163][3] ;
   wire \ram[163][2] ;
   wire \ram[163][1] ;
   wire \ram[163][0] ;
   wire \ram[162][15] ;
   wire \ram[162][14] ;
   wire \ram[162][13] ;
   wire \ram[162][12] ;
   wire \ram[162][11] ;
   wire \ram[162][10] ;
   wire \ram[162][9] ;
   wire \ram[162][8] ;
   wire \ram[162][7] ;
   wire \ram[162][6] ;
   wire \ram[162][5] ;
   wire \ram[162][4] ;
   wire \ram[162][3] ;
   wire \ram[162][2] ;
   wire \ram[162][1] ;
   wire \ram[162][0] ;
   wire \ram[161][15] ;
   wire \ram[161][14] ;
   wire \ram[161][13] ;
   wire \ram[161][12] ;
   wire \ram[161][11] ;
   wire \ram[161][10] ;
   wire \ram[161][9] ;
   wire \ram[161][8] ;
   wire \ram[161][7] ;
   wire \ram[161][6] ;
   wire \ram[161][5] ;
   wire \ram[161][4] ;
   wire \ram[161][3] ;
   wire \ram[161][2] ;
   wire \ram[161][1] ;
   wire \ram[161][0] ;
   wire \ram[160][15] ;
   wire \ram[160][14] ;
   wire \ram[160][13] ;
   wire \ram[160][12] ;
   wire \ram[160][11] ;
   wire \ram[160][10] ;
   wire \ram[160][9] ;
   wire \ram[160][8] ;
   wire \ram[160][7] ;
   wire \ram[160][6] ;
   wire \ram[160][5] ;
   wire \ram[160][4] ;
   wire \ram[160][3] ;
   wire \ram[160][2] ;
   wire \ram[160][1] ;
   wire \ram[160][0] ;
   wire \ram[159][15] ;
   wire \ram[159][14] ;
   wire \ram[159][13] ;
   wire \ram[159][12] ;
   wire \ram[159][11] ;
   wire \ram[159][10] ;
   wire \ram[159][9] ;
   wire \ram[159][8] ;
   wire \ram[159][7] ;
   wire \ram[159][6] ;
   wire \ram[159][5] ;
   wire \ram[159][4] ;
   wire \ram[159][3] ;
   wire \ram[159][2] ;
   wire \ram[159][1] ;
   wire \ram[159][0] ;
   wire \ram[158][15] ;
   wire \ram[158][14] ;
   wire \ram[158][13] ;
   wire \ram[158][12] ;
   wire \ram[158][11] ;
   wire \ram[158][10] ;
   wire \ram[158][9] ;
   wire \ram[158][8] ;
   wire \ram[158][7] ;
   wire \ram[158][6] ;
   wire \ram[158][5] ;
   wire \ram[158][4] ;
   wire \ram[158][3] ;
   wire \ram[158][2] ;
   wire \ram[158][1] ;
   wire \ram[158][0] ;
   wire \ram[157][15] ;
   wire \ram[157][14] ;
   wire \ram[157][13] ;
   wire \ram[157][12] ;
   wire \ram[157][11] ;
   wire \ram[157][10] ;
   wire \ram[157][9] ;
   wire \ram[157][8] ;
   wire \ram[157][7] ;
   wire \ram[157][6] ;
   wire \ram[157][5] ;
   wire \ram[157][4] ;
   wire \ram[157][3] ;
   wire \ram[157][2] ;
   wire \ram[157][1] ;
   wire \ram[157][0] ;
   wire \ram[156][15] ;
   wire \ram[156][14] ;
   wire \ram[156][13] ;
   wire \ram[156][12] ;
   wire \ram[156][11] ;
   wire \ram[156][10] ;
   wire \ram[156][9] ;
   wire \ram[156][8] ;
   wire \ram[156][7] ;
   wire \ram[156][6] ;
   wire \ram[156][5] ;
   wire \ram[156][4] ;
   wire \ram[156][3] ;
   wire \ram[156][2] ;
   wire \ram[156][1] ;
   wire \ram[156][0] ;
   wire \ram[155][15] ;
   wire \ram[155][14] ;
   wire \ram[155][13] ;
   wire \ram[155][12] ;
   wire \ram[155][11] ;
   wire \ram[155][10] ;
   wire \ram[155][9] ;
   wire \ram[155][8] ;
   wire \ram[155][7] ;
   wire \ram[155][6] ;
   wire \ram[155][5] ;
   wire \ram[155][4] ;
   wire \ram[155][3] ;
   wire \ram[155][2] ;
   wire \ram[155][1] ;
   wire \ram[155][0] ;
   wire \ram[154][15] ;
   wire \ram[154][14] ;
   wire \ram[154][13] ;
   wire \ram[154][12] ;
   wire \ram[154][11] ;
   wire \ram[154][10] ;
   wire \ram[154][9] ;
   wire \ram[154][8] ;
   wire \ram[154][7] ;
   wire \ram[154][6] ;
   wire \ram[154][5] ;
   wire \ram[154][4] ;
   wire \ram[154][3] ;
   wire \ram[154][2] ;
   wire \ram[154][1] ;
   wire \ram[154][0] ;
   wire \ram[153][15] ;
   wire \ram[153][14] ;
   wire \ram[153][13] ;
   wire \ram[153][12] ;
   wire \ram[153][11] ;
   wire \ram[153][10] ;
   wire \ram[153][9] ;
   wire \ram[153][8] ;
   wire \ram[153][7] ;
   wire \ram[153][6] ;
   wire \ram[153][5] ;
   wire \ram[153][4] ;
   wire \ram[153][3] ;
   wire \ram[153][2] ;
   wire \ram[153][1] ;
   wire \ram[153][0] ;
   wire \ram[152][15] ;
   wire \ram[152][14] ;
   wire \ram[152][13] ;
   wire \ram[152][12] ;
   wire \ram[152][11] ;
   wire \ram[152][10] ;
   wire \ram[152][9] ;
   wire \ram[152][8] ;
   wire \ram[152][7] ;
   wire \ram[152][6] ;
   wire \ram[152][5] ;
   wire \ram[152][4] ;
   wire \ram[152][3] ;
   wire \ram[152][2] ;
   wire \ram[152][1] ;
   wire \ram[152][0] ;
   wire \ram[151][15] ;
   wire \ram[151][14] ;
   wire \ram[151][13] ;
   wire \ram[151][12] ;
   wire \ram[151][11] ;
   wire \ram[151][10] ;
   wire \ram[151][9] ;
   wire \ram[151][8] ;
   wire \ram[151][7] ;
   wire \ram[151][6] ;
   wire \ram[151][5] ;
   wire \ram[151][4] ;
   wire \ram[151][3] ;
   wire \ram[151][2] ;
   wire \ram[151][1] ;
   wire \ram[151][0] ;
   wire \ram[150][15] ;
   wire \ram[150][14] ;
   wire \ram[150][13] ;
   wire \ram[150][12] ;
   wire \ram[150][11] ;
   wire \ram[150][10] ;
   wire \ram[150][9] ;
   wire \ram[150][8] ;
   wire \ram[150][7] ;
   wire \ram[150][6] ;
   wire \ram[150][5] ;
   wire \ram[150][4] ;
   wire \ram[150][3] ;
   wire \ram[150][2] ;
   wire \ram[150][1] ;
   wire \ram[150][0] ;
   wire \ram[149][15] ;
   wire \ram[149][14] ;
   wire \ram[149][13] ;
   wire \ram[149][12] ;
   wire \ram[149][11] ;
   wire \ram[149][10] ;
   wire \ram[149][9] ;
   wire \ram[149][8] ;
   wire \ram[149][7] ;
   wire \ram[149][6] ;
   wire \ram[149][5] ;
   wire \ram[149][4] ;
   wire \ram[149][3] ;
   wire \ram[149][2] ;
   wire \ram[149][1] ;
   wire \ram[149][0] ;
   wire \ram[148][15] ;
   wire \ram[148][14] ;
   wire \ram[148][13] ;
   wire \ram[148][12] ;
   wire \ram[148][11] ;
   wire \ram[148][10] ;
   wire \ram[148][9] ;
   wire \ram[148][8] ;
   wire \ram[148][7] ;
   wire \ram[148][6] ;
   wire \ram[148][5] ;
   wire \ram[148][4] ;
   wire \ram[148][3] ;
   wire \ram[148][2] ;
   wire \ram[148][1] ;
   wire \ram[148][0] ;
   wire \ram[147][15] ;
   wire \ram[147][14] ;
   wire \ram[147][13] ;
   wire \ram[147][12] ;
   wire \ram[147][11] ;
   wire \ram[147][10] ;
   wire \ram[147][9] ;
   wire \ram[147][8] ;
   wire \ram[147][7] ;
   wire \ram[147][6] ;
   wire \ram[147][5] ;
   wire \ram[147][4] ;
   wire \ram[147][3] ;
   wire \ram[147][2] ;
   wire \ram[147][1] ;
   wire \ram[147][0] ;
   wire \ram[146][15] ;
   wire \ram[146][14] ;
   wire \ram[146][13] ;
   wire \ram[146][12] ;
   wire \ram[146][11] ;
   wire \ram[146][10] ;
   wire \ram[146][9] ;
   wire \ram[146][8] ;
   wire \ram[146][7] ;
   wire \ram[146][6] ;
   wire \ram[146][5] ;
   wire \ram[146][4] ;
   wire \ram[146][3] ;
   wire \ram[146][2] ;
   wire \ram[146][1] ;
   wire \ram[146][0] ;
   wire \ram[145][15] ;
   wire \ram[145][14] ;
   wire \ram[145][13] ;
   wire \ram[145][12] ;
   wire \ram[145][11] ;
   wire \ram[145][10] ;
   wire \ram[145][9] ;
   wire \ram[145][8] ;
   wire \ram[145][7] ;
   wire \ram[145][6] ;
   wire \ram[145][5] ;
   wire \ram[145][4] ;
   wire \ram[145][3] ;
   wire \ram[145][2] ;
   wire \ram[145][1] ;
   wire \ram[145][0] ;
   wire \ram[144][15] ;
   wire \ram[144][14] ;
   wire \ram[144][13] ;
   wire \ram[144][12] ;
   wire \ram[144][11] ;
   wire \ram[144][10] ;
   wire \ram[144][9] ;
   wire \ram[144][8] ;
   wire \ram[144][7] ;
   wire \ram[144][6] ;
   wire \ram[144][5] ;
   wire \ram[144][4] ;
   wire \ram[144][3] ;
   wire \ram[144][2] ;
   wire \ram[144][1] ;
   wire \ram[144][0] ;
   wire \ram[143][15] ;
   wire \ram[143][14] ;
   wire \ram[143][13] ;
   wire \ram[143][12] ;
   wire \ram[143][11] ;
   wire \ram[143][10] ;
   wire \ram[143][9] ;
   wire \ram[143][8] ;
   wire \ram[143][7] ;
   wire \ram[143][6] ;
   wire \ram[143][5] ;
   wire \ram[143][4] ;
   wire \ram[143][3] ;
   wire \ram[143][2] ;
   wire \ram[143][1] ;
   wire \ram[143][0] ;
   wire \ram[142][15] ;
   wire \ram[142][14] ;
   wire \ram[142][13] ;
   wire \ram[142][12] ;
   wire \ram[142][11] ;
   wire \ram[142][10] ;
   wire \ram[142][9] ;
   wire \ram[142][8] ;
   wire \ram[142][7] ;
   wire \ram[142][6] ;
   wire \ram[142][5] ;
   wire \ram[142][4] ;
   wire \ram[142][3] ;
   wire \ram[142][2] ;
   wire \ram[142][1] ;
   wire \ram[142][0] ;
   wire \ram[141][15] ;
   wire \ram[141][14] ;
   wire \ram[141][13] ;
   wire \ram[141][12] ;
   wire \ram[141][11] ;
   wire \ram[141][10] ;
   wire \ram[141][9] ;
   wire \ram[141][8] ;
   wire \ram[141][7] ;
   wire \ram[141][6] ;
   wire \ram[141][5] ;
   wire \ram[141][4] ;
   wire \ram[141][3] ;
   wire \ram[141][2] ;
   wire \ram[141][1] ;
   wire \ram[141][0] ;
   wire \ram[140][15] ;
   wire \ram[140][14] ;
   wire \ram[140][13] ;
   wire \ram[140][12] ;
   wire \ram[140][11] ;
   wire \ram[140][10] ;
   wire \ram[140][9] ;
   wire \ram[140][8] ;
   wire \ram[140][7] ;
   wire \ram[140][6] ;
   wire \ram[140][5] ;
   wire \ram[140][4] ;
   wire \ram[140][3] ;
   wire \ram[140][2] ;
   wire \ram[140][1] ;
   wire \ram[140][0] ;
   wire \ram[139][15] ;
   wire \ram[139][14] ;
   wire \ram[139][13] ;
   wire \ram[139][12] ;
   wire \ram[139][11] ;
   wire \ram[139][10] ;
   wire \ram[139][9] ;
   wire \ram[139][8] ;
   wire \ram[139][7] ;
   wire \ram[139][6] ;
   wire \ram[139][5] ;
   wire \ram[139][4] ;
   wire \ram[139][3] ;
   wire \ram[139][2] ;
   wire \ram[139][1] ;
   wire \ram[139][0] ;
   wire \ram[138][15] ;
   wire \ram[138][14] ;
   wire \ram[138][13] ;
   wire \ram[138][12] ;
   wire \ram[138][11] ;
   wire \ram[138][10] ;
   wire \ram[138][9] ;
   wire \ram[138][8] ;
   wire \ram[138][7] ;
   wire \ram[138][6] ;
   wire \ram[138][5] ;
   wire \ram[138][4] ;
   wire \ram[138][3] ;
   wire \ram[138][2] ;
   wire \ram[138][1] ;
   wire \ram[138][0] ;
   wire \ram[137][15] ;
   wire \ram[137][14] ;
   wire \ram[137][13] ;
   wire \ram[137][12] ;
   wire \ram[137][11] ;
   wire \ram[137][10] ;
   wire \ram[137][9] ;
   wire \ram[137][8] ;
   wire \ram[137][7] ;
   wire \ram[137][6] ;
   wire \ram[137][5] ;
   wire \ram[137][4] ;
   wire \ram[137][3] ;
   wire \ram[137][2] ;
   wire \ram[137][1] ;
   wire \ram[137][0] ;
   wire \ram[136][15] ;
   wire \ram[136][14] ;
   wire \ram[136][13] ;
   wire \ram[136][12] ;
   wire \ram[136][11] ;
   wire \ram[136][10] ;
   wire \ram[136][9] ;
   wire \ram[136][8] ;
   wire \ram[136][7] ;
   wire \ram[136][6] ;
   wire \ram[136][5] ;
   wire \ram[136][4] ;
   wire \ram[136][3] ;
   wire \ram[136][2] ;
   wire \ram[136][1] ;
   wire \ram[136][0] ;
   wire \ram[135][15] ;
   wire \ram[135][14] ;
   wire \ram[135][13] ;
   wire \ram[135][12] ;
   wire \ram[135][11] ;
   wire \ram[135][10] ;
   wire \ram[135][9] ;
   wire \ram[135][8] ;
   wire \ram[135][7] ;
   wire \ram[135][6] ;
   wire \ram[135][5] ;
   wire \ram[135][4] ;
   wire \ram[135][3] ;
   wire \ram[135][2] ;
   wire \ram[135][1] ;
   wire \ram[135][0] ;
   wire \ram[134][15] ;
   wire \ram[134][14] ;
   wire \ram[134][13] ;
   wire \ram[134][12] ;
   wire \ram[134][11] ;
   wire \ram[134][10] ;
   wire \ram[134][9] ;
   wire \ram[134][8] ;
   wire \ram[134][7] ;
   wire \ram[134][6] ;
   wire \ram[134][5] ;
   wire \ram[134][4] ;
   wire \ram[134][3] ;
   wire \ram[134][2] ;
   wire \ram[134][1] ;
   wire \ram[134][0] ;
   wire \ram[133][15] ;
   wire \ram[133][14] ;
   wire \ram[133][13] ;
   wire \ram[133][12] ;
   wire \ram[133][11] ;
   wire \ram[133][10] ;
   wire \ram[133][9] ;
   wire \ram[133][8] ;
   wire \ram[133][7] ;
   wire \ram[133][6] ;
   wire \ram[133][5] ;
   wire \ram[133][4] ;
   wire \ram[133][3] ;
   wire \ram[133][2] ;
   wire \ram[133][1] ;
   wire \ram[133][0] ;
   wire \ram[132][15] ;
   wire \ram[132][14] ;
   wire \ram[132][13] ;
   wire \ram[132][12] ;
   wire \ram[132][11] ;
   wire \ram[132][10] ;
   wire \ram[132][9] ;
   wire \ram[132][8] ;
   wire \ram[132][7] ;
   wire \ram[132][6] ;
   wire \ram[132][5] ;
   wire \ram[132][4] ;
   wire \ram[132][3] ;
   wire \ram[132][2] ;
   wire \ram[132][1] ;
   wire \ram[132][0] ;
   wire \ram[131][15] ;
   wire \ram[131][14] ;
   wire \ram[131][13] ;
   wire \ram[131][12] ;
   wire \ram[131][11] ;
   wire \ram[131][10] ;
   wire \ram[131][9] ;
   wire \ram[131][8] ;
   wire \ram[131][7] ;
   wire \ram[131][6] ;
   wire \ram[131][5] ;
   wire \ram[131][4] ;
   wire \ram[131][3] ;
   wire \ram[131][2] ;
   wire \ram[131][1] ;
   wire \ram[131][0] ;
   wire \ram[130][15] ;
   wire \ram[130][14] ;
   wire \ram[130][13] ;
   wire \ram[130][12] ;
   wire \ram[130][11] ;
   wire \ram[130][10] ;
   wire \ram[130][9] ;
   wire \ram[130][8] ;
   wire \ram[130][7] ;
   wire \ram[130][6] ;
   wire \ram[130][5] ;
   wire \ram[130][4] ;
   wire \ram[130][3] ;
   wire \ram[130][2] ;
   wire \ram[130][1] ;
   wire \ram[130][0] ;
   wire \ram[129][15] ;
   wire \ram[129][14] ;
   wire \ram[129][13] ;
   wire \ram[129][12] ;
   wire \ram[129][11] ;
   wire \ram[129][10] ;
   wire \ram[129][9] ;
   wire \ram[129][8] ;
   wire \ram[129][7] ;
   wire \ram[129][6] ;
   wire \ram[129][5] ;
   wire \ram[129][4] ;
   wire \ram[129][3] ;
   wire \ram[129][2] ;
   wire \ram[129][1] ;
   wire \ram[129][0] ;
   wire \ram[128][15] ;
   wire \ram[128][14] ;
   wire \ram[128][13] ;
   wire \ram[128][12] ;
   wire \ram[128][11] ;
   wire \ram[128][10] ;
   wire \ram[128][9] ;
   wire \ram[128][8] ;
   wire \ram[128][7] ;
   wire \ram[128][6] ;
   wire \ram[128][5] ;
   wire \ram[128][4] ;
   wire \ram[128][3] ;
   wire \ram[128][2] ;
   wire \ram[128][1] ;
   wire \ram[128][0] ;
   wire \ram[127][15] ;
   wire \ram[127][14] ;
   wire \ram[127][13] ;
   wire \ram[127][12] ;
   wire \ram[127][11] ;
   wire \ram[127][10] ;
   wire \ram[127][9] ;
   wire \ram[127][8] ;
   wire \ram[127][7] ;
   wire \ram[127][6] ;
   wire \ram[127][5] ;
   wire \ram[127][4] ;
   wire \ram[127][3] ;
   wire \ram[127][2] ;
   wire \ram[127][1] ;
   wire \ram[127][0] ;
   wire \ram[126][15] ;
   wire \ram[126][14] ;
   wire \ram[126][13] ;
   wire \ram[126][12] ;
   wire \ram[126][11] ;
   wire \ram[126][10] ;
   wire \ram[126][9] ;
   wire \ram[126][8] ;
   wire \ram[126][7] ;
   wire \ram[126][6] ;
   wire \ram[126][5] ;
   wire \ram[126][4] ;
   wire \ram[126][3] ;
   wire \ram[126][2] ;
   wire \ram[126][1] ;
   wire \ram[126][0] ;
   wire \ram[125][15] ;
   wire \ram[125][14] ;
   wire \ram[125][13] ;
   wire \ram[125][12] ;
   wire \ram[125][11] ;
   wire \ram[125][10] ;
   wire \ram[125][9] ;
   wire \ram[125][8] ;
   wire \ram[125][7] ;
   wire \ram[125][6] ;
   wire \ram[125][5] ;
   wire \ram[125][4] ;
   wire \ram[125][3] ;
   wire \ram[125][2] ;
   wire \ram[125][1] ;
   wire \ram[125][0] ;
   wire \ram[124][15] ;
   wire \ram[124][14] ;
   wire \ram[124][13] ;
   wire \ram[124][12] ;
   wire \ram[124][11] ;
   wire \ram[124][10] ;
   wire \ram[124][9] ;
   wire \ram[124][8] ;
   wire \ram[124][7] ;
   wire \ram[124][6] ;
   wire \ram[124][5] ;
   wire \ram[124][4] ;
   wire \ram[124][3] ;
   wire \ram[124][2] ;
   wire \ram[124][1] ;
   wire \ram[124][0] ;
   wire \ram[123][15] ;
   wire \ram[123][14] ;
   wire \ram[123][13] ;
   wire \ram[123][12] ;
   wire \ram[123][11] ;
   wire \ram[123][10] ;
   wire \ram[123][9] ;
   wire \ram[123][8] ;
   wire \ram[123][7] ;
   wire \ram[123][6] ;
   wire \ram[123][5] ;
   wire \ram[123][4] ;
   wire \ram[123][3] ;
   wire \ram[123][2] ;
   wire \ram[123][1] ;
   wire \ram[123][0] ;
   wire \ram[122][15] ;
   wire \ram[122][14] ;
   wire \ram[122][13] ;
   wire \ram[122][12] ;
   wire \ram[122][11] ;
   wire \ram[122][10] ;
   wire \ram[122][9] ;
   wire \ram[122][8] ;
   wire \ram[122][7] ;
   wire \ram[122][6] ;
   wire \ram[122][5] ;
   wire \ram[122][4] ;
   wire \ram[122][3] ;
   wire \ram[122][2] ;
   wire \ram[122][1] ;
   wire \ram[122][0] ;
   wire \ram[121][15] ;
   wire \ram[121][14] ;
   wire \ram[121][13] ;
   wire \ram[121][12] ;
   wire \ram[121][11] ;
   wire \ram[121][10] ;
   wire \ram[121][9] ;
   wire \ram[121][8] ;
   wire \ram[121][7] ;
   wire \ram[121][6] ;
   wire \ram[121][5] ;
   wire \ram[121][4] ;
   wire \ram[121][3] ;
   wire \ram[121][2] ;
   wire \ram[121][1] ;
   wire \ram[121][0] ;
   wire \ram[120][15] ;
   wire \ram[120][14] ;
   wire \ram[120][13] ;
   wire \ram[120][12] ;
   wire \ram[120][11] ;
   wire \ram[120][10] ;
   wire \ram[120][9] ;
   wire \ram[120][8] ;
   wire \ram[120][7] ;
   wire \ram[120][6] ;
   wire \ram[120][5] ;
   wire \ram[120][4] ;
   wire \ram[120][3] ;
   wire \ram[120][2] ;
   wire \ram[120][1] ;
   wire \ram[120][0] ;
   wire \ram[119][15] ;
   wire \ram[119][14] ;
   wire \ram[119][13] ;
   wire \ram[119][12] ;
   wire \ram[119][11] ;
   wire \ram[119][10] ;
   wire \ram[119][9] ;
   wire \ram[119][8] ;
   wire \ram[119][7] ;
   wire \ram[119][6] ;
   wire \ram[119][5] ;
   wire \ram[119][4] ;
   wire \ram[119][3] ;
   wire \ram[119][2] ;
   wire \ram[119][1] ;
   wire \ram[119][0] ;
   wire \ram[118][15] ;
   wire \ram[118][14] ;
   wire \ram[118][13] ;
   wire \ram[118][12] ;
   wire \ram[118][11] ;
   wire \ram[118][10] ;
   wire \ram[118][9] ;
   wire \ram[118][8] ;
   wire \ram[118][7] ;
   wire \ram[118][6] ;
   wire \ram[118][5] ;
   wire \ram[118][4] ;
   wire \ram[118][3] ;
   wire \ram[118][2] ;
   wire \ram[118][1] ;
   wire \ram[118][0] ;
   wire \ram[117][15] ;
   wire \ram[117][14] ;
   wire \ram[117][13] ;
   wire \ram[117][12] ;
   wire \ram[117][11] ;
   wire \ram[117][10] ;
   wire \ram[117][9] ;
   wire \ram[117][8] ;
   wire \ram[117][7] ;
   wire \ram[117][6] ;
   wire \ram[117][5] ;
   wire \ram[117][4] ;
   wire \ram[117][3] ;
   wire \ram[117][2] ;
   wire \ram[117][1] ;
   wire \ram[117][0] ;
   wire \ram[116][15] ;
   wire \ram[116][14] ;
   wire \ram[116][13] ;
   wire \ram[116][12] ;
   wire \ram[116][11] ;
   wire \ram[116][10] ;
   wire \ram[116][9] ;
   wire \ram[116][8] ;
   wire \ram[116][7] ;
   wire \ram[116][6] ;
   wire \ram[116][5] ;
   wire \ram[116][4] ;
   wire \ram[116][3] ;
   wire \ram[116][2] ;
   wire \ram[116][1] ;
   wire \ram[116][0] ;
   wire \ram[115][15] ;
   wire \ram[115][14] ;
   wire \ram[115][13] ;
   wire \ram[115][12] ;
   wire \ram[115][11] ;
   wire \ram[115][10] ;
   wire \ram[115][9] ;
   wire \ram[115][8] ;
   wire \ram[115][7] ;
   wire \ram[115][6] ;
   wire \ram[115][5] ;
   wire \ram[115][4] ;
   wire \ram[115][3] ;
   wire \ram[115][2] ;
   wire \ram[115][1] ;
   wire \ram[115][0] ;
   wire \ram[114][15] ;
   wire \ram[114][14] ;
   wire \ram[114][13] ;
   wire \ram[114][12] ;
   wire \ram[114][11] ;
   wire \ram[114][10] ;
   wire \ram[114][9] ;
   wire \ram[114][8] ;
   wire \ram[114][7] ;
   wire \ram[114][6] ;
   wire \ram[114][5] ;
   wire \ram[114][4] ;
   wire \ram[114][3] ;
   wire \ram[114][2] ;
   wire \ram[114][1] ;
   wire \ram[114][0] ;
   wire \ram[113][15] ;
   wire \ram[113][14] ;
   wire \ram[113][13] ;
   wire \ram[113][12] ;
   wire \ram[113][11] ;
   wire \ram[113][10] ;
   wire \ram[113][9] ;
   wire \ram[113][8] ;
   wire \ram[113][7] ;
   wire \ram[113][6] ;
   wire \ram[113][5] ;
   wire \ram[113][4] ;
   wire \ram[113][3] ;
   wire \ram[113][2] ;
   wire \ram[113][1] ;
   wire \ram[113][0] ;
   wire \ram[112][15] ;
   wire \ram[112][14] ;
   wire \ram[112][13] ;
   wire \ram[112][12] ;
   wire \ram[112][11] ;
   wire \ram[112][10] ;
   wire \ram[112][9] ;
   wire \ram[112][8] ;
   wire \ram[112][7] ;
   wire \ram[112][6] ;
   wire \ram[112][5] ;
   wire \ram[112][4] ;
   wire \ram[112][3] ;
   wire \ram[112][2] ;
   wire \ram[112][1] ;
   wire \ram[112][0] ;
   wire \ram[111][15] ;
   wire \ram[111][14] ;
   wire \ram[111][13] ;
   wire \ram[111][12] ;
   wire \ram[111][11] ;
   wire \ram[111][10] ;
   wire \ram[111][9] ;
   wire \ram[111][8] ;
   wire \ram[111][7] ;
   wire \ram[111][6] ;
   wire \ram[111][5] ;
   wire \ram[111][4] ;
   wire \ram[111][3] ;
   wire \ram[111][2] ;
   wire \ram[111][1] ;
   wire \ram[111][0] ;
   wire \ram[110][15] ;
   wire \ram[110][14] ;
   wire \ram[110][13] ;
   wire \ram[110][12] ;
   wire \ram[110][11] ;
   wire \ram[110][10] ;
   wire \ram[110][9] ;
   wire \ram[110][8] ;
   wire \ram[110][7] ;
   wire \ram[110][6] ;
   wire \ram[110][5] ;
   wire \ram[110][4] ;
   wire \ram[110][3] ;
   wire \ram[110][2] ;
   wire \ram[110][1] ;
   wire \ram[110][0] ;
   wire \ram[109][15] ;
   wire \ram[109][14] ;
   wire \ram[109][13] ;
   wire \ram[109][12] ;
   wire \ram[109][11] ;
   wire \ram[109][10] ;
   wire \ram[109][9] ;
   wire \ram[109][8] ;
   wire \ram[109][7] ;
   wire \ram[109][6] ;
   wire \ram[109][5] ;
   wire \ram[109][4] ;
   wire \ram[109][3] ;
   wire \ram[109][2] ;
   wire \ram[109][1] ;
   wire \ram[109][0] ;
   wire \ram[108][15] ;
   wire \ram[108][14] ;
   wire \ram[108][13] ;
   wire \ram[108][12] ;
   wire \ram[108][11] ;
   wire \ram[108][10] ;
   wire \ram[108][9] ;
   wire \ram[108][8] ;
   wire \ram[108][7] ;
   wire \ram[108][6] ;
   wire \ram[108][5] ;
   wire \ram[108][4] ;
   wire \ram[108][3] ;
   wire \ram[108][2] ;
   wire \ram[108][1] ;
   wire \ram[108][0] ;
   wire \ram[107][15] ;
   wire \ram[107][14] ;
   wire \ram[107][13] ;
   wire \ram[107][12] ;
   wire \ram[107][11] ;
   wire \ram[107][10] ;
   wire \ram[107][9] ;
   wire \ram[107][8] ;
   wire \ram[107][7] ;
   wire \ram[107][6] ;
   wire \ram[107][5] ;
   wire \ram[107][4] ;
   wire \ram[107][3] ;
   wire \ram[107][2] ;
   wire \ram[107][1] ;
   wire \ram[107][0] ;
   wire \ram[106][15] ;
   wire \ram[106][14] ;
   wire \ram[106][13] ;
   wire \ram[106][12] ;
   wire \ram[106][11] ;
   wire \ram[106][10] ;
   wire \ram[106][9] ;
   wire \ram[106][8] ;
   wire \ram[106][7] ;
   wire \ram[106][6] ;
   wire \ram[106][5] ;
   wire \ram[106][4] ;
   wire \ram[106][3] ;
   wire \ram[106][2] ;
   wire \ram[106][1] ;
   wire \ram[106][0] ;
   wire \ram[105][15] ;
   wire \ram[105][14] ;
   wire \ram[105][13] ;
   wire \ram[105][12] ;
   wire \ram[105][11] ;
   wire \ram[105][10] ;
   wire \ram[105][9] ;
   wire \ram[105][8] ;
   wire \ram[105][7] ;
   wire \ram[105][6] ;
   wire \ram[105][5] ;
   wire \ram[105][4] ;
   wire \ram[105][3] ;
   wire \ram[105][2] ;
   wire \ram[105][1] ;
   wire \ram[105][0] ;
   wire \ram[104][15] ;
   wire \ram[104][14] ;
   wire \ram[104][13] ;
   wire \ram[104][12] ;
   wire \ram[104][11] ;
   wire \ram[104][10] ;
   wire \ram[104][9] ;
   wire \ram[104][8] ;
   wire \ram[104][7] ;
   wire \ram[104][6] ;
   wire \ram[104][5] ;
   wire \ram[104][4] ;
   wire \ram[104][3] ;
   wire \ram[104][2] ;
   wire \ram[104][1] ;
   wire \ram[104][0] ;
   wire \ram[103][15] ;
   wire \ram[103][14] ;
   wire \ram[103][13] ;
   wire \ram[103][12] ;
   wire \ram[103][11] ;
   wire \ram[103][10] ;
   wire \ram[103][9] ;
   wire \ram[103][8] ;
   wire \ram[103][7] ;
   wire \ram[103][6] ;
   wire \ram[103][5] ;
   wire \ram[103][4] ;
   wire \ram[103][3] ;
   wire \ram[103][2] ;
   wire \ram[103][1] ;
   wire \ram[103][0] ;
   wire \ram[102][15] ;
   wire \ram[102][14] ;
   wire \ram[102][13] ;
   wire \ram[102][12] ;
   wire \ram[102][11] ;
   wire \ram[102][10] ;
   wire \ram[102][9] ;
   wire \ram[102][8] ;
   wire \ram[102][7] ;
   wire \ram[102][6] ;
   wire \ram[102][5] ;
   wire \ram[102][4] ;
   wire \ram[102][3] ;
   wire \ram[102][2] ;
   wire \ram[102][1] ;
   wire \ram[102][0] ;
   wire \ram[101][15] ;
   wire \ram[101][14] ;
   wire \ram[101][13] ;
   wire \ram[101][12] ;
   wire \ram[101][11] ;
   wire \ram[101][10] ;
   wire \ram[101][9] ;
   wire \ram[101][8] ;
   wire \ram[101][7] ;
   wire \ram[101][6] ;
   wire \ram[101][5] ;
   wire \ram[101][4] ;
   wire \ram[101][3] ;
   wire \ram[101][2] ;
   wire \ram[101][1] ;
   wire \ram[101][0] ;
   wire \ram[100][15] ;
   wire \ram[100][14] ;
   wire \ram[100][13] ;
   wire \ram[100][12] ;
   wire \ram[100][11] ;
   wire \ram[100][10] ;
   wire \ram[100][9] ;
   wire \ram[100][8] ;
   wire \ram[100][7] ;
   wire \ram[100][6] ;
   wire \ram[100][5] ;
   wire \ram[100][4] ;
   wire \ram[100][3] ;
   wire \ram[100][2] ;
   wire \ram[100][1] ;
   wire \ram[100][0] ;
   wire \ram[99][15] ;
   wire \ram[99][14] ;
   wire \ram[99][13] ;
   wire \ram[99][12] ;
   wire \ram[99][11] ;
   wire \ram[99][10] ;
   wire \ram[99][9] ;
   wire \ram[99][8] ;
   wire \ram[99][7] ;
   wire \ram[99][6] ;
   wire \ram[99][5] ;
   wire \ram[99][4] ;
   wire \ram[99][3] ;
   wire \ram[99][2] ;
   wire \ram[99][1] ;
   wire \ram[99][0] ;
   wire \ram[98][15] ;
   wire \ram[98][14] ;
   wire \ram[98][13] ;
   wire \ram[98][12] ;
   wire \ram[98][11] ;
   wire \ram[98][10] ;
   wire \ram[98][9] ;
   wire \ram[98][8] ;
   wire \ram[98][7] ;
   wire \ram[98][6] ;
   wire \ram[98][5] ;
   wire \ram[98][4] ;
   wire \ram[98][3] ;
   wire \ram[98][2] ;
   wire \ram[98][1] ;
   wire \ram[98][0] ;
   wire \ram[97][15] ;
   wire \ram[97][14] ;
   wire \ram[97][13] ;
   wire \ram[97][12] ;
   wire \ram[97][11] ;
   wire \ram[97][10] ;
   wire \ram[97][9] ;
   wire \ram[97][8] ;
   wire \ram[97][7] ;
   wire \ram[97][6] ;
   wire \ram[97][5] ;
   wire \ram[97][4] ;
   wire \ram[97][3] ;
   wire \ram[97][2] ;
   wire \ram[97][1] ;
   wire \ram[97][0] ;
   wire \ram[96][15] ;
   wire \ram[96][14] ;
   wire \ram[96][13] ;
   wire \ram[96][12] ;
   wire \ram[96][11] ;
   wire \ram[96][10] ;
   wire \ram[96][9] ;
   wire \ram[96][8] ;
   wire \ram[96][7] ;
   wire \ram[96][6] ;
   wire \ram[96][5] ;
   wire \ram[96][4] ;
   wire \ram[96][3] ;
   wire \ram[96][2] ;
   wire \ram[96][1] ;
   wire \ram[96][0] ;
   wire \ram[95][15] ;
   wire \ram[95][14] ;
   wire \ram[95][13] ;
   wire \ram[95][12] ;
   wire \ram[95][11] ;
   wire \ram[95][10] ;
   wire \ram[95][9] ;
   wire \ram[95][8] ;
   wire \ram[95][7] ;
   wire \ram[95][6] ;
   wire \ram[95][5] ;
   wire \ram[95][4] ;
   wire \ram[95][3] ;
   wire \ram[95][2] ;
   wire \ram[95][1] ;
   wire \ram[95][0] ;
   wire \ram[94][15] ;
   wire \ram[94][14] ;
   wire \ram[94][13] ;
   wire \ram[94][12] ;
   wire \ram[94][11] ;
   wire \ram[94][10] ;
   wire \ram[94][9] ;
   wire \ram[94][8] ;
   wire \ram[94][7] ;
   wire \ram[94][6] ;
   wire \ram[94][5] ;
   wire \ram[94][4] ;
   wire \ram[94][3] ;
   wire \ram[94][2] ;
   wire \ram[94][1] ;
   wire \ram[94][0] ;
   wire \ram[93][15] ;
   wire \ram[93][14] ;
   wire \ram[93][13] ;
   wire \ram[93][12] ;
   wire \ram[93][11] ;
   wire \ram[93][10] ;
   wire \ram[93][9] ;
   wire \ram[93][8] ;
   wire \ram[93][7] ;
   wire \ram[93][6] ;
   wire \ram[93][5] ;
   wire \ram[93][4] ;
   wire \ram[93][3] ;
   wire \ram[93][2] ;
   wire \ram[93][1] ;
   wire \ram[93][0] ;
   wire \ram[92][15] ;
   wire \ram[92][14] ;
   wire \ram[92][13] ;
   wire \ram[92][12] ;
   wire \ram[92][11] ;
   wire \ram[92][10] ;
   wire \ram[92][9] ;
   wire \ram[92][8] ;
   wire \ram[92][7] ;
   wire \ram[92][6] ;
   wire \ram[92][5] ;
   wire \ram[92][4] ;
   wire \ram[92][3] ;
   wire \ram[92][2] ;
   wire \ram[92][1] ;
   wire \ram[92][0] ;
   wire \ram[91][15] ;
   wire \ram[91][14] ;
   wire \ram[91][13] ;
   wire \ram[91][12] ;
   wire \ram[91][11] ;
   wire \ram[91][10] ;
   wire \ram[91][9] ;
   wire \ram[91][8] ;
   wire \ram[91][7] ;
   wire \ram[91][6] ;
   wire \ram[91][5] ;
   wire \ram[91][4] ;
   wire \ram[91][3] ;
   wire \ram[91][2] ;
   wire \ram[91][1] ;
   wire \ram[91][0] ;
   wire \ram[90][15] ;
   wire \ram[90][14] ;
   wire \ram[90][13] ;
   wire \ram[90][12] ;
   wire \ram[90][11] ;
   wire \ram[90][10] ;
   wire \ram[90][9] ;
   wire \ram[90][8] ;
   wire \ram[90][7] ;
   wire \ram[90][6] ;
   wire \ram[90][5] ;
   wire \ram[90][4] ;
   wire \ram[90][3] ;
   wire \ram[90][2] ;
   wire \ram[90][1] ;
   wire \ram[90][0] ;
   wire \ram[89][15] ;
   wire \ram[89][14] ;
   wire \ram[89][13] ;
   wire \ram[89][12] ;
   wire \ram[89][11] ;
   wire \ram[89][10] ;
   wire \ram[89][9] ;
   wire \ram[89][8] ;
   wire \ram[89][7] ;
   wire \ram[89][6] ;
   wire \ram[89][5] ;
   wire \ram[89][4] ;
   wire \ram[89][3] ;
   wire \ram[89][2] ;
   wire \ram[89][1] ;
   wire \ram[89][0] ;
   wire \ram[88][15] ;
   wire \ram[88][14] ;
   wire \ram[88][13] ;
   wire \ram[88][12] ;
   wire \ram[88][11] ;
   wire \ram[88][10] ;
   wire \ram[88][9] ;
   wire \ram[88][8] ;
   wire \ram[88][7] ;
   wire \ram[88][6] ;
   wire \ram[88][5] ;
   wire \ram[88][4] ;
   wire \ram[88][3] ;
   wire \ram[88][2] ;
   wire \ram[88][1] ;
   wire \ram[88][0] ;
   wire \ram[87][15] ;
   wire \ram[87][14] ;
   wire \ram[87][13] ;
   wire \ram[87][12] ;
   wire \ram[87][11] ;
   wire \ram[87][10] ;
   wire \ram[87][9] ;
   wire \ram[87][8] ;
   wire \ram[87][7] ;
   wire \ram[87][6] ;
   wire \ram[87][5] ;
   wire \ram[87][4] ;
   wire \ram[87][3] ;
   wire \ram[87][2] ;
   wire \ram[87][1] ;
   wire \ram[87][0] ;
   wire \ram[86][15] ;
   wire \ram[86][14] ;
   wire \ram[86][13] ;
   wire \ram[86][12] ;
   wire \ram[86][11] ;
   wire \ram[86][10] ;
   wire \ram[86][9] ;
   wire \ram[86][8] ;
   wire \ram[86][7] ;
   wire \ram[86][6] ;
   wire \ram[86][5] ;
   wire \ram[86][4] ;
   wire \ram[86][3] ;
   wire \ram[86][2] ;
   wire \ram[86][1] ;
   wire \ram[86][0] ;
   wire \ram[85][15] ;
   wire \ram[85][14] ;
   wire \ram[85][13] ;
   wire \ram[85][12] ;
   wire \ram[85][11] ;
   wire \ram[85][10] ;
   wire \ram[85][9] ;
   wire \ram[85][8] ;
   wire \ram[85][7] ;
   wire \ram[85][6] ;
   wire \ram[85][5] ;
   wire \ram[85][4] ;
   wire \ram[85][3] ;
   wire \ram[85][2] ;
   wire \ram[85][1] ;
   wire \ram[85][0] ;
   wire \ram[84][15] ;
   wire \ram[84][14] ;
   wire \ram[84][13] ;
   wire \ram[84][12] ;
   wire \ram[84][11] ;
   wire \ram[84][10] ;
   wire \ram[84][9] ;
   wire \ram[84][8] ;
   wire \ram[84][7] ;
   wire \ram[84][6] ;
   wire \ram[84][5] ;
   wire \ram[84][4] ;
   wire \ram[84][3] ;
   wire \ram[84][2] ;
   wire \ram[84][1] ;
   wire \ram[84][0] ;
   wire \ram[83][15] ;
   wire \ram[83][14] ;
   wire \ram[83][13] ;
   wire \ram[83][12] ;
   wire \ram[83][11] ;
   wire \ram[83][10] ;
   wire \ram[83][9] ;
   wire \ram[83][8] ;
   wire \ram[83][7] ;
   wire \ram[83][6] ;
   wire \ram[83][5] ;
   wire \ram[83][4] ;
   wire \ram[83][3] ;
   wire \ram[83][2] ;
   wire \ram[83][1] ;
   wire \ram[83][0] ;
   wire \ram[82][15] ;
   wire \ram[82][14] ;
   wire \ram[82][13] ;
   wire \ram[82][12] ;
   wire \ram[82][11] ;
   wire \ram[82][10] ;
   wire \ram[82][9] ;
   wire \ram[82][8] ;
   wire \ram[82][7] ;
   wire \ram[82][6] ;
   wire \ram[82][5] ;
   wire \ram[82][4] ;
   wire \ram[82][3] ;
   wire \ram[82][2] ;
   wire \ram[82][1] ;
   wire \ram[82][0] ;
   wire \ram[81][15] ;
   wire \ram[81][14] ;
   wire \ram[81][13] ;
   wire \ram[81][12] ;
   wire \ram[81][11] ;
   wire \ram[81][10] ;
   wire \ram[81][9] ;
   wire \ram[81][8] ;
   wire \ram[81][7] ;
   wire \ram[81][6] ;
   wire \ram[81][5] ;
   wire \ram[81][4] ;
   wire \ram[81][3] ;
   wire \ram[81][2] ;
   wire \ram[81][1] ;
   wire \ram[81][0] ;
   wire \ram[80][15] ;
   wire \ram[80][14] ;
   wire \ram[80][13] ;
   wire \ram[80][12] ;
   wire \ram[80][11] ;
   wire \ram[80][10] ;
   wire \ram[80][9] ;
   wire \ram[80][8] ;
   wire \ram[80][7] ;
   wire \ram[80][6] ;
   wire \ram[80][5] ;
   wire \ram[80][4] ;
   wire \ram[80][3] ;
   wire \ram[80][2] ;
   wire \ram[80][1] ;
   wire \ram[80][0] ;
   wire \ram[79][15] ;
   wire \ram[79][14] ;
   wire \ram[79][13] ;
   wire \ram[79][12] ;
   wire \ram[79][11] ;
   wire \ram[79][10] ;
   wire \ram[79][9] ;
   wire \ram[79][8] ;
   wire \ram[79][7] ;
   wire \ram[79][6] ;
   wire \ram[79][5] ;
   wire \ram[79][4] ;
   wire \ram[79][3] ;
   wire \ram[79][2] ;
   wire \ram[79][1] ;
   wire \ram[79][0] ;
   wire \ram[78][15] ;
   wire \ram[78][14] ;
   wire \ram[78][13] ;
   wire \ram[78][12] ;
   wire \ram[78][11] ;
   wire \ram[78][10] ;
   wire \ram[78][9] ;
   wire \ram[78][8] ;
   wire \ram[78][7] ;
   wire \ram[78][6] ;
   wire \ram[78][5] ;
   wire \ram[78][4] ;
   wire \ram[78][3] ;
   wire \ram[78][2] ;
   wire \ram[78][1] ;
   wire \ram[78][0] ;
   wire \ram[77][15] ;
   wire \ram[77][14] ;
   wire \ram[77][13] ;
   wire \ram[77][12] ;
   wire \ram[77][11] ;
   wire \ram[77][10] ;
   wire \ram[77][9] ;
   wire \ram[77][8] ;
   wire \ram[77][7] ;
   wire \ram[77][6] ;
   wire \ram[77][5] ;
   wire \ram[77][4] ;
   wire \ram[77][3] ;
   wire \ram[77][2] ;
   wire \ram[77][1] ;
   wire \ram[77][0] ;
   wire \ram[76][15] ;
   wire \ram[76][14] ;
   wire \ram[76][13] ;
   wire \ram[76][12] ;
   wire \ram[76][11] ;
   wire \ram[76][10] ;
   wire \ram[76][9] ;
   wire \ram[76][8] ;
   wire \ram[76][7] ;
   wire \ram[76][6] ;
   wire \ram[76][5] ;
   wire \ram[76][4] ;
   wire \ram[76][3] ;
   wire \ram[76][2] ;
   wire \ram[76][1] ;
   wire \ram[76][0] ;
   wire \ram[75][15] ;
   wire \ram[75][14] ;
   wire \ram[75][13] ;
   wire \ram[75][12] ;
   wire \ram[75][11] ;
   wire \ram[75][10] ;
   wire \ram[75][9] ;
   wire \ram[75][8] ;
   wire \ram[75][7] ;
   wire \ram[75][6] ;
   wire \ram[75][5] ;
   wire \ram[75][4] ;
   wire \ram[75][3] ;
   wire \ram[75][2] ;
   wire \ram[75][1] ;
   wire \ram[75][0] ;
   wire \ram[74][15] ;
   wire \ram[74][14] ;
   wire \ram[74][13] ;
   wire \ram[74][12] ;
   wire \ram[74][11] ;
   wire \ram[74][10] ;
   wire \ram[74][9] ;
   wire \ram[74][8] ;
   wire \ram[74][7] ;
   wire \ram[74][6] ;
   wire \ram[74][5] ;
   wire \ram[74][4] ;
   wire \ram[74][3] ;
   wire \ram[74][2] ;
   wire \ram[74][1] ;
   wire \ram[74][0] ;
   wire \ram[73][15] ;
   wire \ram[73][14] ;
   wire \ram[73][13] ;
   wire \ram[73][12] ;
   wire \ram[73][11] ;
   wire \ram[73][10] ;
   wire \ram[73][9] ;
   wire \ram[73][8] ;
   wire \ram[73][7] ;
   wire \ram[73][6] ;
   wire \ram[73][5] ;
   wire \ram[73][4] ;
   wire \ram[73][3] ;
   wire \ram[73][2] ;
   wire \ram[73][1] ;
   wire \ram[73][0] ;
   wire \ram[72][15] ;
   wire \ram[72][14] ;
   wire \ram[72][13] ;
   wire \ram[72][12] ;
   wire \ram[72][11] ;
   wire \ram[72][10] ;
   wire \ram[72][9] ;
   wire \ram[72][8] ;
   wire \ram[72][7] ;
   wire \ram[72][6] ;
   wire \ram[72][5] ;
   wire \ram[72][4] ;
   wire \ram[72][3] ;
   wire \ram[72][2] ;
   wire \ram[72][1] ;
   wire \ram[72][0] ;
   wire \ram[71][15] ;
   wire \ram[71][14] ;
   wire \ram[71][13] ;
   wire \ram[71][12] ;
   wire \ram[71][11] ;
   wire \ram[71][10] ;
   wire \ram[71][9] ;
   wire \ram[71][8] ;
   wire \ram[71][7] ;
   wire \ram[71][6] ;
   wire \ram[71][5] ;
   wire \ram[71][4] ;
   wire \ram[71][3] ;
   wire \ram[71][2] ;
   wire \ram[71][1] ;
   wire \ram[71][0] ;
   wire \ram[70][15] ;
   wire \ram[70][14] ;
   wire \ram[70][13] ;
   wire \ram[70][12] ;
   wire \ram[70][11] ;
   wire \ram[70][10] ;
   wire \ram[70][9] ;
   wire \ram[70][8] ;
   wire \ram[70][7] ;
   wire \ram[70][6] ;
   wire \ram[70][5] ;
   wire \ram[70][4] ;
   wire \ram[70][3] ;
   wire \ram[70][2] ;
   wire \ram[70][1] ;
   wire \ram[70][0] ;
   wire \ram[69][15] ;
   wire \ram[69][14] ;
   wire \ram[69][13] ;
   wire \ram[69][12] ;
   wire \ram[69][11] ;
   wire \ram[69][10] ;
   wire \ram[69][9] ;
   wire \ram[69][8] ;
   wire \ram[69][7] ;
   wire \ram[69][6] ;
   wire \ram[69][5] ;
   wire \ram[69][4] ;
   wire \ram[69][3] ;
   wire \ram[69][2] ;
   wire \ram[69][1] ;
   wire \ram[69][0] ;
   wire \ram[68][15] ;
   wire \ram[68][14] ;
   wire \ram[68][13] ;
   wire \ram[68][12] ;
   wire \ram[68][11] ;
   wire \ram[68][10] ;
   wire \ram[68][9] ;
   wire \ram[68][8] ;
   wire \ram[68][7] ;
   wire \ram[68][6] ;
   wire \ram[68][5] ;
   wire \ram[68][4] ;
   wire \ram[68][3] ;
   wire \ram[68][2] ;
   wire \ram[68][1] ;
   wire \ram[68][0] ;
   wire \ram[67][15] ;
   wire \ram[67][14] ;
   wire \ram[67][13] ;
   wire \ram[67][12] ;
   wire \ram[67][11] ;
   wire \ram[67][10] ;
   wire \ram[67][9] ;
   wire \ram[67][8] ;
   wire \ram[67][7] ;
   wire \ram[67][6] ;
   wire \ram[67][5] ;
   wire \ram[67][4] ;
   wire \ram[67][3] ;
   wire \ram[67][2] ;
   wire \ram[67][1] ;
   wire \ram[67][0] ;
   wire \ram[66][15] ;
   wire \ram[66][14] ;
   wire \ram[66][13] ;
   wire \ram[66][12] ;
   wire \ram[66][11] ;
   wire \ram[66][10] ;
   wire \ram[66][9] ;
   wire \ram[66][8] ;
   wire \ram[66][7] ;
   wire \ram[66][6] ;
   wire \ram[66][5] ;
   wire \ram[66][4] ;
   wire \ram[66][3] ;
   wire \ram[66][2] ;
   wire \ram[66][1] ;
   wire \ram[66][0] ;
   wire \ram[65][15] ;
   wire \ram[65][14] ;
   wire \ram[65][13] ;
   wire \ram[65][12] ;
   wire \ram[65][11] ;
   wire \ram[65][10] ;
   wire \ram[65][9] ;
   wire \ram[65][8] ;
   wire \ram[65][7] ;
   wire \ram[65][6] ;
   wire \ram[65][5] ;
   wire \ram[65][4] ;
   wire \ram[65][3] ;
   wire \ram[65][2] ;
   wire \ram[65][1] ;
   wire \ram[65][0] ;
   wire \ram[64][15] ;
   wire \ram[64][14] ;
   wire \ram[64][13] ;
   wire \ram[64][12] ;
   wire \ram[64][11] ;
   wire \ram[64][10] ;
   wire \ram[64][9] ;
   wire \ram[64][8] ;
   wire \ram[64][7] ;
   wire \ram[64][6] ;
   wire \ram[64][5] ;
   wire \ram[64][4] ;
   wire \ram[64][3] ;
   wire \ram[64][2] ;
   wire \ram[64][1] ;
   wire \ram[64][0] ;
   wire \ram[63][15] ;
   wire \ram[63][14] ;
   wire \ram[63][13] ;
   wire \ram[63][12] ;
   wire \ram[63][11] ;
   wire \ram[63][10] ;
   wire \ram[63][9] ;
   wire \ram[63][8] ;
   wire \ram[63][7] ;
   wire \ram[63][6] ;
   wire \ram[63][5] ;
   wire \ram[63][4] ;
   wire \ram[63][3] ;
   wire \ram[63][2] ;
   wire \ram[63][1] ;
   wire \ram[63][0] ;
   wire \ram[62][15] ;
   wire \ram[62][14] ;
   wire \ram[62][13] ;
   wire \ram[62][12] ;
   wire \ram[62][11] ;
   wire \ram[62][10] ;
   wire \ram[62][9] ;
   wire \ram[62][8] ;
   wire \ram[62][7] ;
   wire \ram[62][6] ;
   wire \ram[62][5] ;
   wire \ram[62][4] ;
   wire \ram[62][3] ;
   wire \ram[62][2] ;
   wire \ram[62][1] ;
   wire \ram[62][0] ;
   wire \ram[61][15] ;
   wire \ram[61][14] ;
   wire \ram[61][13] ;
   wire \ram[61][12] ;
   wire \ram[61][11] ;
   wire \ram[61][10] ;
   wire \ram[61][9] ;
   wire \ram[61][8] ;
   wire \ram[61][7] ;
   wire \ram[61][6] ;
   wire \ram[61][5] ;
   wire \ram[61][4] ;
   wire \ram[61][3] ;
   wire \ram[61][2] ;
   wire \ram[61][1] ;
   wire \ram[61][0] ;
   wire \ram[60][15] ;
   wire \ram[60][14] ;
   wire \ram[60][13] ;
   wire \ram[60][12] ;
   wire \ram[60][11] ;
   wire \ram[60][10] ;
   wire \ram[60][9] ;
   wire \ram[60][8] ;
   wire \ram[60][7] ;
   wire \ram[60][6] ;
   wire \ram[60][5] ;
   wire \ram[60][4] ;
   wire \ram[60][3] ;
   wire \ram[60][2] ;
   wire \ram[60][1] ;
   wire \ram[60][0] ;
   wire \ram[59][15] ;
   wire \ram[59][14] ;
   wire \ram[59][13] ;
   wire \ram[59][12] ;
   wire \ram[59][11] ;
   wire \ram[59][10] ;
   wire \ram[59][9] ;
   wire \ram[59][8] ;
   wire \ram[59][7] ;
   wire \ram[59][6] ;
   wire \ram[59][5] ;
   wire \ram[59][4] ;
   wire \ram[59][3] ;
   wire \ram[59][2] ;
   wire \ram[59][1] ;
   wire \ram[59][0] ;
   wire \ram[58][15] ;
   wire \ram[58][14] ;
   wire \ram[58][13] ;
   wire \ram[58][12] ;
   wire \ram[58][11] ;
   wire \ram[58][10] ;
   wire \ram[58][9] ;
   wire \ram[58][8] ;
   wire \ram[58][7] ;
   wire \ram[58][6] ;
   wire \ram[58][5] ;
   wire \ram[58][4] ;
   wire \ram[58][3] ;
   wire \ram[58][2] ;
   wire \ram[58][1] ;
   wire \ram[58][0] ;
   wire \ram[57][15] ;
   wire \ram[57][14] ;
   wire \ram[57][13] ;
   wire \ram[57][12] ;
   wire \ram[57][11] ;
   wire \ram[57][10] ;
   wire \ram[57][9] ;
   wire \ram[57][8] ;
   wire \ram[57][7] ;
   wire \ram[57][6] ;
   wire \ram[57][5] ;
   wire \ram[57][4] ;
   wire \ram[57][3] ;
   wire \ram[57][2] ;
   wire \ram[57][1] ;
   wire \ram[57][0] ;
   wire \ram[56][15] ;
   wire \ram[56][14] ;
   wire \ram[56][13] ;
   wire \ram[56][12] ;
   wire \ram[56][11] ;
   wire \ram[56][10] ;
   wire \ram[56][9] ;
   wire \ram[56][8] ;
   wire \ram[56][7] ;
   wire \ram[56][6] ;
   wire \ram[56][5] ;
   wire \ram[56][4] ;
   wire \ram[56][3] ;
   wire \ram[56][2] ;
   wire \ram[56][1] ;
   wire \ram[56][0] ;
   wire \ram[55][15] ;
   wire \ram[55][14] ;
   wire \ram[55][13] ;
   wire \ram[55][12] ;
   wire \ram[55][11] ;
   wire \ram[55][10] ;
   wire \ram[55][9] ;
   wire \ram[55][8] ;
   wire \ram[55][7] ;
   wire \ram[55][6] ;
   wire \ram[55][5] ;
   wire \ram[55][4] ;
   wire \ram[55][3] ;
   wire \ram[55][2] ;
   wire \ram[55][1] ;
   wire \ram[55][0] ;
   wire \ram[54][15] ;
   wire \ram[54][14] ;
   wire \ram[54][13] ;
   wire \ram[54][12] ;
   wire \ram[54][11] ;
   wire \ram[54][10] ;
   wire \ram[54][9] ;
   wire \ram[54][8] ;
   wire \ram[54][7] ;
   wire \ram[54][6] ;
   wire \ram[54][5] ;
   wire \ram[54][4] ;
   wire \ram[54][3] ;
   wire \ram[54][2] ;
   wire \ram[54][1] ;
   wire \ram[54][0] ;
   wire \ram[53][15] ;
   wire \ram[53][14] ;
   wire \ram[53][13] ;
   wire \ram[53][12] ;
   wire \ram[53][11] ;
   wire \ram[53][10] ;
   wire \ram[53][9] ;
   wire \ram[53][8] ;
   wire \ram[53][7] ;
   wire \ram[53][6] ;
   wire \ram[53][5] ;
   wire \ram[53][4] ;
   wire \ram[53][3] ;
   wire \ram[53][2] ;
   wire \ram[53][1] ;
   wire \ram[53][0] ;
   wire \ram[52][15] ;
   wire \ram[52][14] ;
   wire \ram[52][13] ;
   wire \ram[52][12] ;
   wire \ram[52][11] ;
   wire \ram[52][10] ;
   wire \ram[52][9] ;
   wire \ram[52][8] ;
   wire \ram[52][7] ;
   wire \ram[52][6] ;
   wire \ram[52][5] ;
   wire \ram[52][4] ;
   wire \ram[52][3] ;
   wire \ram[52][2] ;
   wire \ram[52][1] ;
   wire \ram[52][0] ;
   wire \ram[51][15] ;
   wire \ram[51][14] ;
   wire \ram[51][13] ;
   wire \ram[51][12] ;
   wire \ram[51][11] ;
   wire \ram[51][10] ;
   wire \ram[51][9] ;
   wire \ram[51][8] ;
   wire \ram[51][7] ;
   wire \ram[51][6] ;
   wire \ram[51][5] ;
   wire \ram[51][4] ;
   wire \ram[51][3] ;
   wire \ram[51][2] ;
   wire \ram[51][1] ;
   wire \ram[51][0] ;
   wire \ram[50][15] ;
   wire \ram[50][14] ;
   wire \ram[50][13] ;
   wire \ram[50][12] ;
   wire \ram[50][11] ;
   wire \ram[50][10] ;
   wire \ram[50][9] ;
   wire \ram[50][8] ;
   wire \ram[50][7] ;
   wire \ram[50][6] ;
   wire \ram[50][5] ;
   wire \ram[50][4] ;
   wire \ram[50][3] ;
   wire \ram[50][2] ;
   wire \ram[50][1] ;
   wire \ram[50][0] ;
   wire \ram[49][15] ;
   wire \ram[49][14] ;
   wire \ram[49][13] ;
   wire \ram[49][12] ;
   wire \ram[49][11] ;
   wire \ram[49][10] ;
   wire \ram[49][9] ;
   wire \ram[49][8] ;
   wire \ram[49][7] ;
   wire \ram[49][6] ;
   wire \ram[49][5] ;
   wire \ram[49][4] ;
   wire \ram[49][3] ;
   wire \ram[49][2] ;
   wire \ram[49][1] ;
   wire \ram[49][0] ;
   wire \ram[48][15] ;
   wire \ram[48][14] ;
   wire \ram[48][13] ;
   wire \ram[48][12] ;
   wire \ram[48][11] ;
   wire \ram[48][10] ;
   wire \ram[48][9] ;
   wire \ram[48][8] ;
   wire \ram[48][7] ;
   wire \ram[48][6] ;
   wire \ram[48][5] ;
   wire \ram[48][4] ;
   wire \ram[48][3] ;
   wire \ram[48][2] ;
   wire \ram[48][1] ;
   wire \ram[48][0] ;
   wire \ram[47][15] ;
   wire \ram[47][14] ;
   wire \ram[47][13] ;
   wire \ram[47][12] ;
   wire \ram[47][11] ;
   wire \ram[47][10] ;
   wire \ram[47][9] ;
   wire \ram[47][8] ;
   wire \ram[47][7] ;
   wire \ram[47][6] ;
   wire \ram[47][5] ;
   wire \ram[47][4] ;
   wire \ram[47][3] ;
   wire \ram[47][2] ;
   wire \ram[47][1] ;
   wire \ram[47][0] ;
   wire \ram[46][15] ;
   wire \ram[46][14] ;
   wire \ram[46][13] ;
   wire \ram[46][12] ;
   wire \ram[46][11] ;
   wire \ram[46][10] ;
   wire \ram[46][9] ;
   wire \ram[46][8] ;
   wire \ram[46][7] ;
   wire \ram[46][6] ;
   wire \ram[46][5] ;
   wire \ram[46][4] ;
   wire \ram[46][3] ;
   wire \ram[46][2] ;
   wire \ram[46][1] ;
   wire \ram[46][0] ;
   wire \ram[45][15] ;
   wire \ram[45][14] ;
   wire \ram[45][13] ;
   wire \ram[45][12] ;
   wire \ram[45][11] ;
   wire \ram[45][10] ;
   wire \ram[45][9] ;
   wire \ram[45][8] ;
   wire \ram[45][7] ;
   wire \ram[45][6] ;
   wire \ram[45][5] ;
   wire \ram[45][4] ;
   wire \ram[45][3] ;
   wire \ram[45][2] ;
   wire \ram[45][1] ;
   wire \ram[45][0] ;
   wire \ram[44][15] ;
   wire \ram[44][14] ;
   wire \ram[44][13] ;
   wire \ram[44][12] ;
   wire \ram[44][11] ;
   wire \ram[44][10] ;
   wire \ram[44][9] ;
   wire \ram[44][8] ;
   wire \ram[44][7] ;
   wire \ram[44][6] ;
   wire \ram[44][5] ;
   wire \ram[44][4] ;
   wire \ram[44][3] ;
   wire \ram[44][2] ;
   wire \ram[44][1] ;
   wire \ram[44][0] ;
   wire \ram[43][15] ;
   wire \ram[43][14] ;
   wire \ram[43][13] ;
   wire \ram[43][12] ;
   wire \ram[43][11] ;
   wire \ram[43][10] ;
   wire \ram[43][9] ;
   wire \ram[43][8] ;
   wire \ram[43][7] ;
   wire \ram[43][6] ;
   wire \ram[43][5] ;
   wire \ram[43][4] ;
   wire \ram[43][3] ;
   wire \ram[43][2] ;
   wire \ram[43][1] ;
   wire \ram[43][0] ;
   wire \ram[42][15] ;
   wire \ram[42][14] ;
   wire \ram[42][13] ;
   wire \ram[42][12] ;
   wire \ram[42][11] ;
   wire \ram[42][10] ;
   wire \ram[42][9] ;
   wire \ram[42][8] ;
   wire \ram[42][7] ;
   wire \ram[42][6] ;
   wire \ram[42][5] ;
   wire \ram[42][4] ;
   wire \ram[42][3] ;
   wire \ram[42][2] ;
   wire \ram[42][1] ;
   wire \ram[42][0] ;
   wire \ram[41][15] ;
   wire \ram[41][14] ;
   wire \ram[41][13] ;
   wire \ram[41][12] ;
   wire \ram[41][11] ;
   wire \ram[41][10] ;
   wire \ram[41][9] ;
   wire \ram[41][8] ;
   wire \ram[41][7] ;
   wire \ram[41][6] ;
   wire \ram[41][5] ;
   wire \ram[41][4] ;
   wire \ram[41][3] ;
   wire \ram[41][2] ;
   wire \ram[41][1] ;
   wire \ram[41][0] ;
   wire \ram[40][15] ;
   wire \ram[40][14] ;
   wire \ram[40][13] ;
   wire \ram[40][12] ;
   wire \ram[40][11] ;
   wire \ram[40][10] ;
   wire \ram[40][9] ;
   wire \ram[40][8] ;
   wire \ram[40][7] ;
   wire \ram[40][6] ;
   wire \ram[40][5] ;
   wire \ram[40][4] ;
   wire \ram[40][3] ;
   wire \ram[40][2] ;
   wire \ram[40][1] ;
   wire \ram[40][0] ;
   wire \ram[39][15] ;
   wire \ram[39][14] ;
   wire \ram[39][13] ;
   wire \ram[39][12] ;
   wire \ram[39][11] ;
   wire \ram[39][10] ;
   wire \ram[39][9] ;
   wire \ram[39][8] ;
   wire \ram[39][7] ;
   wire \ram[39][6] ;
   wire \ram[39][5] ;
   wire \ram[39][4] ;
   wire \ram[39][3] ;
   wire \ram[39][2] ;
   wire \ram[39][1] ;
   wire \ram[39][0] ;
   wire \ram[38][15] ;
   wire \ram[38][14] ;
   wire \ram[38][13] ;
   wire \ram[38][12] ;
   wire \ram[38][11] ;
   wire \ram[38][10] ;
   wire \ram[38][9] ;
   wire \ram[38][8] ;
   wire \ram[38][7] ;
   wire \ram[38][6] ;
   wire \ram[38][5] ;
   wire \ram[38][4] ;
   wire \ram[38][3] ;
   wire \ram[38][2] ;
   wire \ram[38][1] ;
   wire \ram[38][0] ;
   wire \ram[37][15] ;
   wire \ram[37][14] ;
   wire \ram[37][13] ;
   wire \ram[37][12] ;
   wire \ram[37][11] ;
   wire \ram[37][10] ;
   wire \ram[37][9] ;
   wire \ram[37][8] ;
   wire \ram[37][7] ;
   wire \ram[37][6] ;
   wire \ram[37][5] ;
   wire \ram[37][4] ;
   wire \ram[37][3] ;
   wire \ram[37][2] ;
   wire \ram[37][1] ;
   wire \ram[37][0] ;
   wire \ram[36][15] ;
   wire \ram[36][14] ;
   wire \ram[36][13] ;
   wire \ram[36][12] ;
   wire \ram[36][11] ;
   wire \ram[36][10] ;
   wire \ram[36][9] ;
   wire \ram[36][8] ;
   wire \ram[36][7] ;
   wire \ram[36][6] ;
   wire \ram[36][5] ;
   wire \ram[36][4] ;
   wire \ram[36][3] ;
   wire \ram[36][2] ;
   wire \ram[36][1] ;
   wire \ram[36][0] ;
   wire \ram[35][15] ;
   wire \ram[35][14] ;
   wire \ram[35][13] ;
   wire \ram[35][12] ;
   wire \ram[35][11] ;
   wire \ram[35][10] ;
   wire \ram[35][9] ;
   wire \ram[35][8] ;
   wire \ram[35][7] ;
   wire \ram[35][6] ;
   wire \ram[35][5] ;
   wire \ram[35][4] ;
   wire \ram[35][3] ;
   wire \ram[35][2] ;
   wire \ram[35][1] ;
   wire \ram[35][0] ;
   wire \ram[34][15] ;
   wire \ram[34][14] ;
   wire \ram[34][13] ;
   wire \ram[34][12] ;
   wire \ram[34][11] ;
   wire \ram[34][10] ;
   wire \ram[34][9] ;
   wire \ram[34][8] ;
   wire \ram[34][7] ;
   wire \ram[34][6] ;
   wire \ram[34][5] ;
   wire \ram[34][4] ;
   wire \ram[34][3] ;
   wire \ram[34][2] ;
   wire \ram[34][1] ;
   wire \ram[34][0] ;
   wire \ram[33][15] ;
   wire \ram[33][14] ;
   wire \ram[33][13] ;
   wire \ram[33][12] ;
   wire \ram[33][11] ;
   wire \ram[33][10] ;
   wire \ram[33][9] ;
   wire \ram[33][8] ;
   wire \ram[33][7] ;
   wire \ram[33][6] ;
   wire \ram[33][5] ;
   wire \ram[33][4] ;
   wire \ram[33][3] ;
   wire \ram[33][2] ;
   wire \ram[33][1] ;
   wire \ram[33][0] ;
   wire \ram[32][15] ;
   wire \ram[32][14] ;
   wire \ram[32][13] ;
   wire \ram[32][12] ;
   wire \ram[32][11] ;
   wire \ram[32][10] ;
   wire \ram[32][9] ;
   wire \ram[32][8] ;
   wire \ram[32][7] ;
   wire \ram[32][6] ;
   wire \ram[32][5] ;
   wire \ram[32][4] ;
   wire \ram[32][3] ;
   wire \ram[32][2] ;
   wire \ram[32][1] ;
   wire \ram[32][0] ;
   wire \ram[31][15] ;
   wire \ram[31][14] ;
   wire \ram[31][13] ;
   wire \ram[31][12] ;
   wire \ram[31][11] ;
   wire \ram[31][10] ;
   wire \ram[31][9] ;
   wire \ram[31][8] ;
   wire \ram[31][7] ;
   wire \ram[31][6] ;
   wire \ram[31][5] ;
   wire \ram[31][4] ;
   wire \ram[31][3] ;
   wire \ram[31][2] ;
   wire \ram[31][1] ;
   wire \ram[31][0] ;
   wire \ram[30][15] ;
   wire \ram[30][14] ;
   wire \ram[30][13] ;
   wire \ram[30][12] ;
   wire \ram[30][11] ;
   wire \ram[30][10] ;
   wire \ram[30][9] ;
   wire \ram[30][8] ;
   wire \ram[30][7] ;
   wire \ram[30][6] ;
   wire \ram[30][5] ;
   wire \ram[30][4] ;
   wire \ram[30][3] ;
   wire \ram[30][2] ;
   wire \ram[30][1] ;
   wire \ram[30][0] ;
   wire \ram[29][15] ;
   wire \ram[29][14] ;
   wire \ram[29][13] ;
   wire \ram[29][12] ;
   wire \ram[29][11] ;
   wire \ram[29][10] ;
   wire \ram[29][9] ;
   wire \ram[29][8] ;
   wire \ram[29][7] ;
   wire \ram[29][6] ;
   wire \ram[29][5] ;
   wire \ram[29][4] ;
   wire \ram[29][3] ;
   wire \ram[29][2] ;
   wire \ram[29][1] ;
   wire \ram[29][0] ;
   wire \ram[28][15] ;
   wire \ram[28][14] ;
   wire \ram[28][13] ;
   wire \ram[28][12] ;
   wire \ram[28][11] ;
   wire \ram[28][10] ;
   wire \ram[28][9] ;
   wire \ram[28][8] ;
   wire \ram[28][7] ;
   wire \ram[28][6] ;
   wire \ram[28][5] ;
   wire \ram[28][4] ;
   wire \ram[28][3] ;
   wire \ram[28][2] ;
   wire \ram[28][1] ;
   wire \ram[28][0] ;
   wire \ram[27][15] ;
   wire \ram[27][14] ;
   wire \ram[27][13] ;
   wire \ram[27][12] ;
   wire \ram[27][11] ;
   wire \ram[27][10] ;
   wire \ram[27][9] ;
   wire \ram[27][8] ;
   wire \ram[27][7] ;
   wire \ram[27][6] ;
   wire \ram[27][5] ;
   wire \ram[27][4] ;
   wire \ram[27][3] ;
   wire \ram[27][2] ;
   wire \ram[27][1] ;
   wire \ram[27][0] ;
   wire \ram[26][15] ;
   wire \ram[26][14] ;
   wire \ram[26][13] ;
   wire \ram[26][12] ;
   wire \ram[26][11] ;
   wire \ram[26][10] ;
   wire \ram[26][9] ;
   wire \ram[26][8] ;
   wire \ram[26][7] ;
   wire \ram[26][6] ;
   wire \ram[26][5] ;
   wire \ram[26][4] ;
   wire \ram[26][3] ;
   wire \ram[26][2] ;
   wire \ram[26][1] ;
   wire \ram[26][0] ;
   wire \ram[25][15] ;
   wire \ram[25][14] ;
   wire \ram[25][13] ;
   wire \ram[25][12] ;
   wire \ram[25][11] ;
   wire \ram[25][10] ;
   wire \ram[25][9] ;
   wire \ram[25][8] ;
   wire \ram[25][7] ;
   wire \ram[25][6] ;
   wire \ram[25][5] ;
   wire \ram[25][4] ;
   wire \ram[25][3] ;
   wire \ram[25][2] ;
   wire \ram[25][1] ;
   wire \ram[25][0] ;
   wire \ram[24][15] ;
   wire \ram[24][14] ;
   wire \ram[24][13] ;
   wire \ram[24][12] ;
   wire \ram[24][11] ;
   wire \ram[24][10] ;
   wire \ram[24][9] ;
   wire \ram[24][8] ;
   wire \ram[24][7] ;
   wire \ram[24][6] ;
   wire \ram[24][5] ;
   wire \ram[24][4] ;
   wire \ram[24][3] ;
   wire \ram[24][2] ;
   wire \ram[24][1] ;
   wire \ram[24][0] ;
   wire \ram[23][15] ;
   wire \ram[23][14] ;
   wire \ram[23][13] ;
   wire \ram[23][12] ;
   wire \ram[23][11] ;
   wire \ram[23][10] ;
   wire \ram[23][9] ;
   wire \ram[23][8] ;
   wire \ram[23][7] ;
   wire \ram[23][6] ;
   wire \ram[23][5] ;
   wire \ram[23][4] ;
   wire \ram[23][3] ;
   wire \ram[23][2] ;
   wire \ram[23][1] ;
   wire \ram[23][0] ;
   wire \ram[22][15] ;
   wire \ram[22][14] ;
   wire \ram[22][13] ;
   wire \ram[22][12] ;
   wire \ram[22][11] ;
   wire \ram[22][10] ;
   wire \ram[22][9] ;
   wire \ram[22][8] ;
   wire \ram[22][7] ;
   wire \ram[22][6] ;
   wire \ram[22][5] ;
   wire \ram[22][4] ;
   wire \ram[22][3] ;
   wire \ram[22][2] ;
   wire \ram[22][1] ;
   wire \ram[22][0] ;
   wire \ram[21][15] ;
   wire \ram[21][14] ;
   wire \ram[21][13] ;
   wire \ram[21][12] ;
   wire \ram[21][11] ;
   wire \ram[21][10] ;
   wire \ram[21][9] ;
   wire \ram[21][8] ;
   wire \ram[21][7] ;
   wire \ram[21][6] ;
   wire \ram[21][5] ;
   wire \ram[21][4] ;
   wire \ram[21][3] ;
   wire \ram[21][2] ;
   wire \ram[21][1] ;
   wire \ram[21][0] ;
   wire \ram[20][15] ;
   wire \ram[20][14] ;
   wire \ram[20][13] ;
   wire \ram[20][12] ;
   wire \ram[20][11] ;
   wire \ram[20][10] ;
   wire \ram[20][9] ;
   wire \ram[20][8] ;
   wire \ram[20][7] ;
   wire \ram[20][6] ;
   wire \ram[20][5] ;
   wire \ram[20][4] ;
   wire \ram[20][3] ;
   wire \ram[20][2] ;
   wire \ram[20][1] ;
   wire \ram[20][0] ;
   wire \ram[19][15] ;
   wire \ram[19][14] ;
   wire \ram[19][13] ;
   wire \ram[19][12] ;
   wire \ram[19][11] ;
   wire \ram[19][10] ;
   wire \ram[19][9] ;
   wire \ram[19][8] ;
   wire \ram[19][7] ;
   wire \ram[19][6] ;
   wire \ram[19][5] ;
   wire \ram[19][4] ;
   wire \ram[19][3] ;
   wire \ram[19][2] ;
   wire \ram[19][1] ;
   wire \ram[19][0] ;
   wire \ram[18][15] ;
   wire \ram[18][14] ;
   wire \ram[18][13] ;
   wire \ram[18][12] ;
   wire \ram[18][11] ;
   wire \ram[18][10] ;
   wire \ram[18][9] ;
   wire \ram[18][8] ;
   wire \ram[18][7] ;
   wire \ram[18][6] ;
   wire \ram[18][5] ;
   wire \ram[18][4] ;
   wire \ram[18][3] ;
   wire \ram[18][2] ;
   wire \ram[18][1] ;
   wire \ram[18][0] ;
   wire \ram[17][15] ;
   wire \ram[17][14] ;
   wire \ram[17][13] ;
   wire \ram[17][12] ;
   wire \ram[17][11] ;
   wire \ram[17][10] ;
   wire \ram[17][9] ;
   wire \ram[17][8] ;
   wire \ram[17][7] ;
   wire \ram[17][6] ;
   wire \ram[17][5] ;
   wire \ram[17][4] ;
   wire \ram[17][3] ;
   wire \ram[17][2] ;
   wire \ram[17][1] ;
   wire \ram[17][0] ;
   wire \ram[16][15] ;
   wire \ram[16][14] ;
   wire \ram[16][13] ;
   wire \ram[16][12] ;
   wire \ram[16][11] ;
   wire \ram[16][10] ;
   wire \ram[16][9] ;
   wire \ram[16][8] ;
   wire \ram[16][7] ;
   wire \ram[16][6] ;
   wire \ram[16][5] ;
   wire \ram[16][4] ;
   wire \ram[16][3] ;
   wire \ram[16][2] ;
   wire \ram[16][1] ;
   wire \ram[16][0] ;
   wire \ram[15][15] ;
   wire \ram[15][14] ;
   wire \ram[15][13] ;
   wire \ram[15][12] ;
   wire \ram[15][11] ;
   wire \ram[15][10] ;
   wire \ram[15][9] ;
   wire \ram[15][8] ;
   wire \ram[15][7] ;
   wire \ram[15][6] ;
   wire \ram[15][5] ;
   wire \ram[15][4] ;
   wire \ram[15][3] ;
   wire \ram[15][2] ;
   wire \ram[15][1] ;
   wire \ram[15][0] ;
   wire \ram[14][15] ;
   wire \ram[14][14] ;
   wire \ram[14][13] ;
   wire \ram[14][12] ;
   wire \ram[14][11] ;
   wire \ram[14][10] ;
   wire \ram[14][9] ;
   wire \ram[14][8] ;
   wire \ram[14][7] ;
   wire \ram[14][6] ;
   wire \ram[14][5] ;
   wire \ram[14][4] ;
   wire \ram[14][3] ;
   wire \ram[14][2] ;
   wire \ram[14][1] ;
   wire \ram[14][0] ;
   wire \ram[13][15] ;
   wire \ram[13][14] ;
   wire \ram[13][13] ;
   wire \ram[13][12] ;
   wire \ram[13][11] ;
   wire \ram[13][10] ;
   wire \ram[13][9] ;
   wire \ram[13][8] ;
   wire \ram[13][7] ;
   wire \ram[13][6] ;
   wire \ram[13][5] ;
   wire \ram[13][4] ;
   wire \ram[13][3] ;
   wire \ram[13][2] ;
   wire \ram[13][1] ;
   wire \ram[13][0] ;
   wire \ram[12][15] ;
   wire \ram[12][14] ;
   wire \ram[12][13] ;
   wire \ram[12][12] ;
   wire \ram[12][11] ;
   wire \ram[12][10] ;
   wire \ram[12][9] ;
   wire \ram[12][8] ;
   wire \ram[12][7] ;
   wire \ram[12][6] ;
   wire \ram[12][5] ;
   wire \ram[12][4] ;
   wire \ram[12][3] ;
   wire \ram[12][2] ;
   wire \ram[12][1] ;
   wire \ram[12][0] ;
   wire \ram[11][15] ;
   wire \ram[11][14] ;
   wire \ram[11][13] ;
   wire \ram[11][12] ;
   wire \ram[11][11] ;
   wire \ram[11][10] ;
   wire \ram[11][9] ;
   wire \ram[11][8] ;
   wire \ram[11][7] ;
   wire \ram[11][6] ;
   wire \ram[11][5] ;
   wire \ram[11][4] ;
   wire \ram[11][3] ;
   wire \ram[11][2] ;
   wire \ram[11][1] ;
   wire \ram[11][0] ;
   wire \ram[10][15] ;
   wire \ram[10][14] ;
   wire \ram[10][13] ;
   wire \ram[10][12] ;
   wire \ram[10][11] ;
   wire \ram[10][10] ;
   wire \ram[10][9] ;
   wire \ram[10][8] ;
   wire \ram[10][7] ;
   wire \ram[10][6] ;
   wire \ram[10][5] ;
   wire \ram[10][4] ;
   wire \ram[10][3] ;
   wire \ram[10][2] ;
   wire \ram[10][1] ;
   wire \ram[10][0] ;
   wire \ram[9][15] ;
   wire \ram[9][14] ;
   wire \ram[9][13] ;
   wire \ram[9][12] ;
   wire \ram[9][11] ;
   wire \ram[9][10] ;
   wire \ram[9][9] ;
   wire \ram[9][8] ;
   wire \ram[9][7] ;
   wire \ram[9][6] ;
   wire \ram[9][5] ;
   wire \ram[9][4] ;
   wire \ram[9][3] ;
   wire \ram[9][2] ;
   wire \ram[9][1] ;
   wire \ram[9][0] ;
   wire \ram[8][15] ;
   wire \ram[8][14] ;
   wire \ram[8][13] ;
   wire \ram[8][12] ;
   wire \ram[8][11] ;
   wire \ram[8][10] ;
   wire \ram[8][9] ;
   wire \ram[8][8] ;
   wire \ram[8][7] ;
   wire \ram[8][6] ;
   wire \ram[8][5] ;
   wire \ram[8][4] ;
   wire \ram[8][3] ;
   wire \ram[8][2] ;
   wire \ram[8][1] ;
   wire \ram[8][0] ;
   wire \ram[7][15] ;
   wire \ram[7][14] ;
   wire \ram[7][13] ;
   wire \ram[7][12] ;
   wire \ram[7][11] ;
   wire \ram[7][10] ;
   wire \ram[7][9] ;
   wire \ram[7][8] ;
   wire \ram[7][7] ;
   wire \ram[7][6] ;
   wire \ram[7][5] ;
   wire \ram[7][4] ;
   wire \ram[7][3] ;
   wire \ram[7][2] ;
   wire \ram[7][1] ;
   wire \ram[7][0] ;
   wire \ram[6][15] ;
   wire \ram[6][14] ;
   wire \ram[6][13] ;
   wire \ram[6][12] ;
   wire \ram[6][11] ;
   wire \ram[6][10] ;
   wire \ram[6][9] ;
   wire \ram[6][8] ;
   wire \ram[6][7] ;
   wire \ram[6][6] ;
   wire \ram[6][5] ;
   wire \ram[6][4] ;
   wire \ram[6][3] ;
   wire \ram[6][2] ;
   wire \ram[6][1] ;
   wire \ram[6][0] ;
   wire \ram[5][15] ;
   wire \ram[5][14] ;
   wire \ram[5][13] ;
   wire \ram[5][12] ;
   wire \ram[5][11] ;
   wire \ram[5][10] ;
   wire \ram[5][9] ;
   wire \ram[5][8] ;
   wire \ram[5][7] ;
   wire \ram[5][6] ;
   wire \ram[5][5] ;
   wire \ram[5][4] ;
   wire \ram[5][3] ;
   wire \ram[5][2] ;
   wire \ram[5][1] ;
   wire \ram[5][0] ;
   wire \ram[4][15] ;
   wire \ram[4][14] ;
   wire \ram[4][13] ;
   wire \ram[4][12] ;
   wire \ram[4][11] ;
   wire \ram[4][10] ;
   wire \ram[4][9] ;
   wire \ram[4][8] ;
   wire \ram[4][7] ;
   wire \ram[4][6] ;
   wire \ram[4][5] ;
   wire \ram[4][4] ;
   wire \ram[4][3] ;
   wire \ram[4][2] ;
   wire \ram[4][1] ;
   wire \ram[4][0] ;
   wire \ram[3][15] ;
   wire \ram[3][14] ;
   wire \ram[3][13] ;
   wire \ram[3][12] ;
   wire \ram[3][11] ;
   wire \ram[3][10] ;
   wire \ram[3][9] ;
   wire \ram[3][8] ;
   wire \ram[3][7] ;
   wire \ram[3][6] ;
   wire \ram[3][5] ;
   wire \ram[3][4] ;
   wire \ram[3][3] ;
   wire \ram[3][2] ;
   wire \ram[3][1] ;
   wire \ram[3][0] ;
   wire \ram[2][15] ;
   wire \ram[2][14] ;
   wire \ram[2][13] ;
   wire \ram[2][12] ;
   wire \ram[2][11] ;
   wire \ram[2][10] ;
   wire \ram[2][9] ;
   wire \ram[2][8] ;
   wire \ram[2][7] ;
   wire \ram[2][6] ;
   wire \ram[2][5] ;
   wire \ram[2][4] ;
   wire \ram[2][3] ;
   wire \ram[2][2] ;
   wire \ram[2][1] ;
   wire \ram[2][0] ;
   wire \ram[1][15] ;
   wire \ram[1][14] ;
   wire \ram[1][13] ;
   wire \ram[1][12] ;
   wire \ram[1][11] ;
   wire \ram[1][10] ;
   wire \ram[1][9] ;
   wire \ram[1][8] ;
   wire \ram[1][7] ;
   wire \ram[1][6] ;
   wire \ram[1][5] ;
   wire \ram[1][4] ;
   wire \ram[1][3] ;
   wire \ram[1][2] ;
   wire \ram[1][1] ;
   wire \ram[1][0] ;
   wire \ram[0][15] ;
   wire \ram[0][14] ;
   wire \ram[0][13] ;
   wire \ram[0][12] ;
   wire \ram[0][11] ;
   wire \ram[0][10] ;
   wire \ram[0][9] ;
   wire \ram[0][8] ;
   wire \ram[0][7] ;
   wire \ram[0][6] ;
   wire \ram[0][5] ;
   wire \ram[0][4] ;
   wire \ram[0][3] ;
   wire \ram[0][2] ;
   wire \ram[0][1] ;
   wire \ram[0][0] ;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3368;
   wire n3369;
   wire n3370;
   wire n3371;
   wire n3372;
   wire n3373;
   wire n3374;
   wire n3375;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3412;
   wire n3413;
   wire n3414;
   wire n3415;
   wire n3416;
   wire n3417;
   wire n3418;
   wire n3419;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3459;
   wire n3460;
   wire n3461;
   wire n3462;
   wire n3463;
   wire n3464;
   wire n3465;
   wire n3466;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n3594;
   wire n3595;
   wire n3596;
   wire n3597;
   wire n3598;
   wire n3599;
   wire n3600;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3619;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3630;
   wire n3631;
   wire n3632;
   wire n3633;
   wire n3634;
   wire n3635;
   wire n3636;
   wire n3637;
   wire n3638;
   wire n3639;
   wire n3640;
   wire n3641;
   wire n3642;
   wire n3643;
   wire n3644;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3648;
   wire n3649;
   wire n3650;
   wire n3651;
   wire n3652;
   wire n3653;
   wire n3654;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3658;
   wire n3659;
   wire n3660;
   wire n3661;
   wire n3662;
   wire n3663;
   wire n3664;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3668;
   wire n3669;
   wire n3670;
   wire n3671;
   wire n3672;
   wire n3673;
   wire n3674;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3679;
   wire n3680;
   wire n3681;
   wire n3682;
   wire n3683;
   wire n3684;
   wire n3685;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3689;
   wire n3690;
   wire n3691;
   wire n3692;
   wire n3693;
   wire n3694;
   wire n3695;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3699;
   wire n3700;
   wire n3701;
   wire n3702;
   wire n3703;
   wire n3704;
   wire n3705;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3709;
   wire n3710;
   wire n3711;
   wire n3712;
   wire n3713;
   wire n3714;
   wire n3715;
   wire n3716;
   wire n3717;
   wire n3718;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3759;
   wire n3760;
   wire n3761;
   wire n3762;
   wire n3763;
   wire n3764;
   wire n3765;
   wire n3766;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3770;
   wire n3771;
   wire n3772;
   wire n3773;
   wire n3774;
   wire n3775;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3779;
   wire n3780;
   wire n3781;
   wire n3782;
   wire n3783;
   wire n3784;
   wire n3785;
   wire n3786;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3790;
   wire n3791;
   wire n3792;
   wire n3793;
   wire n3794;
   wire n3795;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3799;
   wire n3800;
   wire n3801;
   wire n3802;
   wire n3803;
   wire n3804;
   wire n3805;
   wire n3806;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3810;
   wire n3811;
   wire n3812;
   wire n3813;
   wire n3814;
   wire n3815;
   wire n3816;
   wire n3817;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3821;
   wire n3822;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3836;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire n3844;
   wire n3845;
   wire n3846;
   wire n3847;
   wire n3848;
   wire n3849;
   wire n3850;
   wire n3851;
   wire n3852;
   wire n3853;
   wire n3854;
   wire n3855;
   wire n3856;
   wire n3857;
   wire n3858;
   wire n3859;
   wire n3860;
   wire n3861;
   wire n3862;
   wire n3863;
   wire n3864;
   wire n3865;
   wire n3866;
   wire n3867;
   wire n3868;
   wire n3869;
   wire n3870;
   wire n3871;
   wire n3872;
   wire n3873;
   wire n3874;
   wire n3875;
   wire n3876;
   wire n3877;
   wire n3878;
   wire n3879;
   wire n3880;
   wire n3881;
   wire n3882;
   wire n3883;
   wire n3884;
   wire n3885;
   wire n3886;
   wire n3887;
   wire n3888;
   wire n3889;
   wire n3890;
   wire n3891;
   wire n3892;
   wire n3893;
   wire n3894;
   wire n3895;
   wire n3896;
   wire n3897;
   wire n3898;
   wire n3899;
   wire n3900;
   wire n3901;
   wire n3902;
   wire n3903;
   wire n3904;
   wire n3905;
   wire n3906;
   wire n3907;
   wire n3908;
   wire n3909;
   wire n3910;
   wire n3911;
   wire n3912;
   wire n3913;
   wire n3914;
   wire n3915;
   wire n3916;
   wire n3917;
   wire n3918;
   wire n3919;
   wire n3920;
   wire n3921;
   wire n3922;
   wire n3923;
   wire n3924;
   wire n3925;
   wire n3926;
   wire n3927;
   wire n3928;
   wire n3929;
   wire n3930;
   wire n3931;
   wire n3932;
   wire n3933;
   wire n3934;
   wire n3935;
   wire n3936;
   wire n3937;
   wire n3938;
   wire n3939;
   wire n3940;
   wire n3941;
   wire n3942;
   wire n3943;
   wire n3944;
   wire n3945;
   wire n3946;
   wire n3947;
   wire n3948;
   wire n3949;
   wire n3950;
   wire n3951;
   wire n3952;
   wire n3953;
   wire n3954;
   wire n3955;
   wire n3956;
   wire n3957;
   wire n3958;
   wire n3959;
   wire n3960;
   wire n3961;
   wire n3962;
   wire n3963;
   wire n3964;
   wire n3965;
   wire n3966;
   wire n3967;
   wire n3968;
   wire n3969;
   wire n3970;
   wire n3971;
   wire n3972;
   wire n3973;
   wire n3974;
   wire n3975;
   wire n3976;
   wire n3977;
   wire n3978;
   wire n3979;
   wire n3980;
   wire n3981;
   wire n3982;
   wire n3983;
   wire n3984;
   wire n3985;
   wire n3986;
   wire n3987;
   wire n3988;
   wire n3989;
   wire n3990;
   wire n3991;
   wire n3992;
   wire n3993;
   wire n3994;
   wire n3995;
   wire n3996;
   wire n3997;
   wire n3998;
   wire n3999;
   wire n4000;
   wire n4001;
   wire n4002;
   wire n4003;
   wire n4004;
   wire n4005;
   wire n4006;
   wire n4007;
   wire n4008;
   wire n4009;
   wire n4010;
   wire n4011;
   wire n4012;
   wire n4013;
   wire n4014;
   wire n4015;
   wire n4016;
   wire n4017;
   wire n4018;
   wire n4019;
   wire n4020;
   wire n4021;
   wire n4022;
   wire n4023;
   wire n4024;
   wire n4025;
   wire n4026;
   wire n4027;
   wire n4028;
   wire n4029;
   wire n4030;
   wire n4031;
   wire n4032;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4036;
   wire n4037;
   wire n4038;
   wire n4039;
   wire n4040;
   wire n4041;
   wire n4042;
   wire n4043;
   wire n4044;
   wire n4045;
   wire n4046;
   wire n4047;
   wire n4048;
   wire n4049;
   wire n4050;
   wire n4051;
   wire n4052;
   wire n4053;
   wire n4054;
   wire n4055;
   wire n4056;
   wire n4057;
   wire n4058;
   wire n4059;
   wire n4060;
   wire n4061;
   wire n4062;
   wire n4063;
   wire n4064;
   wire n4065;
   wire n4066;
   wire n4067;
   wire n4068;
   wire n4069;
   wire n4070;
   wire n4071;
   wire n4072;
   wire n4073;
   wire n4074;
   wire n4075;
   wire n4076;
   wire n4077;
   wire n4078;
   wire n4079;
   wire n4080;
   wire n4081;
   wire n4082;
   wire n4083;
   wire n4084;
   wire n4085;
   wire n4086;
   wire n4087;
   wire n4088;
   wire n4089;
   wire n4090;
   wire n4091;
   wire n4092;
   wire n4093;
   wire n4094;
   wire n4095;
   wire n4096;
   wire n4097;
   wire n4098;
   wire n4099;
   wire n4100;
   wire n4101;
   wire n4102;
   wire n4103;
   wire n4104;
   wire n4105;
   wire n4106;
   wire n4107;
   wire n4108;
   wire n4109;
   wire n4110;
   wire n4111;
   wire n4112;
   wire n4113;
   wire n4114;
   wire n4115;
   wire n4116;
   wire n4117;
   wire n4118;
   wire n4119;
   wire n4120;
   wire n4121;
   wire n4122;
   wire n4123;
   wire n4124;
   wire n4125;
   wire n4126;
   wire n4127;
   wire n4128;
   wire n4129;
   wire n4130;
   wire n4131;
   wire n4132;
   wire n4133;
   wire n4134;
   wire n4135;
   wire n4136;
   wire n4137;
   wire n4138;
   wire n4139;
   wire n4140;
   wire n4141;
   wire n4142;
   wire n4143;
   wire n4144;
   wire n4145;
   wire n4146;
   wire n4147;
   wire n4148;
   wire n4149;
   wire n4150;
   wire n4151;
   wire n4152;
   wire n4153;
   wire n4154;
   wire n4155;
   wire n4156;
   wire n4157;
   wire n4158;
   wire n4159;
   wire n4160;
   wire n4161;
   wire n4162;
   wire n4163;
   wire n4164;
   wire n4165;
   wire n4166;
   wire n4167;
   wire n4168;
   wire n4169;
   wire n4170;
   wire n4171;
   wire n4172;
   wire n4173;
   wire n4174;
   wire n4175;
   wire n4176;
   wire n4177;
   wire n4178;
   wire n4179;
   wire n4180;
   wire n4181;
   wire n4182;
   wire n4183;
   wire n4184;
   wire n4185;
   wire n4186;
   wire n4187;
   wire n4188;
   wire n4189;
   wire n4190;
   wire n4191;
   wire n4192;
   wire n4193;
   wire n4194;
   wire n4195;
   wire n4196;
   wire n4197;
   wire n4198;
   wire n4199;
   wire n4200;
   wire n4201;
   wire n4202;
   wire n4203;
   wire n4204;
   wire n4205;
   wire n4206;
   wire n4207;
   wire n4208;
   wire n4209;
   wire n4210;
   wire n4211;
   wire n4212;
   wire n4213;
   wire n4214;
   wire n4215;
   wire n4216;
   wire n4217;
   wire n4218;
   wire n4219;
   wire n4220;
   wire n4221;
   wire n4222;
   wire n4223;
   wire n4224;
   wire n4225;
   wire n4226;
   wire n4227;
   wire n4228;
   wire n4229;
   wire n4230;
   wire n4231;
   wire n4232;
   wire n4233;
   wire n4234;
   wire n4235;
   wire n4236;
   wire n4237;
   wire n4238;
   wire n4239;
   wire n4240;
   wire n4241;
   wire n4242;
   wire n4243;
   wire n4244;
   wire n4245;
   wire n4246;
   wire n4247;
   wire n4248;
   wire n4249;
   wire n4250;
   wire n4251;
   wire n4252;
   wire n4253;
   wire n4254;
   wire n4255;
   wire n4256;
   wire n4257;
   wire n4258;
   wire n4259;
   wire n4260;
   wire n4261;
   wire n4262;
   wire n4263;
   wire n4264;
   wire n4265;
   wire n4266;
   wire n4267;
   wire n4268;
   wire n4269;
   wire n4270;
   wire n4271;
   wire n4272;
   wire n4273;
   wire n4274;
   wire n4275;
   wire n4276;
   wire n4277;
   wire n4278;
   wire n4279;
   wire n4280;
   wire n4281;
   wire n4282;
   wire n4283;
   wire n4284;
   wire n4285;
   wire n4286;
   wire n4287;
   wire n4288;
   wire n4289;
   wire n4290;
   wire n4291;
   wire n4292;
   wire n4293;
   wire n4294;
   wire n4295;
   wire n4296;
   wire n4297;
   wire n4298;
   wire n4299;
   wire n4300;
   wire n4301;
   wire n4302;
   wire n4303;
   wire n4304;
   wire n4305;
   wire n4306;
   wire n4307;
   wire n4308;
   wire n4309;
   wire n4310;
   wire n4311;
   wire n4312;
   wire n4313;
   wire n4314;
   wire n4315;
   wire n4316;
   wire n4317;
   wire n4318;
   wire n4319;
   wire n4320;
   wire n4321;
   wire n4322;
   wire n4323;
   wire n4324;
   wire n4325;
   wire n4326;
   wire n4327;
   wire n4328;
   wire n4329;
   wire n4330;
   wire n4331;
   wire n4332;
   wire n4333;
   wire n4334;
   wire n4335;
   wire n4336;
   wire n4337;
   wire n4338;
   wire n4339;
   wire n4340;
   wire n4341;
   wire n4342;
   wire n4343;
   wire n4344;
   wire n4345;
   wire n4346;
   wire n4347;
   wire n4348;
   wire n4349;
   wire n4350;
   wire n4351;
   wire n4352;
   wire n4353;
   wire n4354;
   wire n4355;
   wire n4356;
   wire n4357;
   wire n4358;
   wire n4359;
   wire n4360;
   wire n4361;
   wire n4362;
   wire n4363;
   wire n4364;
   wire n4365;
   wire n4366;
   wire n4367;
   wire n4368;
   wire n4369;
   wire n4370;
   wire n4371;
   wire n4372;
   wire n4373;
   wire n4374;
   wire n4375;
   wire n4376;
   wire n4377;
   wire n4378;
   wire n4379;
   wire n4380;
   wire n4381;
   wire n4382;
   wire n4383;
   wire n4384;
   wire n4385;
   wire n4386;
   wire n4387;
   wire n4388;
   wire n4389;
   wire n4390;
   wire n4391;
   wire n4392;
   wire n4393;
   wire n4394;
   wire n4395;
   wire n4396;
   wire n4397;
   wire n4398;
   wire n4399;
   wire n4400;
   wire n4401;
   wire n4402;
   wire n4403;
   wire n4404;
   wire n4405;
   wire n4406;
   wire n4407;
   wire n4408;
   wire n4409;
   wire n4410;
   wire n4411;
   wire n4412;
   wire n4413;
   wire n4414;
   wire n4415;
   wire n4416;
   wire n4417;
   wire n4418;
   wire n4419;
   wire n4420;
   wire n4421;
   wire n4422;
   wire n4423;
   wire n4424;
   wire n4425;
   wire n4426;
   wire n4427;
   wire n4428;
   wire n4429;
   wire n4430;
   wire n4431;
   wire n4432;
   wire n4433;
   wire n4434;
   wire n4435;
   wire n4436;
   wire n4437;
   wire n4438;
   wire n4439;
   wire n4440;
   wire n4441;
   wire n4442;
   wire n4443;
   wire n4444;
   wire n4445;
   wire n4446;
   wire n4447;
   wire n4448;
   wire n4449;
   wire n4450;
   wire n4451;
   wire n4452;
   wire n4453;
   wire n4454;
   wire n4455;
   wire n4456;
   wire n4457;
   wire n4458;
   wire n4459;
   wire n4460;
   wire n4461;
   wire n4462;
   wire n4463;
   wire n4464;
   wire n4465;
   wire n4466;
   wire n4467;
   wire n4468;
   wire n4469;
   wire n4470;
   wire n4471;
   wire n4472;
   wire n4473;
   wire n4474;
   wire n4475;
   wire n4476;
   wire n4477;
   wire n4478;
   wire n4479;
   wire n4480;
   wire n4481;
   wire n4482;
   wire n4483;
   wire n4484;
   wire n4485;
   wire n4486;
   wire n4487;
   wire n4488;
   wire n4489;
   wire n4490;
   wire n4491;
   wire n4492;
   wire n4493;
   wire n4494;
   wire n4495;
   wire n4496;
   wire n4497;
   wire n4498;
   wire n4499;
   wire n4500;
   wire n4501;
   wire n4502;
   wire n4503;
   wire n4504;
   wire n4505;
   wire n4506;
   wire n4507;
   wire n4508;
   wire n4509;
   wire n4510;
   wire n4511;
   wire n4512;
   wire n4513;
   wire n4514;
   wire n4515;
   wire n4516;
   wire n4517;
   wire n4518;
   wire n4519;
   wire n4520;
   wire n4521;
   wire n4522;
   wire n4523;
   wire n4524;
   wire n4525;
   wire n4526;
   wire n4527;
   wire n4528;
   wire n4529;
   wire n4530;
   wire n4531;
   wire n4532;
   wire n4533;
   wire n4534;
   wire n4535;
   wire n4536;
   wire n4537;
   wire n4538;
   wire n4539;
   wire n4540;
   wire n4541;
   wire n4542;
   wire n4543;
   wire n4544;
   wire n4545;
   wire n4546;
   wire n4547;
   wire n4548;
   wire n4549;
   wire n4550;
   wire n4551;
   wire n4552;
   wire n4553;
   wire n4554;
   wire n4555;
   wire n4556;
   wire n4557;
   wire n4558;
   wire n4559;
   wire n4560;
   wire n4561;
   wire n4562;
   wire n4563;
   wire n4564;
   wire n4565;
   wire n4566;
   wire n4567;
   wire n4568;
   wire n4569;
   wire n4570;
   wire n4571;
   wire n4572;
   wire n4573;
   wire n4574;
   wire n4575;
   wire n4576;
   wire n4577;
   wire n4578;
   wire n4579;
   wire n4580;
   wire n4581;
   wire n4582;
   wire n4583;
   wire n4584;
   wire n4585;
   wire n4586;
   wire n4587;
   wire n4588;
   wire n4589;
   wire n4590;
   wire n4591;
   wire n4592;
   wire n4593;
   wire n4594;
   wire n4595;
   wire n4596;
   wire n4597;
   wire n4598;
   wire n4599;
   wire n4600;
   wire n4601;
   wire n4602;
   wire n4603;
   wire n4604;
   wire n4605;
   wire n4606;
   wire n4607;
   wire n4608;
   wire n4609;
   wire n4610;
   wire n4611;
   wire n4612;
   wire n4613;
   wire n4614;
   wire n4615;
   wire n4616;
   wire n4617;
   wire n4618;
   wire n4619;
   wire n4620;
   wire n4621;
   wire n4622;
   wire n4623;
   wire n4624;
   wire n4625;
   wire n4626;
   wire n4627;
   wire n4628;
   wire n4629;
   wire n4630;
   wire n4631;
   wire n4632;
   wire n4633;
   wire n4634;
   wire n4635;
   wire n4636;
   wire n4637;
   wire n4638;
   wire n4639;
   wire n4640;
   wire n4641;
   wire n4642;
   wire n4643;
   wire n4644;
   wire n4645;
   wire n4646;
   wire n4647;
   wire n4648;
   wire n4649;
   wire n4650;
   wire n4651;
   wire n4652;
   wire n4653;
   wire n4654;
   wire n4655;
   wire n4656;
   wire n4657;
   wire n4658;
   wire n4659;
   wire n4660;
   wire n4661;
   wire n4662;
   wire n4663;
   wire n4664;
   wire n4665;
   wire n4666;
   wire n4667;
   wire n4668;
   wire n4669;
   wire n4670;
   wire n4671;
   wire n4672;
   wire n4673;
   wire n4674;
   wire n4675;
   wire n4676;
   wire n4677;
   wire n6304;
   wire n6305;
   wire n6306;
   wire n6307;
   wire n6308;
   wire n6309;
   wire n6310;
   wire n6311;
   wire n6312;
   wire n6313;
   wire n6314;
   wire n6315;
   wire n6316;
   wire n6317;
   wire n6318;
   wire n6319;
   wire n6320;
   wire n6321;
   wire n6322;
   wire n6323;
   wire n6324;
   wire n6325;
   wire n6326;
   wire n6327;
   wire n6328;
   wire n6329;
   wire n6330;
   wire n6331;
   wire n6332;
   wire n6333;
   wire n6334;
   wire n6335;
   wire n6336;
   wire n6337;
   wire n6338;
   wire n6339;
   wire n6340;
   wire n6341;
   wire n6342;
   wire n6343;
   wire n6344;
   wire n6345;
   wire n6346;
   wire n6347;
   wire n6348;
   wire n6349;
   wire n6350;
   wire n6351;
   wire n6352;
   wire n6353;
   wire n6354;
   wire n6355;
   wire n6356;
   wire n6357;
   wire n6358;
   wire n6359;
   wire n6360;
   wire n6361;
   wire n6362;
   wire n6363;
   wire n6364;
   wire n6365;
   wire n6366;
   wire n6367;
   wire n6368;
   wire n6369;
   wire n6370;
   wire n6371;
   wire n6372;
   wire n6373;
   wire n6374;
   wire n6375;
   wire n6376;
   wire n6377;
   wire n6378;
   wire n6379;
   wire n6380;
   wire n6381;
   wire n6382;
   wire n6383;
   wire n6384;
   wire n6385;
   wire n6386;
   wire n6387;
   wire n6388;
   wire n6389;
   wire n6390;
   wire n6391;
   wire n6392;
   wire n6393;
   wire n6394;
   wire n6395;
   wire n6396;
   wire n6397;
   wire n6398;
   wire n6399;
   wire n6400;
   wire n6401;
   wire n6402;
   wire n6403;
   wire n6404;
   wire n6405;
   wire n6406;
   wire n6407;
   wire n6408;
   wire n6409;
   wire n6410;
   wire n6411;
   wire n6412;
   wire n6413;
   wire n6414;
   wire n6415;
   wire n6416;
   wire n6417;
   wire n6418;
   wire n6419;
   wire n6420;
   wire n6421;
   wire n6422;
   wire n6423;
   wire n6424;
   wire n6425;
   wire n6426;
   wire n6427;
   wire n6428;
   wire n6429;
   wire n6430;
   wire n6431;
   wire n6432;
   wire n6433;
   wire n6434;
   wire n6435;
   wire n6436;
   wire n6437;
   wire n6438;
   wire n6439;
   wire n6440;
   wire n6441;
   wire n6442;
   wire n6443;
   wire n6444;
   wire n6445;
   wire n6446;
   wire n6447;
   wire n6448;
   wire n6449;
   wire n6450;
   wire n6451;
   wire n6452;
   wire n6453;
   wire n6454;
   wire n6455;
   wire n6456;
   wire n6457;
   wire n6458;
   wire n6459;
   wire n6460;
   wire n6461;
   wire n6462;
   wire n6463;
   wire n6464;
   wire n6465;
   wire n6466;
   wire n6467;
   wire n6468;
   wire n6469;
   wire n6470;
   wire n6471;
   wire n6472;
   wire n6473;
   wire n6474;
   wire n6475;
   wire n6476;
   wire n6477;
   wire n6478;
   wire n6479;
   wire n6480;
   wire n6481;
   wire n6482;
   wire n6483;
   wire n6484;
   wire n6485;
   wire n6486;
   wire n6487;
   wire n6488;
   wire n6489;
   wire n6490;
   wire n6491;
   wire n6492;
   wire n6493;
   wire n6494;
   wire n6495;
   wire n6496;
   wire n6497;
   wire n6498;
   wire n6499;
   wire n6500;
   wire n6501;
   wire n6502;
   wire n6503;
   wire n6504;
   wire n6505;
   wire n6506;
   wire n6507;
   wire n6508;
   wire n6509;
   wire n6510;
   wire n6511;
   wire n6512;
   wire n6513;
   wire n6514;
   wire n6515;
   wire n6516;
   wire n6517;
   wire n6518;
   wire n6519;
   wire n6520;
   wire n6521;
   wire n6522;
   wire n6523;
   wire n6524;
   wire n6525;
   wire n6526;
   wire n6527;
   wire n6528;
   wire n6529;
   wire n6530;
   wire n6531;
   wire n6532;
   wire n6533;
   wire n6534;
   wire n6535;
   wire n6536;
   wire n6537;
   wire n6538;
   wire n6539;
   wire n6540;
   wire n6541;
   wire n6542;
   wire n6543;
   wire n6544;
   wire n6545;
   wire n6546;
   wire n6547;
   wire n6548;
   wire n6549;
   wire n6550;
   wire n6551;
   wire n6552;
   wire n6553;
   wire n6554;
   wire n6555;
   wire n6556;
   wire n6557;
   wire n6558;
   wire n6559;
   wire n6560;
   wire n6561;
   wire n6562;
   wire n6563;
   wire n6564;
   wire n6565;
   wire n6566;
   wire n6567;
   wire n6568;
   wire n6569;
   wire n6570;
   wire n6571;
   wire n6572;
   wire n6573;
   wire n6574;
   wire n6575;
   wire n6576;
   wire n6577;
   wire n6578;
   wire n6579;
   wire n6580;
   wire n6581;
   wire n6582;
   wire n6583;
   wire n6584;
   wire n6585;
   wire n6586;
   wire n6587;
   wire n6588;
   wire n6589;
   wire n6590;
   wire n6591;
   wire n6592;
   wire n6593;
   wire n6594;
   wire n6595;
   wire n6596;
   wire n6597;
   wire n6598;
   wire n6599;
   wire n6600;
   wire n6601;
   wire n6602;
   wire n6603;
   wire n6604;
   wire n6605;
   wire n6606;
   wire n6607;
   wire n6608;
   wire n6609;
   wire n6610;
   wire n6611;
   wire n6612;
   wire n6613;
   wire n6614;
   wire n6615;
   wire n6616;
   wire n6617;
   wire n6618;
   wire n6619;
   wire n6620;
   wire n6621;
   wire n6622;
   wire n6623;
   wire n6624;
   wire n6625;
   wire n6626;
   wire n6627;
   wire n6628;
   wire n6629;
   wire n6630;
   wire n6631;
   wire n6632;
   wire n6633;
   wire n6634;
   wire n6635;
   wire n6636;
   wire n6637;
   wire n6638;
   wire n6639;
   wire n6640;
   wire n6641;
   wire n6642;
   wire n6643;
   wire n6644;
   wire n6645;
   wire n6646;
   wire n6647;
   wire n6648;
   wire n6649;
   wire n6650;
   wire n6651;
   wire n6652;
   wire n6653;
   wire n6654;
   wire n6655;
   wire n6656;
   wire n6657;
   wire n6658;
   wire n6659;
   wire n6660;
   wire n6661;
   wire n6662;
   wire n6663;
   wire n6664;
   wire n6665;
   wire n6666;
   wire n6667;
   wire n6668;
   wire n6669;
   wire n6670;
   wire n6671;
   wire n6672;
   wire n6673;
   wire n6674;
   wire n6675;
   wire n6676;
   wire n6677;
   wire n6678;
   wire n6679;
   wire n6680;
   wire n6681;
   wire n6682;
   wire n6683;
   wire n6684;
   wire n6685;
   wire n6686;
   wire n6687;
   wire n6688;
   wire n6689;
   wire n6690;
   wire n6691;
   wire n6692;
   wire n6693;
   wire n6694;
   wire n6695;
   wire n6696;
   wire n6697;
   wire n6698;
   wire n6699;
   wire n6700;
   wire n6701;
   wire n6702;
   wire n6703;
   wire n6704;
   wire n6705;
   wire n6706;
   wire n6707;
   wire n6708;
   wire n6709;
   wire n6710;
   wire n6711;
   wire n6712;
   wire n6713;
   wire n6714;
   wire n6715;
   wire n6716;
   wire n6717;
   wire n6718;
   wire n6719;
   wire n6720;
   wire n6721;
   wire n6722;
   wire n6723;
   wire n6724;
   wire n6725;
   wire n6726;
   wire n6727;
   wire n6728;
   wire n6729;
   wire n6730;
   wire n6731;
   wire n6732;
   wire n6733;
   wire n6734;
   wire n6735;
   wire n6736;
   wire n6737;
   wire n6738;
   wire n6739;
   wire n6740;
   wire n6741;
   wire n6742;
   wire n6743;
   wire n6744;
   wire n6745;
   wire n6746;
   wire n6747;
   wire n6748;
   wire n6749;
   wire n6750;
   wire n6751;
   wire n6752;
   wire n6753;
   wire n6754;
   wire n6755;
   wire n6756;
   wire n6757;
   wire n6758;
   wire n6759;
   wire n6760;
   wire n6761;
   wire n6762;
   wire n6763;
   wire n6764;
   wire n6765;
   wire n6766;
   wire n6767;
   wire n6768;
   wire n6769;
   wire n6770;
   wire n6771;
   wire n6772;
   wire n6773;
   wire n6774;
   wire n6775;
   wire n6776;
   wire n6777;
   wire n6778;
   wire n6779;
   wire n6780;
   wire n6781;
   wire n6782;
   wire n6783;
   wire n6784;
   wire n6785;
   wire n6786;
   wire n6787;
   wire n6788;
   wire n6789;
   wire n6790;
   wire n6791;
   wire n6792;
   wire n6793;
   wire n6794;
   wire n6795;
   wire n6796;
   wire n6797;
   wire n6798;
   wire n6799;
   wire n6800;
   wire n6801;
   wire n6802;
   wire n6803;
   wire n6804;
   wire n6805;
   wire n6806;
   wire n6807;
   wire n6808;
   wire n6809;
   wire n6810;
   wire n6811;
   wire n6812;
   wire n6813;
   wire n6814;
   wire n6815;
   wire n6816;
   wire n6817;
   wire n6818;
   wire n6819;
   wire n6820;
   wire n6821;
   wire n6822;
   wire n6823;
   wire n6824;
   wire n6825;
   wire n6826;
   wire n6827;
   wire n6828;
   wire n6829;
   wire n6830;
   wire n6831;
   wire n6832;
   wire n6833;
   wire n6834;
   wire n6835;
   wire n6836;
   wire n6837;
   wire n6838;
   wire n6839;
   wire n6840;
   wire n6841;
   wire n6842;
   wire n6843;
   wire n6844;
   wire n6845;
   wire n6846;
   wire n6847;
   wire n6848;
   wire n6849;
   wire n6850;
   wire n6851;
   wire n6852;
   wire n6853;
   wire n6854;
   wire n6855;
   wire n6856;
   wire n6857;
   wire n6858;
   wire n6859;
   wire n6860;
   wire n6861;
   wire n6862;
   wire n6863;
   wire n6864;
   wire n6865;
   wire n6866;
   wire n6867;
   wire n6868;
   wire n6869;
   wire n6870;
   wire n6871;
   wire n6872;
   wire n6873;
   wire n6874;
   wire n6875;
   wire n6876;
   wire n6877;
   wire n6878;
   wire n6879;
   wire n6880;
   wire n6881;
   wire n6882;
   wire n6883;
   wire n6884;
   wire n6885;
   wire n6886;
   wire n6887;
   wire n6888;
   wire n6889;
   wire n6890;
   wire n6891;
   wire n6892;
   wire n6893;
   wire n6894;
   wire n6895;
   wire n6896;
   wire n6897;
   wire n6898;
   wire n6899;
   wire n6900;
   wire n6901;
   wire n6902;
   wire n6903;
   wire n6904;
   wire n6905;
   wire n6906;
   wire n6907;
   wire n6908;
   wire n6909;
   wire n6910;
   wire n6911;
   wire n6912;
   wire n6913;
   wire n6914;
   wire n6915;
   wire n6916;
   wire n6917;
   wire n6918;
   wire n6919;
   wire n6920;
   wire n6921;
   wire n6922;
   wire n6923;
   wire n6924;
   wire n6925;
   wire n6926;
   wire n6927;
   wire n6928;
   wire n6929;
   wire n6930;
   wire n6931;
   wire n6932;
   wire n6933;
   wire n6934;
   wire n6935;
   wire n6936;
   wire n6937;
   wire n6938;
   wire n6939;
   wire n6940;
   wire n6941;
   wire n6942;
   wire n6943;
   wire n6944;
   wire n6945;
   wire n6946;
   wire n6947;
   wire n6948;
   wire n6949;
   wire n6950;
   wire n6951;
   wire n6952;
   wire n6953;
   wire n6954;
   wire n6955;
   wire n6956;
   wire n6957;
   wire n6958;
   wire n6959;
   wire n6960;
   wire n6961;
   wire n6962;
   wire n6963;
   wire n6964;
   wire n6965;
   wire n6966;
   wire n6967;
   wire n6968;
   wire n6969;
   wire n6970;
   wire n6971;
   wire n6972;
   wire n6973;
   wire n6974;
   wire n6975;
   wire n6976;
   wire n6977;
   wire n6978;
   wire n6979;
   wire n6980;
   wire n6981;
   wire n6982;
   wire n6983;
   wire n6984;
   wire n6985;
   wire n6986;
   wire n6987;
   wire n6988;
   wire n6989;
   wire n6990;
   wire n6991;
   wire n6992;
   wire n6993;
   wire n6994;
   wire n6995;
   wire n6996;
   wire n6997;
   wire n6998;
   wire n6999;
   wire n7000;
   wire n7001;
   wire n7002;
   wire n7003;
   wire n7004;
   wire n7005;
   wire n7006;
   wire n7007;
   wire n7008;
   wire n7009;
   wire n7010;
   wire n7011;
   wire n7012;
   wire n7013;
   wire n7014;
   wire n7015;
   wire n7016;
   wire n7017;
   wire n7018;
   wire n7019;
   wire n7020;
   wire n7021;
   wire n7022;
   wire n7023;
   wire n7024;
   wire n7025;
   wire n7026;
   wire n7027;
   wire n7028;
   wire n7029;
   wire n7030;
   wire n7031;
   wire n7032;
   wire n7033;
   wire n7034;
   wire n7035;
   wire n7036;
   wire n7037;
   wire n7038;
   wire n7039;
   wire n7040;
   wire n7041;
   wire n7042;
   wire n7043;
   wire n7044;
   wire n7045;
   wire n7046;
   wire n7047;
   wire n7048;
   wire n7049;
   wire n7050;
   wire n7051;
   wire n7052;
   wire n7053;
   wire n7054;
   wire n7055;
   wire n7056;
   wire n7057;
   wire n7058;
   wire n7059;
   wire n7060;
   wire n7061;
   wire n7062;
   wire n7063;
   wire n7064;
   wire n7065;
   wire n7066;
   wire n7067;
   wire n7068;
   wire n7069;
   wire n7070;
   wire n7071;
   wire n7072;
   wire n7073;
   wire n7074;
   wire n7075;
   wire n7076;
   wire n7077;
   wire n7078;
   wire n7079;
   wire n7080;
   wire n7081;
   wire n7082;
   wire n7083;
   wire n7084;
   wire n7085;
   wire n7086;
   wire n7087;
   wire n7088;
   wire n7089;
   wire n7090;
   wire n7091;
   wire n7092;
   wire n7093;
   wire n7094;
   wire n7095;
   wire n7096;
   wire n7097;
   wire n7098;
   wire n7099;
   wire n7100;
   wire n7101;
   wire n7102;
   wire n7103;
   wire n7104;
   wire n7105;
   wire n7106;
   wire n7107;
   wire n7108;
   wire n7109;
   wire n7110;
   wire n7111;
   wire n7112;
   wire n7113;
   wire n7114;
   wire n7115;
   wire n7116;
   wire n7117;
   wire n7118;
   wire n7119;
   wire n7120;
   wire n7121;
   wire n7122;
   wire n7123;
   wire n7124;
   wire n7125;
   wire n7126;
   wire n7127;
   wire n7128;
   wire n7129;
   wire n7130;
   wire n7131;
   wire n7132;
   wire n7133;
   wire n7134;
   wire n7135;
   wire n7136;
   wire n7137;
   wire n7138;
   wire n7139;
   wire n7140;
   wire n7141;
   wire n7142;
   wire n7143;
   wire n7144;
   wire n7145;
   wire n7146;
   wire n7147;
   wire n7148;
   wire n7149;
   wire n7150;
   wire n7151;
   wire n7152;
   wire n7153;
   wire n7154;
   wire n7155;
   wire n7156;
   wire n7157;
   wire n7158;
   wire n7159;
   wire n7160;
   wire n7161;
   wire n7162;
   wire n7163;
   wire n7164;
   wire n7165;
   wire n7166;
   wire n7167;
   wire n7168;
   wire n7169;
   wire n7170;
   wire n7171;
   wire n7172;
   wire n7173;
   wire n7174;
   wire n7175;
   wire n7176;
   wire n7177;
   wire n7178;
   wire n7179;
   wire n7180;
   wire n7181;
   wire n7182;
   wire n7183;
   wire n7184;
   wire n7185;
   wire n7186;
   wire n7187;
   wire n7188;
   wire n7189;
   wire n7190;
   wire n7191;
   wire n7192;
   wire n7193;
   wire n7194;
   wire n7195;
   wire n7196;
   wire n7197;
   wire n7198;
   wire n7199;
   wire n7200;
   wire n7201;
   wire n7202;
   wire n7203;
   wire n7204;
   wire n7205;
   wire n7206;
   wire n7207;
   wire n7208;
   wire n7209;
   wire n7210;
   wire n7211;
   wire n7212;
   wire n7213;
   wire n7214;
   wire n7215;
   wire n7216;
   wire n7217;
   wire n7218;
   wire n7219;
   wire n7220;
   wire n7221;
   wire n7222;
   wire n7223;
   wire n7224;
   wire n7225;
   wire n7226;
   wire n7227;
   wire n7228;
   wire n7229;
   wire n7230;
   wire n7231;
   wire n7232;
   wire n7233;
   wire n7234;
   wire n7235;
   wire n7236;
   wire n7237;
   wire n7238;
   wire n7239;
   wire n7240;
   wire n7241;
   wire n7242;
   wire n7243;
   wire n7244;
   wire n7245;
   wire n7246;
   wire n7247;
   wire n7248;
   wire n7249;
   wire n7250;
   wire n7251;
   wire n7252;
   wire n7253;
   wire n7254;
   wire n7255;
   wire n7256;
   wire n7257;
   wire n7258;
   wire n7259;
   wire n7260;
   wire n7261;
   wire n7262;
   wire n7263;
   wire n7264;
   wire n7265;
   wire n7266;
   wire n7267;
   wire n7268;
   wire n7269;
   wire n7270;
   wire n7271;
   wire n7272;
   wire n7273;
   wire n7274;
   wire n7275;
   wire n7276;
   wire n7277;
   wire n7278;
   wire n7279;
   wire n7280;
   wire n7281;
   wire n7282;
   wire n7283;
   wire n7284;
   wire n7285;
   wire n7286;
   wire n7287;
   wire n7288;
   wire n7289;
   wire n7290;
   wire n7291;
   wire n7292;
   wire n7293;
   wire n7294;
   wire n7295;
   wire n7296;
   wire n7297;
   wire n7298;
   wire n7299;
   wire n7300;
   wire n7301;
   wire n7302;
   wire n7303;
   wire n7304;
   wire n7305;
   wire n7306;
   wire n7307;
   wire n7308;
   wire n7309;
   wire n7310;
   wire n7311;
   wire n7312;
   wire n7313;
   wire n7314;
   wire n7315;
   wire n7316;
   wire n7317;
   wire n7318;
   wire n7319;
   wire n7320;
   wire n7321;
   wire n7322;
   wire n7323;
   wire n7324;
   wire n7325;
   wire n7326;
   wire n7327;
   wire n7328;
   wire n7329;
   wire n7330;
   wire n7331;
   wire n7332;
   wire n7333;
   wire n7334;
   wire n7335;
   wire n7336;
   wire n7337;
   wire n7338;
   wire n7339;
   wire n7340;
   wire n7341;
   wire n7342;
   wire n7343;
   wire n7344;
   wire n7345;
   wire n7346;
   wire n7347;
   wire n7348;
   wire n7349;
   wire n7350;
   wire n7351;
   wire n7352;
   wire n7353;
   wire n7354;
   wire n7355;
   wire n7356;
   wire n7357;
   wire n7358;
   wire n7359;
   wire n7360;
   wire n7361;
   wire n7362;
   wire n7363;
   wire n7364;
   wire n7365;
   wire n7366;
   wire n7367;
   wire n7368;
   wire n7369;
   wire n7370;
   wire n7371;
   wire n7372;
   wire n7373;
   wire n7374;
   wire n7375;
   wire n7376;
   wire n7377;
   wire n7378;
   wire n7379;
   wire n7380;
   wire n7381;
   wire n7382;
   wire n7383;
   wire n7384;
   wire n7385;
   wire n7386;
   wire n7387;
   wire n7388;
   wire n7389;
   wire n7390;
   wire n7391;
   wire n7392;
   wire n7393;
   wire n7394;
   wire n7395;
   wire n7396;
   wire n7397;
   wire n7398;
   wire n7399;
   wire n7400;
   wire n7401;
   wire n7402;
   wire n7403;
   wire n7404;
   wire n7405;
   wire n7406;
   wire n7407;
   wire n7408;
   wire n7409;
   wire n7410;
   wire n7411;
   wire n7412;
   wire n7413;
   wire n7414;
   wire n7415;
   wire n7416;
   wire n7417;
   wire n7418;
   wire n7419;
   wire n7420;
   wire n7421;
   wire n7422;
   wire n7423;
   wire n7424;
   wire n7425;
   wire n7426;
   wire n7427;
   wire n7428;
   wire n7429;
   wire n7430;
   wire n7431;
   wire n7432;
   wire n7433;
   wire n7434;
   wire n7435;
   wire n7436;
   wire n7437;
   wire n7438;
   wire n7439;
   wire n7440;
   wire n7441;
   wire n7442;
   wire n7443;
   wire n7444;
   wire n7445;
   wire n7446;
   wire n7447;
   wire n7448;
   wire n7449;
   wire n7450;
   wire n7451;
   wire n7452;
   wire n7453;
   wire n7454;
   wire n7455;
   wire n7456;
   wire n7457;
   wire n7458;
   wire n7459;
   wire n7460;
   wire n7461;
   wire n7462;
   wire n7463;
   wire n7464;
   wire n7465;
   wire n7466;
   wire n7467;
   wire n7468;
   wire n7469;
   wire n7470;
   wire n7471;
   wire n7472;
   wire n7473;
   wire n7474;
   wire n7475;
   wire n7476;
   wire n7477;
   wire n7478;
   wire n7479;
   wire n7480;
   wire n7481;
   wire n7482;
   wire n7483;
   wire n7484;
   wire n7485;
   wire n7486;
   wire n7487;
   wire n7488;
   wire n7489;
   wire n7490;
   wire n7491;
   wire n7492;
   wire n7493;
   wire n7494;
   wire n7495;
   wire n7496;
   wire n7497;
   wire n7498;
   wire n7499;
   wire n7500;
   wire n7501;
   wire n7502;
   wire n7503;
   wire n7504;
   wire n7505;
   wire n7506;
   wire n7507;
   wire n7508;
   wire n7509;
   wire n7510;
   wire n7511;
   wire n7512;
   wire n7513;
   wire n7514;
   wire n7515;
   wire n7516;
   wire n7517;
   wire n7518;
   wire n7519;
   wire n7520;
   wire n7521;
   wire n7522;
   wire n7523;
   wire n7524;
   wire n7525;
   wire n7526;
   wire n7527;
   wire n7528;
   wire n7529;
   wire n7530;
   wire n7531;
   wire n7532;
   wire n7533;
   wire n7534;
   wire n7535;
   wire n7536;
   wire n7537;
   wire n7538;
   wire n7539;
   wire n7540;
   wire n7541;
   wire n7542;
   wire n7543;
   wire n7544;
   wire n7545;
   wire n7546;
   wire n7547;
   wire n7548;
   wire n7549;
   wire n7550;
   wire n7551;
   wire n7552;
   wire n7553;
   wire n7554;
   wire n7555;
   wire n7556;
   wire n7557;
   wire n7558;
   wire n7559;
   wire n7560;
   wire n7561;
   wire n7562;
   wire n7563;
   wire n7564;
   wire n7565;
   wire n7566;
   wire n7567;
   wire n7568;
   wire n7569;
   wire n7570;
   wire n7571;
   wire n7572;
   wire n7573;
   wire n7574;
   wire n7575;
   wire n7576;
   wire n7577;
   wire n7578;
   wire n7579;
   wire n7580;
   wire n7581;
   wire n7582;
   wire n7583;
   wire n7584;
   wire n7585;
   wire n7586;
   wire n7587;
   wire n7588;
   wire n7589;
   wire n7590;
   wire n7591;
   wire n7592;
   wire n7593;
   wire n7594;
   wire n7595;
   wire n7596;
   wire n7597;
   wire n7598;
   wire n7599;
   wire n7600;
   wire n7601;
   wire n7602;
   wire n7603;
   wire n7604;
   wire n7605;
   wire n7606;
   wire n7607;
   wire n7608;
   wire n7609;
   wire n7610;
   wire n7611;
   wire n7612;
   wire n7613;
   wire n7614;
   wire n7615;
   wire n7616;
   wire n7617;
   wire n7618;
   wire n7619;
   wire n7620;
   wire n7621;
   wire n7622;
   wire n7623;
   wire n7624;
   wire n7625;
   wire n7626;
   wire n7627;
   wire n7628;
   wire n7629;
   wire n7630;
   wire n7631;
   wire n7632;
   wire n7633;
   wire n7634;
   wire n7635;
   wire n7636;
   wire n7637;
   wire n7638;
   wire n7639;
   wire n7640;
   wire n7641;
   wire n7642;
   wire n7643;
   wire n7644;
   wire n7645;
   wire n7646;
   wire n7647;
   wire n7648;
   wire n7649;
   wire n7650;
   wire n7651;
   wire n7652;
   wire n7653;
   wire n7654;
   wire n7655;
   wire n7656;
   wire n7657;
   wire n7658;
   wire n7659;
   wire n7660;
   wire n7661;
   wire n7662;
   wire n7663;
   wire n7664;
   wire n7665;
   wire n7666;
   wire n7667;
   wire n7668;
   wire n7669;
   wire n7670;
   wire n7671;
   wire n7672;
   wire n7673;
   wire n7674;
   wire n7675;
   wire n7676;
   wire n7677;
   wire n7678;
   wire n7679;
   wire n7680;
   wire n7681;
   wire n7682;
   wire n7683;
   wire n7684;
   wire n7685;
   wire n7686;
   wire n7687;
   wire n7688;
   wire n7689;
   wire n7690;
   wire n7691;
   wire n7692;
   wire n7693;
   wire n7694;
   wire n7695;
   wire n7696;
   wire n7697;
   wire n7698;
   wire n7699;
   wire n7700;
   wire n7701;
   wire n7702;
   wire n7703;
   wire n7704;
   wire n7705;
   wire n7706;
   wire n7707;
   wire n7708;
   wire n7709;
   wire n7710;
   wire n7711;
   wire n7712;
   wire n7713;
   wire n7714;
   wire n7715;
   wire n7716;
   wire n7717;
   wire n7718;
   wire n7719;
   wire n7720;
   wire n7721;
   wire n7722;
   wire n7723;
   wire n7724;
   wire n7725;
   wire n7726;
   wire n7727;
   wire n7728;
   wire n7729;
   wire n7730;
   wire n7731;
   wire n7732;
   wire n7733;
   wire n7734;
   wire n7735;
   wire n7736;
   wire n7737;
   wire n7738;
   wire n7739;
   wire n7740;
   wire n7741;
   wire n7742;
   wire n7743;
   wire n7744;
   wire n7745;
   wire n7746;
   wire n7747;
   wire n7748;
   wire n7749;
   wire n7750;
   wire n7751;
   wire n7752;
   wire n7753;
   wire n7754;
   wire n7755;
   wire n7756;
   wire n7757;
   wire n7758;
   wire n7759;
   wire n7760;
   wire n7761;
   wire n7762;
   wire n7763;
   wire n7764;
   wire n7765;
   wire n7766;
   wire n7767;
   wire n7768;
   wire n7769;
   wire n7770;
   wire n7771;
   wire n7772;
   wire n7773;
   wire n7774;
   wire n7775;
   wire n7776;
   wire n7777;
   wire n7778;
   wire n7779;
   wire n7780;
   wire n7781;
   wire n7782;
   wire n7783;
   wire n7784;
   wire n7785;
   wire n7786;
   wire n7787;
   wire n7788;
   wire n7789;
   wire n7790;
   wire n7791;
   wire n7792;
   wire n7793;
   wire n7794;
   wire n7795;
   wire n7796;
   wire n7797;
   wire n7798;
   wire n7799;
   wire n7800;
   wire n7801;
   wire n7802;
   wire n7803;
   wire n7804;
   wire n7805;
   wire n7806;
   wire n7807;
   wire n7808;
   wire n7809;
   wire n7810;
   wire n7811;
   wire n7812;
   wire n7813;
   wire n7814;
   wire n7815;
   wire n7816;
   wire n7817;
   wire n7818;
   wire n7819;
   wire n7820;
   wire n7821;
   wire n7822;
   wire n7823;
   wire n7824;
   wire n7825;
   wire n7826;
   wire n7827;
   wire n7828;
   wire n7829;
   wire n7830;
   wire n7831;
   wire n7832;
   wire n7833;
   wire n7834;
   wire n7835;
   wire n7836;
   wire n7837;
   wire n7838;
   wire n7839;
   wire n7840;
   wire n7841;
   wire n7842;
   wire n7843;
   wire n7844;
   wire n7845;
   wire n7846;
   wire n7847;
   wire n7848;
   wire n7849;
   wire n7850;
   wire n7851;
   wire n7852;
   wire n7853;
   wire n7854;
   wire n7855;
   wire n7856;
   wire n7857;
   wire n7858;
   wire n7859;
   wire n7860;
   wire n7861;
   wire n7862;
   wire n7863;
   wire n7864;
   wire n7865;
   wire n7866;
   wire n7867;
   wire n7868;
   wire n7869;
   wire n7870;
   wire n7871;
   wire n7872;
   wire n7873;
   wire n7874;
   wire n7875;
   wire n7876;
   wire n7877;
   wire n7878;
   wire n7879;
   wire n7880;
   wire n7881;
   wire n7882;
   wire n7883;
   wire n7884;
   wire n7885;
   wire n7886;
   wire n7887;
   wire n7888;
   wire n7889;
   wire n7890;
   wire n7891;
   wire n7892;
   wire n7893;
   wire n7894;
   wire n7895;
   wire n7896;
   wire n7897;
   wire n7898;
   wire n7899;
   wire n7900;
   wire n7901;
   wire n7902;
   wire n7903;
   wire n7904;
   wire n7905;
   wire n7906;
   wire n7907;
   wire n7908;
   wire n7909;
   wire n7910;
   wire n7911;
   wire n7912;
   wire n7913;
   wire n7914;
   wire n7915;
   wire n7916;
   wire n7917;
   wire n7918;
   wire n7919;
   wire n7920;
   wire n7921;
   wire n7922;
   wire n7923;
   wire n7924;
   wire n7925;
   wire n7926;
   wire n7927;
   wire n7928;
   wire n7929;
   wire n7930;
   wire n7931;
   wire n7932;
   wire n7933;
   wire n7934;
   wire n7935;
   wire n7936;
   wire n7937;
   wire n7938;
   wire n7939;
   wire n7940;
   wire n7941;
   wire n7942;
   wire n7943;
   wire n7944;
   wire n7945;
   wire n7946;
   wire n7947;
   wire n7948;
   wire n7949;
   wire n7950;
   wire n7951;
   wire n7952;
   wire n7953;
   wire n7954;
   wire n7955;
   wire n7956;
   wire n7957;
   wire n7958;
   wire n7959;
   wire n7960;
   wire n7961;
   wire n7962;
   wire n7963;
   wire n7964;
   wire n7965;
   wire n7966;
   wire n7967;
   wire n7968;
   wire n7969;
   wire n7970;
   wire n7971;
   wire n7972;
   wire n7973;
   wire n7974;
   wire n7975;
   wire n7976;
   wire n7977;
   wire n7978;
   wire n7979;
   wire n7980;
   wire n7981;
   wire n7982;
   wire n7983;
   wire n7984;
   wire n7985;
   wire n7986;
   wire n7987;
   wire n7988;
   wire n7989;
   wire n7990;
   wire n7991;
   wire n7992;
   wire n7993;
   wire n7994;
   wire n7995;
   wire n7996;
   wire n7997;
   wire n7998;
   wire n7999;
   wire n8000;
   wire n8001;
   wire n8002;
   wire n8003;
   wire n8004;
   wire n8005;
   wire n8006;
   wire n8007;
   wire n8008;
   wire n8009;
   wire n8010;
   wire n8011;
   wire n8012;
   wire n8013;
   wire n8014;
   wire n8015;
   wire n8016;
   wire n8017;
   wire n8018;
   wire n8019;
   wire n8020;
   wire n8021;
   wire n8022;
   wire n8023;
   wire n8024;
   wire n8025;
   wire n8026;
   wire n8027;
   wire n8028;
   wire n8029;
   wire n8030;
   wire n8031;
   wire n8032;
   wire n8033;
   wire n8034;
   wire n8035;
   wire n8036;
   wire n8037;
   wire n8038;
   wire n8039;
   wire n8040;
   wire n8041;
   wire n8042;
   wire n8043;
   wire n8044;
   wire n8045;
   wire n8046;
   wire n8047;
   wire n8048;
   wire n8049;
   wire n8050;
   wire n8051;
   wire n8052;
   wire n8053;
   wire n8054;
   wire n8055;
   wire n8056;
   wire n8057;
   wire n8058;
   wire n8059;
   wire n8060;
   wire n8061;
   wire n8062;
   wire n8063;
   wire n8064;
   wire n8065;
   wire n8066;
   wire n8067;
   wire n8068;
   wire n8069;
   wire n8070;
   wire n8071;
   wire n8072;
   wire n8073;
   wire n8074;
   wire n8075;
   wire n8076;
   wire n8077;
   wire n8078;
   wire n8079;
   wire n8080;
   wire n8081;
   wire n8082;
   wire n8083;
   wire n8084;
   wire n8085;
   wire n8086;
   wire n8087;
   wire n8088;
   wire n8089;
   wire n8090;
   wire n8091;
   wire n8092;
   wire n8093;
   wire n8094;
   wire n8095;
   wire n8096;
   wire n8097;
   wire n8098;
   wire n8099;
   wire n8100;
   wire n8101;
   wire n8102;
   wire n8103;
   wire n8104;
   wire n8105;
   wire n8106;
   wire n8107;
   wire n8108;
   wire n8109;
   wire n8110;
   wire n8111;
   wire n8112;
   wire n8113;
   wire n8114;
   wire n8115;
   wire n8116;
   wire n8117;
   wire n8118;
   wire n8119;
   wire n8120;
   wire n8121;
   wire n8122;
   wire n8123;
   wire n8124;
   wire n8125;
   wire n8126;
   wire n8127;
   wire n8128;
   wire n8129;
   wire n8130;
   wire n8131;
   wire n8132;
   wire n8133;
   wire n8134;
   wire n8135;
   wire n8136;
   wire n8137;
   wire n8138;
   wire n8139;
   wire n8140;
   wire n8141;
   wire n8142;
   wire n8143;
   wire n8144;
   wire n8145;
   wire n8146;
   wire n8147;
   wire n8148;
   wire n8149;
   wire n8150;
   wire n8151;
   wire n8152;
   wire n8153;
   wire n8154;
   wire n8155;
   wire n8156;
   wire n8157;
   wire n8158;
   wire n8159;
   wire n8160;
   wire n8161;
   wire n8162;
   wire n8163;
   wire n8164;
   wire n8165;
   wire n8166;
   wire n8167;
   wire n8168;
   wire n8169;
   wire n8170;
   wire n8171;
   wire n8172;
   wire n8173;
   wire n8174;
   wire n8175;
   wire n8176;
   wire n8177;
   wire n8178;
   wire n8179;
   wire n8180;
   wire n8181;
   wire n8182;
   wire n8183;
   wire n8184;
   wire n8185;
   wire n8186;
   wire n8187;
   wire n8188;
   wire n8189;
   wire n8190;
   wire n8191;
   wire n8192;
   wire n8193;
   wire n8194;
   wire n8195;
   wire n8196;
   wire n8197;
   wire n8198;
   wire n8199;
   wire n8200;
   wire n8201;
   wire n8202;
   wire n8203;
   wire n8204;
   wire n8205;
   wire n8206;
   wire n8207;
   wire n8208;
   wire n8209;
   wire n8210;
   wire n8211;
   wire n8212;
   wire n8213;
   wire n8214;
   wire n8215;
   wire n8216;
   wire n8217;
   wire n8218;
   wire n8219;
   wire n8220;
   wire n8221;
   wire n8222;
   wire n8223;
   wire n8224;
   wire n8225;
   wire n8226;
   wire n8227;
   wire n8228;
   wire n8229;
   wire n8230;
   wire n8231;
   wire n8232;
   wire n8233;
   wire n8234;
   wire n8235;
   wire n8236;
   wire n8237;
   wire n8238;
   wire n8239;
   wire n8240;
   wire n8241;
   wire n8242;
   wire n8243;
   wire n8244;
   wire n8245;
   wire n8246;
   wire n8247;
   wire n8248;
   wire n8249;
   wire n8250;
   wire n8251;
   wire n8252;
   wire n8253;
   wire n8254;
   wire n8255;
   wire n8256;
   wire n8257;
   wire n8258;
   wire n8259;
   wire n8260;
   wire n8261;
   wire n8262;
   wire n8263;
   wire n8264;
   wire n8265;
   wire n8266;
   wire n8267;
   wire n8268;
   wire n8269;
   wire n8270;
   wire n8271;
   wire n8272;
   wire n8273;
   wire n8274;
   wire n8275;
   wire n8276;
   wire n8277;
   wire n8278;
   wire n8279;
   wire n8280;
   wire n8281;
   wire n8282;
   wire n8283;
   wire n8284;
   wire n8285;
   wire n8286;
   wire n8287;
   wire n8288;
   wire n8289;
   wire n8290;
   wire n8291;
   wire n8292;
   wire n8293;
   wire n8294;
   wire n8295;
   wire n8296;
   wire n8297;
   wire n8298;
   wire n8299;
   wire n8300;
   wire n8301;
   wire n8302;
   wire n8303;
   wire n8304;
   wire n8305;
   wire n8306;
   wire n8307;
   wire n8308;
   wire n8309;
   wire n8310;
   wire n8311;
   wire n8312;
   wire n8313;
   wire n8314;
   wire n8315;
   wire n8316;
   wire n8317;
   wire n8318;
   wire n8319;
   wire n8320;
   wire n8321;
   wire n8322;
   wire n8323;
   wire n8324;
   wire n8325;
   wire n8326;
   wire n8327;
   wire n8328;
   wire n8329;
   wire n8330;
   wire n8331;
   wire n8332;
   wire n8333;
   wire n8334;
   wire n8335;
   wire n8336;
   wire n8337;
   wire n8338;
   wire n8339;
   wire n8340;
   wire n8341;
   wire n8342;
   wire n8343;
   wire n8344;
   wire n8345;
   wire n8346;
   wire n8347;
   wire n8348;
   wire n8349;
   wire n8350;
   wire n8351;
   wire n8352;
   wire n8353;
   wire n8354;
   wire n8355;
   wire n8356;
   wire n8357;
   wire n8358;
   wire n8359;
   wire n8360;
   wire n8361;
   wire n8362;
   wire n8363;
   wire n8364;
   wire n8365;
   wire n8366;
   wire n8367;
   wire n8368;
   wire n8369;
   wire n8370;
   wire n8371;
   wire n8372;
   wire n8373;
   wire n8374;
   wire n8375;
   wire n8376;
   wire n8377;
   wire n8378;
   wire n8379;
   wire n8380;
   wire n8381;
   wire n8382;
   wire n8383;
   wire n8384;
   wire n8385;
   wire n8386;
   wire n8387;
   wire n8388;
   wire n8389;
   wire n8390;
   wire n8391;
   wire n8392;
   wire n8393;
   wire n8394;
   wire n8395;
   wire n8396;
   wire n8397;
   wire n8398;
   wire n8399;
   wire n8400;
   wire n8401;
   wire n8402;
   wire n8403;
   wire n8404;
   wire n8405;
   wire n8406;
   wire n8407;
   wire n8408;
   wire n8409;
   wire n8410;
   wire n8411;
   wire n8412;
   wire n8413;
   wire n8414;
   wire n8415;
   wire n8416;
   wire n8417;
   wire n8418;
   wire n8419;
   wire n8420;
   wire n8421;
   wire n8422;
   wire n8423;
   wire n8424;
   wire n8425;
   wire n8426;
   wire n8427;
   wire n8428;
   wire n8429;
   wire n8430;
   wire n8431;
   wire n8432;
   wire n8433;
   wire n8434;
   wire n8435;
   wire n8436;
   wire n8437;
   wire n8438;
   wire n8439;
   wire n8440;
   wire n8441;
   wire n8442;
   wire n8443;
   wire n8444;
   wire n8445;
   wire n8446;
   wire n8447;
   wire n8448;
   wire n8449;
   wire n8450;
   wire n8451;
   wire n8452;
   wire n8453;
   wire n8454;
   wire n8455;
   wire n8456;
   wire n8457;
   wire n8458;
   wire n8459;
   wire n8460;
   wire n8461;
   wire n8462;
   wire n8463;
   wire n8464;
   wire n8465;
   wire n8466;
   wire n8467;
   wire n8468;
   wire n8469;
   wire n8470;
   wire n8471;
   wire n8472;
   wire n8473;
   wire n8474;
   wire n8475;
   wire n8476;
   wire n8477;
   wire n8478;
   wire n8479;
   wire n8480;
   wire n8481;
   wire n8482;
   wire n8483;
   wire n8484;
   wire n8485;
   wire n8486;
   wire n8487;
   wire n8488;
   wire n8489;
   wire n8490;
   wire n8491;
   wire n8492;
   wire n8493;
   wire n8494;
   wire n8495;
   wire n8496;
   wire n8497;
   wire n8498;
   wire n8499;
   wire n8500;
   wire n8501;
   wire n8502;
   wire n8503;
   wire n8504;
   wire n8505;
   wire n8506;
   wire n8507;
   wire n8508;
   wire n8509;
   wire n8510;
   wire n8511;
   wire n8512;
   wire n8513;
   wire n8514;
   wire n8515;
   wire n8516;
   wire n8517;
   wire n8518;
   wire n8519;
   wire n8520;
   wire n8521;
   wire n8522;
   wire n8523;
   wire n8524;
   wire n8525;
   wire n8526;
   wire n8527;
   wire n8528;
   wire n8529;
   wire n8530;
   wire n8531;
   wire n8532;
   wire n8533;
   wire n8534;
   wire n8535;
   wire n8536;
   wire n8537;
   wire n8538;
   wire n8539;
   wire n8540;
   wire n8541;
   wire n8542;
   wire n8543;
   wire n8544;
   wire n8545;
   wire n8546;
   wire n8547;
   wire n8548;
   wire n8549;
   wire n8550;
   wire n8551;
   wire n8552;
   wire n8553;
   wire n8554;
   wire n8555;
   wire n8556;
   wire n8557;
   wire n8558;
   wire n8559;
   wire n8560;
   wire n8561;
   wire n8562;
   wire n8563;
   wire n8564;
   wire n8565;
   wire n8566;
   wire n8567;
   wire n8568;
   wire n8569;
   wire n8570;
   wire n8571;
   wire n8572;
   wire n8573;
   wire n8574;
   wire n8575;
   wire n8576;
   wire n8577;
   wire n8578;
   wire n8579;
   wire n8580;
   wire n8581;
   wire n8582;
   wire n8583;
   wire n8584;
   wire n8585;
   wire n8586;
   wire n8587;
   wire n8588;
   wire n8589;
   wire n8590;
   wire n8591;
   wire n8592;
   wire n8593;
   wire n8594;
   wire n8595;
   wire n8596;
   wire n8597;
   wire n8598;
   wire n8599;
   wire n8600;
   wire n8601;
   wire n8602;
   wire n8603;
   wire n8604;
   wire n8605;
   wire n8606;
   wire n8607;
   wire n8608;
   wire n8609;
   wire n8610;
   wire n8611;
   wire n8612;
   wire n8613;
   wire n8614;
   wire n8615;
   wire n8616;
   wire n8617;
   wire n8618;
   wire n8619;
   wire n8620;
   wire n8621;
   wire n8622;
   wire n8623;
   wire n8624;
   wire n8625;
   wire n8626;
   wire n8627;
   wire n8628;
   wire n8629;
   wire n8630;
   wire n8631;
   wire n8632;
   wire n8633;
   wire n8634;
   wire n8635;
   wire n8636;
   wire n8637;
   wire n8638;
   wire n8639;
   wire n8640;
   wire n8641;
   wire n8642;
   wire n8643;
   wire n8644;
   wire n8645;
   wire n8646;
   wire n8647;
   wire n8648;
   wire n8649;
   wire n8650;
   wire n8651;
   wire n8652;
   wire n8653;
   wire n8654;
   wire n8655;
   wire n8656;
   wire n8657;
   wire n8658;
   wire n8659;
   wire n8660;
   wire n8661;
   wire n8662;
   wire n8663;
   wire n8664;
   wire n8665;
   wire n8666;
   wire n8667;
   wire n8668;
   wire n8669;
   wire n8670;
   wire n8671;
   wire n8672;
   wire n8673;
   wire n8674;
   wire n8675;
   wire n8676;
   wire n8677;
   wire n8678;
   wire n8679;
   wire n8680;
   wire n8681;
   wire n8682;
   wire n8683;
   wire n8684;
   wire n8685;
   wire n8686;
   wire n8687;
   wire n8688;
   wire n8689;
   wire n8690;
   wire n8691;
   wire n8692;
   wire n8693;
   wire n8694;
   wire n8695;
   wire n8696;
   wire n8697;
   wire n8698;
   wire n8699;
   wire n8700;
   wire n8701;
   wire n8702;
   wire n8703;
   wire n8704;
   wire n8705;
   wire n8706;
   wire n8707;
   wire n8708;
   wire n8709;
   wire n8710;
   wire n8711;
   wire n8712;
   wire n8713;
   wire n8714;
   wire n8715;
   wire n8716;
   wire n8717;
   wire n8718;
   wire n8719;
   wire n8720;
   wire n8721;
   wire n8722;
   wire n8723;
   wire n8724;
   wire n8725;
   wire n8726;
   wire n8727;
   wire n8728;
   wire n8729;
   wire n8730;
   wire n8731;
   wire n8732;
   wire n8733;
   wire n8734;
   wire n8735;
   wire n8736;
   wire n8737;
   wire n8738;
   wire n8739;
   wire n8740;
   wire n8741;
   wire n8742;
   wire n8743;
   wire n8744;
   wire n8745;
   wire n8746;
   wire n8747;
   wire n8748;
   wire n8749;
   wire n8750;
   wire n8751;
   wire n8752;
   wire n8753;
   wire n8754;
   wire n8755;
   wire n8756;
   wire n8757;
   wire n8758;
   wire n8759;
   wire n8760;
   wire n8761;
   wire n8762;
   wire n8763;
   wire n8764;
   wire n8765;
   wire n8766;
   wire n8767;
   wire n8768;
   wire n8769;
   wire n8770;
   wire n8771;
   wire n8772;
   wire n8773;
   wire n8774;
   wire n8775;
   wire n8776;
   wire n8777;
   wire n8778;
   wire n8779;
   wire n8780;
   wire n8781;
   wire n8782;
   wire n8783;
   wire n8784;
   wire n8785;
   wire n8786;
   wire n8787;
   wire n8788;
   wire n8789;
   wire n8790;
   wire n8791;
   wire n8792;
   wire n8793;
   wire n8794;
   wire n8795;
   wire n8796;
   wire n8797;
   wire n8798;
   wire n8799;
   wire n8800;
   wire n8801;
   wire n8802;
   wire n8803;
   wire n8804;
   wire n8805;
   wire n8806;
   wire n8807;
   wire n8808;
   wire n8809;
   wire n8810;
   wire n8811;
   wire n8812;
   wire n8813;
   wire n8814;
   wire n8815;
   wire n8816;
   wire n8817;
   wire n8818;
   wire n8819;
   wire n8820;
   wire n8821;
   wire n8822;
   wire n8823;
   wire n8824;
   wire n8825;
   wire n8826;
   wire n8827;
   wire n8828;
   wire n8829;
   wire n8830;
   wire n8831;
   wire n8832;
   wire n8833;
   wire n8834;
   wire n8835;
   wire n8836;
   wire n8837;
   wire n8838;
   wire n8839;
   wire n8840;
   wire n8841;
   wire n8842;
   wire n8843;
   wire n8844;
   wire n8845;
   wire n8846;
   wire n8847;
   wire n8848;
   wire n8849;
   wire n8850;
   wire n8851;
   wire n8852;
   wire n8853;
   wire n8854;
   wire n8855;
   wire n8856;
   wire n8857;
   wire n8858;
   wire n8859;
   wire n8860;
   wire n8861;
   wire n8862;
   wire n8863;
   wire n8864;
   wire n8865;
   wire n8866;
   wire n8867;
   wire n8868;
   wire n8869;
   wire n8870;
   wire n8871;
   wire n8872;
   wire n8873;
   wire n8874;
   wire n8875;
   wire n8876;
   wire n8877;
   wire n8878;
   wire n8879;
   wire n8880;
   wire n8881;
   wire n8882;
   wire n8883;
   wire n8884;
   wire n8885;
   wire n8886;
   wire n8887;
   wire n8888;
   wire n8889;
   wire n8890;
   wire n8891;
   wire n8892;
   wire n8893;
   wire n8894;
   wire n8895;
   wire n8896;
   wire n8897;
   wire n8898;
   wire n8899;
   wire n8900;
   wire n8901;
   wire n8902;
   wire n8903;
   wire n8904;
   wire n8905;
   wire n8906;
   wire n8907;
   wire n8908;
   wire n8909;
   wire n8910;
   wire n8911;
   wire n8912;
   wire n8913;
   wire n8914;
   wire n8915;
   wire n8916;
   wire n8917;
   wire n8918;
   wire n8919;
   wire n8920;
   wire n8921;
   wire n8922;
   wire n8923;
   wire n8924;
   wire n8925;
   wire n8926;
   wire n8927;
   wire n8928;
   wire n8929;
   wire n8930;
   wire n8931;
   wire n8932;
   wire n8933;
   wire n8934;
   wire n8935;
   wire n8936;
   wire n8937;
   wire n8938;
   wire n8939;
   wire n8940;
   wire n8941;
   wire n8942;
   wire n8943;
   wire n8944;
   wire n8945;
   wire n8946;
   wire n8947;
   wire n8948;
   wire n8949;
   wire n8950;
   wire n8951;
   wire n8952;
   wire n8953;
   wire n8954;
   wire n8955;
   wire n8956;
   wire n8957;
   wire n8958;
   wire n8959;
   wire n8960;
   wire n8961;
   wire n8962;
   wire n8963;
   wire n8964;
   wire n8965;
   wire n8966;
   wire n8967;
   wire n8968;
   wire n8969;
   wire n8970;
   wire n8971;
   wire n8972;
   wire n8973;
   wire n8974;
   wire n8975;
   wire n8976;
   wire n8977;
   wire n8978;
   wire n8979;
   wire n8980;
   wire n8981;
   wire n8982;
   wire n8983;
   wire n8984;
   wire n8985;
   wire n8986;
   wire n8987;
   wire n8988;
   wire n8989;
   wire n8990;
   wire n8991;
   wire n8992;
   wire n8993;
   wire n8994;
   wire n8995;
   wire n8996;
   wire n8997;
   wire n8998;
   wire n8999;
   wire n9000;
   wire n9001;
   wire n9002;
   wire n9003;
   wire n9004;
   wire n9005;
   wire n9006;
   wire n9007;
   wire n9008;
   wire n9009;
   wire n9010;
   wire n9011;
   wire n9012;
   wire n9013;
   wire n9014;
   wire n9015;
   wire n9016;
   wire n9017;
   wire n9018;
   wire n9019;
   wire n9020;
   wire n9021;
   wire n9022;
   wire n9023;
   wire n9024;
   wire n9025;
   wire n9026;
   wire n9027;
   wire n9028;
   wire n9029;
   wire n9030;
   wire n9031;
   wire n9032;
   wire n9033;
   wire n9034;
   wire n9035;
   wire n9036;
   wire n9037;
   wire n9038;
   wire n9039;
   wire n9040;
   wire n9041;
   wire n9042;
   wire n9043;
   wire n9044;
   wire n9045;
   wire n9046;
   wire n9047;
   wire n9048;
   wire n9049;
   wire n9050;
   wire n9051;
   wire n9052;
   wire n9053;
   wire n9054;
   wire n9055;
   wire n9056;
   wire n9057;
   wire n9058;
   wire n9059;
   wire n9060;
   wire n9061;
   wire n9062;
   wire n9063;
   wire n9064;
   wire n9065;
   wire n9066;
   wire n9067;
   wire n9068;
   wire n9069;
   wire n9070;
   wire n9071;
   wire n9072;
   wire n9073;
   wire n9074;
   wire n9075;
   wire n9076;
   wire n9077;
   wire n9078;
   wire n9079;
   wire n9080;
   wire n9081;
   wire n9082;
   wire n9083;
   wire n9084;
   wire n9085;
   wire n9086;
   wire n9087;
   wire n9088;
   wire n9089;
   wire n9090;
   wire n9091;
   wire n9092;
   wire n9093;
   wire n9094;
   wire n9095;
   wire n9096;
   wire n9097;
   wire n9098;
   wire n9099;
   wire n9100;
   wire n9101;
   wire n9102;
   wire n9103;
   wire n9104;
   wire n9105;
   wire n9106;
   wire n9107;
   wire n9108;
   wire n9109;
   wire n9110;
   wire n9111;
   wire n9112;
   wire n9113;
   wire n9114;
   wire n9115;
   wire n9116;
   wire n9117;
   wire n9118;
   wire n9119;
   wire n9120;
   wire n9121;
   wire n9122;
   wire n9123;
   wire n9124;
   wire n9125;
   wire n9126;
   wire n9127;
   wire n9128;
   wire n9129;
   wire n9130;
   wire n9131;
   wire n9132;
   wire n9133;
   wire n9134;
   wire n9135;
   wire n9136;
   wire n9137;
   wire n9138;
   wire n9139;
   wire n9140;
   wire n9141;
   wire n9142;
   wire n9143;
   wire n9144;
   wire n9145;
   wire n9146;
   wire n9147;
   wire n9148;
   wire n9149;
   wire n9150;
   wire n9151;
   wire n9152;
   wire n9153;
   wire n9154;
   wire n9155;
   wire n9156;
   wire n9157;
   wire n9158;
   wire n9159;
   wire n9160;
   wire n9161;
   wire n9162;
   wire n9163;
   wire n9164;
   wire n9165;
   wire n9166;
   wire n9167;
   wire n9168;
   wire n9169;
   wire n9170;
   wire n9171;
   wire n9172;
   wire n9173;
   wire n9174;
   wire n9175;
   wire n9176;
   wire n9177;
   wire n9178;
   wire n9179;
   wire n9180;
   wire n9181;
   wire n9182;
   wire n9183;
   wire n9184;
   wire n9185;
   wire n9186;
   wire n9187;
   wire n9188;
   wire n9189;
   wire n9190;
   wire n9191;
   wire n9192;
   wire n9193;
   wire n9194;
   wire n9195;
   wire n9196;
   wire n9197;
   wire n9198;
   wire n9199;
   wire n9200;
   wire n9201;
   wire n9202;
   wire n9203;
   wire n9204;
   wire n9205;
   wire n9206;
   wire n9207;
   wire n9208;
   wire n9209;
   wire n9210;
   wire n9211;
   wire n9212;
   wire n9213;
   wire n9214;
   wire n9215;
   wire n9216;
   wire n9217;
   wire n9218;
   wire n9219;
   wire n9220;
   wire n9221;
   wire n9222;
   wire n9223;
   wire n9224;
   wire n9225;
   wire n9226;
   wire n9227;
   wire n9228;
   wire n9229;
   wire n9230;
   wire n9231;
   wire n9232;
   wire n9233;
   wire n9234;
   wire n9235;
   wire n9236;
   wire n9237;
   wire n9238;
   wire n9239;
   wire n9240;
   wire n9241;
   wire n9242;
   wire n9243;
   wire n9244;
   wire n9245;
   wire n9246;
   wire n9247;
   wire n9248;
   wire n9249;
   wire n9250;
   wire n9251;
   wire n9252;
   wire n9253;
   wire n9254;
   wire n9255;
   wire n9256;
   wire n9257;
   wire n9258;
   wire n9259;
   wire n9260;
   wire n9261;
   wire n9262;
   wire n9263;
   wire n9264;
   wire n9265;
   wire n9266;
   wire n9267;
   wire n9268;
   wire n9269;
   wire n9270;
   wire n9271;
   wire n9272;
   wire n9273;
   wire n9274;
   wire n9275;
   wire n9276;
   wire n9277;
   wire n9278;
   wire n9279;
   wire n9280;
   wire n9281;
   wire n9282;
   wire n9283;
   wire n9284;
   wire n9285;
   wire n9286;
   wire n9287;
   wire n9288;
   wire n9289;
   wire n9290;
   wire n9291;
   wire n9292;
   wire n9293;
   wire n9294;
   wire n9295;
   wire n9296;
   wire n9297;
   wire n9298;
   wire n9299;
   wire n9300;
   wire n9301;
   wire n9302;
   wire n9303;
   wire n9304;
   wire n9305;
   wire n9306;
   wire n9307;
   wire n9308;
   wire n9309;
   wire n9310;
   wire n9311;
   wire n9312;
   wire n9313;
   wire n9314;
   wire n9315;
   wire n9316;
   wire n9317;
   wire n9318;
   wire n9319;
   wire n9320;
   wire n9321;
   wire n9322;
   wire n9323;
   wire n9324;
   wire n9325;
   wire n9326;
   wire n9327;
   wire n9328;
   wire n9329;
   wire n9330;
   wire n9331;
   wire n9332;
   wire n9333;
   wire n9334;
   wire n9335;
   wire n9336;
   wire n9337;
   wire n9338;
   wire n9339;
   wire n9340;
   wire n9341;
   wire n9342;
   wire n9343;
   wire n9344;
   wire n9345;
   wire n9346;
   wire n9347;
   wire n9348;
   wire n9349;
   wire n9350;
   wire n9351;
   wire n9352;
   wire n9353;
   wire n9354;
   wire n9355;
   wire n9356;
   wire n9357;
   wire n9358;
   wire n9359;
   wire n9360;
   wire n9361;
   wire n9362;
   wire n9363;
   wire n9364;
   wire n9365;
   wire n9366;
   wire n9367;
   wire n9368;
   wire n9369;
   wire n9370;
   wire n9371;
   wire n9372;
   wire n9373;
   wire n9374;
   wire n9375;
   wire n9376;
   wire n9377;
   wire n9378;
   wire n9379;
   wire n9380;
   wire n9381;
   wire n9382;
   wire n9383;
   wire n9384;
   wire n9385;
   wire n9386;
   wire n9387;
   wire n9388;
   wire n9389;
   wire n9390;
   wire n9391;
   wire n9392;
   wire n9393;
   wire n9394;
   wire n9395;
   wire n9396;
   wire n9397;
   wire n9398;
   wire n9399;
   wire n9400;
   wire n9401;
   wire n9402;
   wire n9403;
   wire n9404;
   wire n9405;
   wire n9406;
   wire n9407;
   wire n9408;
   wire n9409;
   wire n9410;
   wire n9411;
   wire n9412;
   wire n9413;
   wire n9414;
   wire n9415;
   wire n9416;
   wire n9417;
   wire n9418;
   wire n9419;
   wire n9420;
   wire n9421;
   wire n9422;
   wire n9423;
   wire n9424;
   wire n9425;
   wire n9426;
   wire n9427;
   wire n9428;
   wire n9429;
   wire n9430;
   wire n9431;
   wire n9432;
   wire n9433;
   wire n9434;
   wire n9435;
   wire n9436;
   wire n9437;
   wire n9438;
   wire n9439;
   wire n9440;
   wire n9441;
   wire n9442;
   wire n9443;
   wire n9444;
   wire n9445;
   wire n9446;
   wire n9447;
   wire n9448;
   wire n9449;
   wire n9450;
   wire n9451;
   wire n9452;
   wire n9453;
   wire n9454;
   wire n9455;
   wire n9456;
   wire n9457;
   wire n9458;
   wire n9459;
   wire n9460;
   wire n9461;
   wire n9462;
   wire n9463;
   wire n9464;
   wire n9465;
   wire n9466;
   wire n9467;
   wire n9468;
   wire n9469;
   wire n9470;
   wire n9471;
   wire n9472;
   wire n9473;
   wire n9474;
   wire n9475;
   wire n9476;
   wire n9477;
   wire n9478;
   wire n9479;
   wire n9480;
   wire n9481;
   wire n9482;
   wire n9483;
   wire n9484;
   wire n9485;
   wire n9486;
   wire n9487;
   wire n9488;
   wire n9489;
   wire n9490;
   wire n9491;
   wire n9492;
   wire n9493;
   wire n9494;
   wire n9495;
   wire n9496;
   wire n9497;
   wire n9498;
   wire n9499;
   wire n9500;
   wire n9501;
   wire n9502;
   wire n9503;
   wire n9504;
   wire n9505;
   wire n9506;
   wire n9507;
   wire n9508;
   wire n9509;
   wire n9510;
   wire n9511;
   wire n9512;
   wire n9513;
   wire n9514;
   wire n9515;
   wire n9516;
   wire n9517;
   wire n9518;
   wire n9519;
   wire n9520;
   wire n9521;
   wire n9522;
   wire n9523;
   wire n9524;
   wire n9525;
   wire n9526;
   wire n9527;
   wire n9528;
   wire n9529;
   wire n9530;
   wire n9531;
   wire n9532;
   wire n9533;
   wire n9534;
   wire n9535;
   wire n9536;
   wire n9537;
   wire n9538;
   wire n9539;
   wire n9540;
   wire n9541;
   wire n9542;
   wire n9543;
   wire n9544;
   wire n9545;
   wire n9546;
   wire n9547;
   wire n9548;
   wire n9549;
   wire n9550;
   wire n9551;
   wire n9552;
   wire n9553;
   wire n9554;
   wire n9555;
   wire n9556;
   wire n9557;
   wire n9558;
   wire n9559;
   wire n9560;
   wire n9561;
   wire n9562;
   wire n9563;
   wire n9564;
   wire n9565;
   wire n9566;
   wire n9567;
   wire n9568;
   wire n9569;
   wire n9570;
   wire n9571;
   wire n9572;
   wire n9573;
   wire n9574;
   wire n9575;
   wire n9576;
   wire n9577;
   wire n9578;
   wire n9579;
   wire n9580;
   wire n9581;
   wire n9582;
   wire n9583;
   wire n9584;
   wire n9585;
   wire n9586;
   wire n9587;
   wire n9588;
   wire n9589;
   wire n9590;
   wire n9591;
   wire n9592;
   wire n9593;
   wire n9594;
   wire n9595;
   wire n9596;
   wire n9597;
   wire n9598;
   wire n9599;
   wire n9600;
   wire n9601;
   wire n9602;
   wire n9603;
   wire n9604;
   wire n9605;
   wire n9606;
   wire n9607;
   wire n9608;
   wire n9609;
   wire n9610;
   wire n9611;
   wire n9612;
   wire n9613;
   wire n9614;
   wire n9615;
   wire n9616;
   wire n9617;
   wire n9618;
   wire n9619;
   wire n9620;
   wire n9621;
   wire n9622;
   wire n9623;
   wire n9624;
   wire n9625;
   wire n9626;
   wire n9627;
   wire n9628;
   wire n9629;
   wire n9630;
   wire n9631;
   wire n9632;
   wire n9633;
   wire n9634;
   wire n9635;
   wire n9636;
   wire n9637;
   wire n9638;
   wire n9639;
   wire n9640;
   wire n9641;
   wire n9642;
   wire n9643;
   wire n9644;
   wire n9645;
   wire n9646;
   wire n9647;
   wire n9648;
   wire n9649;
   wire n9650;
   wire n9651;
   wire n9652;
   wire n9653;
   wire n9654;
   wire n9655;
   wire n9656;
   wire n9657;
   wire n9658;
   wire n9659;
   wire n9660;
   wire n9661;
   wire n9662;
   wire n9663;
   wire n9664;
   wire n9665;
   wire n9666;
   wire n9667;
   wire n9668;
   wire n9669;
   wire n9670;
   wire n9671;
   wire n9672;
   wire n9673;
   wire n9674;
   wire n9675;
   wire n9676;
   wire n9677;
   wire n9678;
   wire n9679;
   wire n9680;
   wire n9681;
   wire n9682;
   wire n9683;
   wire n9684;
   wire n9685;
   wire n9686;
   wire n9687;
   wire n9688;
   wire n9689;
   wire n9690;
   wire n9691;
   wire n9692;
   wire n9693;
   wire n9694;
   wire n9695;
   wire n9696;
   wire n9697;
   wire n9698;
   wire n9699;
   wire n9700;
   wire n9701;
   wire n9702;
   wire n9703;
   wire n9704;
   wire n9705;
   wire n9706;
   wire n9707;
   wire n9708;
   wire n9709;
   wire n9710;
   wire n9711;
   wire n9712;
   wire n9713;
   wire n9714;
   wire n9715;
   wire n9716;
   wire n9717;
   wire n9718;
   wire n9719;
   wire n9720;
   wire n9721;
   wire n9722;
   wire n9723;
   wire n9724;
   wire n9725;
   wire n9726;
   wire n9727;
   wire n9728;
   wire n9729;
   wire n9730;
   wire n9731;
   wire n9732;
   wire n9733;
   wire n9734;
   wire n9735;
   wire n9736;
   wire n9737;
   wire n9738;
   wire n9739;
   wire n9740;
   wire n9741;
   wire n9742;
   wire n9743;
   wire n9744;
   wire n9745;
   wire n9746;
   wire n9747;
   wire n9748;
   wire n9749;
   wire n9750;
   wire n9751;
   wire n9752;
   wire n9753;
   wire n9754;
   wire n9755;
   wire n9756;
   wire n9757;
   wire n9758;
   wire n9759;
   wire n9760;
   wire n9761;
   wire n9762;
   wire n9763;
   wire n9764;
   wire n9765;
   wire n9766;
   wire n9767;
   wire n9768;
   wire n9769;
   wire n9770;
   wire n9771;
   wire n9772;
   wire n9773;
   wire n9774;
   wire n9775;
   wire n9776;
   wire n9777;
   wire n9778;
   wire n9779;
   wire n9780;
   wire n9781;
   wire n9782;
   wire n9783;
   wire n9784;
   wire n9785;
   wire n9786;
   wire n9787;
   wire n9788;
   wire n9789;
   wire n9790;
   wire n9791;
   wire n9792;
   wire n9793;
   wire n9794;
   wire n9795;
   wire n9796;
   wire n9797;
   wire n9798;
   wire n9799;
   wire n9800;
   wire n9801;
   wire n9802;
   wire n9803;
   wire n9804;
   wire n9805;
   wire n9806;
   wire n9807;
   wire n9808;
   wire n9809;
   wire n9810;
   wire n9811;
   wire n9812;
   wire n9813;
   wire n9814;
   wire n9815;
   wire n9816;
   wire n9817;
   wire n9818;
   wire n9819;
   wire n9820;
   wire n9821;
   wire n9822;
   wire n9823;
   wire n9824;
   wire n9825;
   wire n9826;
   wire n9827;
   wire n9828;
   wire n9829;
   wire n9830;
   wire n9831;
   wire n9832;
   wire n9833;
   wire n9834;
   wire n9835;
   wire n9836;
   wire n9837;
   wire n9838;
   wire n9839;
   wire n9840;
   wire n9841;
   wire n9842;
   wire n9843;
   wire n9844;
   wire n9845;
   wire n9846;
   wire n9847;
   wire n9848;
   wire n9849;
   wire n9850;
   wire n9851;
   wire n9852;
   wire n9853;
   wire n9854;
   wire n9855;
   wire n9856;
   wire n9857;
   wire n9858;
   wire n9859;
   wire n9860;
   wire n9861;
   wire n9862;
   wire n9863;
   wire n9864;
   wire n9865;
   wire n9866;
   wire n9867;
   wire n9868;
   wire n9869;
   wire n9870;
   wire n9871;
   wire n9872;
   wire n9873;
   wire n9874;
   wire n9875;
   wire n9876;
   wire n9877;
   wire n9878;
   wire n9879;
   wire n9880;
   wire n9881;
   wire n9882;
   wire n9883;
   wire n9884;
   wire n9885;
   wire n9886;
   wire n9887;
   wire n9888;
   wire n9889;
   wire n9890;
   wire n9891;
   wire n9892;
   wire n9893;
   wire n9894;
   wire n9895;
   wire n9896;
   wire n9897;
   wire n9898;
   wire n9899;
   wire n9900;
   wire n9901;
   wire n9902;
   wire n9903;
   wire n9904;
   wire n9905;
   wire n9906;
   wire n9907;
   wire n9908;
   wire n9909;
   wire n9910;
   wire n9911;
   wire n9912;
   wire n9913;
   wire n9914;
   wire n9915;
   wire n9916;
   wire n9917;
   wire n9918;
   wire n9919;
   wire n9920;
   wire n9921;
   wire n9922;
   wire n9923;
   wire n9924;
   wire n9925;
   wire n9926;
   wire n9927;
   wire n9928;
   wire n9929;
   wire n9930;
   wire n9931;
   wire n9932;
   wire n9933;
   wire n9934;
   wire n9935;
   wire n9936;
   wire n9937;
   wire n9938;
   wire n9939;
   wire n9940;
   wire n9941;
   wire n9942;
   wire n9943;
   wire n9944;
   wire n9945;
   wire n9946;
   wire n9947;
   wire n9948;
   wire n9949;
   wire n9950;
   wire n9951;
   wire n9952;
   wire n9953;
   wire n9954;
   wire n9955;
   wire n9956;
   wire n9957;
   wire n9958;
   wire n9959;
   wire n9960;
   wire n9961;
   wire n9962;
   wire n9963;
   wire n9964;
   wire n9965;
   wire n9966;
   wire n9967;
   wire n9968;
   wire n9969;
   wire n9970;
   wire n9971;
   wire n9972;
   wire n9973;
   wire n9974;
   wire n9975;
   wire n9976;
   wire n9977;
   wire n9978;
   wire n9979;
   wire n9980;
   wire n9981;
   wire n9982;
   wire n9983;
   wire n9984;
   wire n9985;
   wire n9986;
   wire n9987;
   wire n9988;
   wire n9989;
   wire n9990;
   wire n9991;
   wire n9992;
   wire n9993;
   wire n9994;
   wire n9995;
   wire n9996;
   wire n9997;
   wire n9998;
   wire n9999;
   wire n10000;
   wire n10001;
   wire n10002;
   wire n10003;
   wire n10004;
   wire n10005;
   wire n10006;
   wire n10007;
   wire n10008;
   wire n10009;
   wire n10010;
   wire n10011;
   wire n10012;
   wire n10013;
   wire n10014;
   wire n10015;
   wire n10016;
   wire n10017;
   wire n10018;
   wire n10019;
   wire n10020;
   wire n10021;
   wire n10022;
   wire n10023;
   wire n10024;
   wire n10025;
   wire n10026;
   wire n10027;
   wire n10028;
   wire n10029;
   wire n10030;
   wire n10031;
   wire n10032;
   wire n10033;
   wire n10034;
   wire n10035;
   wire n10036;
   wire n10037;
   wire n10038;
   wire n10039;
   wire n10040;
   wire n10041;
   wire n10042;
   wire n10043;
   wire n10044;
   wire n10045;
   wire n10046;
   wire n10047;
   wire n10048;
   wire n10049;
   wire n10050;
   wire n10051;
   wire n10052;
   wire n10053;
   wire n10054;
   wire n10055;
   wire n10056;
   wire n10057;
   wire n10058;
   wire n10059;
   wire n10060;
   wire n10061;
   wire n10062;
   wire n10063;
   wire n10064;
   wire n10065;
   wire n10066;
   wire n10067;
   wire n10068;
   wire n10069;
   wire n10070;
   wire n10071;
   wire n10072;
   wire n10073;
   wire n10074;
   wire n10075;
   wire n10076;
   wire n10077;
   wire n10078;
   wire n10079;
   wire n10080;
   wire n10081;
   wire n10082;
   wire n10083;
   wire n10084;
   wire n10085;
   wire n10086;
   wire n10087;
   wire n10088;
   wire n10089;
   wire n10090;
   wire n10091;
   wire n10092;
   wire n10093;
   wire n10094;
   wire n10095;
   wire n10096;
   wire n10097;
   wire n10098;
   wire n10099;
   wire n10100;
   wire n10101;
   wire n10102;
   wire n10103;
   wire n10104;
   wire n10105;
   wire n10106;
   wire n10107;
   wire n10108;
   wire n10109;
   wire n10110;
   wire n10111;
   wire n10112;
   wire n10113;
   wire n10114;
   wire n10115;
   wire n10116;
   wire n10117;
   wire n10118;
   wire n10119;
   wire n10120;
   wire n10121;
   wire n10122;
   wire n10123;
   wire n10124;
   wire n10125;
   wire n10126;
   wire n10127;
   wire n10128;
   wire n10129;
   wire n10130;
   wire n10131;
   wire n10132;
   wire n10133;
   wire n10134;
   wire n10135;
   wire n10136;
   wire n10137;
   wire n10138;
   wire n10139;
   wire n10140;
   wire n10141;
   wire n10142;
   wire n10143;
   wire n10144;
   wire n10145;
   wire n10146;
   wire n10147;
   wire n10148;
   wire n10149;
   wire n10150;
   wire n10151;
   wire n10152;
   wire n10153;
   wire n10154;
   wire n10155;
   wire n10156;
   wire n10157;
   wire n10158;
   wire n10159;
   wire n10160;
   wire n10161;
   wire n10162;
   wire n10163;
   wire n10164;
   wire n10165;
   wire n10166;
   wire n10167;
   wire n10168;
   wire n10169;
   wire n10170;
   wire n10171;
   wire n10172;
   wire n10173;
   wire n10174;
   wire n10175;
   wire n10176;
   wire n10177;
   wire n10178;
   wire n10179;
   wire n10180;
   wire n10181;
   wire n10182;
   wire n10183;
   wire n10184;
   wire n10185;
   wire n10186;
   wire n10187;
   wire n10188;
   wire n10189;
   wire n10190;
   wire n10191;
   wire n10192;
   wire n10193;
   wire n10194;
   wire n10195;
   wire n10196;
   wire n10197;
   wire n10198;
   wire n10199;
   wire n10200;
   wire n10201;
   wire n10202;
   wire n10203;
   wire n10204;
   wire n10205;
   wire n10206;
   wire n10207;
   wire n10208;
   wire n10209;
   wire n10210;
   wire n10211;
   wire n10212;
   wire n10213;
   wire n10214;
   wire n10215;
   wire n10216;
   wire n10217;
   wire n10218;
   wire n10219;
   wire n10220;
   wire n10221;
   wire n10222;
   wire n10223;
   wire n10224;
   wire n10225;
   wire n10226;
   wire n10227;
   wire n10228;
   wire n10229;
   wire n10230;
   wire n10231;
   wire n10232;
   wire n10233;
   wire n10234;
   wire n10235;
   wire n10236;
   wire n10237;
   wire n10238;
   wire n10239;
   wire n10240;
   wire n10241;
   wire n10242;
   wire n10243;
   wire n10244;
   wire n10245;
   wire n10246;
   wire n10247;
   wire n10248;
   wire n10249;
   wire n10250;
   wire n10251;
   wire n10252;
   wire n10253;
   wire n10254;
   wire n10255;
   wire n10256;
   wire n10257;
   wire n10258;
   wire n10259;
   wire n10260;
   wire n10261;
   wire n10262;
   wire n10263;
   wire n10264;
   wire n10265;
   wire n10266;
   wire n10267;
   wire n10268;
   wire n10269;
   wire n10270;
   wire n10271;
   wire n10272;
   wire n10273;
   wire n10274;
   wire n10275;
   wire n10276;
   wire n10277;
   wire n10278;
   wire n10279;
   wire n10280;
   wire n10281;
   wire n10282;
   wire n10283;
   wire n10284;
   wire n10285;
   wire n10286;
   wire n10287;
   wire n10288;
   wire n10289;
   wire n10290;
   wire n10291;
   wire n10292;
   wire n10293;
   wire n10294;
   wire n10295;
   wire n10296;
   wire n10297;
   wire n10298;
   wire n10299;
   wire n10300;
   wire n10301;
   wire n10302;
   wire n10303;
   wire n10304;
   wire n10305;
   wire n10306;
   wire n10307;
   wire n10308;
   wire n10309;
   wire n10310;
   wire n10311;
   wire n10312;
   wire n10313;
   wire n10314;
   wire n10315;
   wire n10316;
   wire n10317;
   wire n10318;
   wire n10319;
   wire n10320;
   wire n10321;
   wire n10322;
   wire n10323;
   wire n10324;
   wire n10325;
   wire n10326;
   wire n10327;
   wire n10328;
   wire n10329;
   wire n10330;
   wire n10331;
   wire n10332;
   wire n10333;
   wire n10334;
   wire n10335;
   wire n10336;
   wire n10337;
   wire n10338;
   wire n10339;
   wire n10340;
   wire n10341;
   wire n10342;
   wire n10343;
   wire n10344;
   wire n10345;
   wire n10346;
   wire n10347;
   wire n10348;
   wire n10349;
   wire n10350;
   wire n10351;
   wire n10352;
   wire n10353;
   wire n10354;
   wire n10355;
   wire n10356;
   wire n10357;
   wire n10358;
   wire n10359;
   wire n10360;
   wire n10361;
   wire n10362;
   wire n10363;
   wire n10364;
   wire n10365;
   wire n10366;
   wire n10367;
   wire n10368;
   wire n10369;
   wire n10370;
   wire n10371;
   wire n10372;
   wire n10373;
   wire n10374;
   wire n10375;
   wire n10376;
   wire n10377;
   wire n10378;
   wire n10379;
   wire n10380;
   wire n10381;
   wire n10382;
   wire n10383;
   wire n10384;
   wire n10385;
   wire n10386;
   wire n10387;
   wire n10388;
   wire n10389;
   wire n10390;
   wire n10391;
   wire n10392;
   wire n10393;
   wire n10394;
   wire n10395;
   wire n10396;
   wire n10397;
   wire n10398;
   wire n10399;
   wire n10400;
   wire n10401;
   wire n10402;
   wire n10403;
   wire n10404;
   wire n10405;
   wire n10406;
   wire n10407;
   wire n10408;
   wire n10409;
   wire n10410;
   wire n10411;
   wire n10412;
   wire n10413;
   wire n10414;
   wire n10415;
   wire n10416;
   wire n10417;
   wire n10418;
   wire n10419;
   wire n10420;
   wire n10421;
   wire n10422;
   wire n10423;
   wire n10424;
   wire n10425;
   wire n10426;
   wire n10427;
   wire n10428;
   wire n10429;
   wire n10430;
   wire n10431;
   wire n10432;
   wire n10433;
   wire n10434;
   wire n10435;
   wire n10436;
   wire n10437;
   wire n10438;
   wire n10439;
   wire n10440;
   wire n10441;
   wire n10442;
   wire n10443;
   wire n10444;
   wire n10445;
   wire n10446;
   wire n10447;
   wire n10448;
   wire n10449;
   wire n10450;
   wire n10451;
   wire n10452;
   wire n10453;
   wire n10454;
   wire n10455;
   wire n10456;
   wire n10457;
   wire n10458;
   wire n10459;
   wire n10460;
   wire n10461;
   wire n10462;
   wire n10463;
   wire n10464;
   wire n10465;
   wire n10466;
   wire n10467;
   wire n10468;
   wire n10469;
   wire n10470;
   wire n10471;
   wire n10472;
   wire n10473;
   wire n10474;
   wire n10475;
   wire n10476;
   wire n10477;
   wire n10478;
   wire n10479;
   wire n10480;
   wire n10481;
   wire n10482;
   wire n10483;
   wire n10484;
   wire n10485;
   wire n10486;
   wire n10487;
   wire n10488;
   wire n10489;
   wire n10490;
   wire n10491;
   wire n10492;
   wire n10493;
   wire n10494;
   wire n10495;
   wire n10496;
   wire n10497;
   wire n10498;
   wire n10499;
   wire n10500;
   wire n10501;
   wire n10502;
   wire n10503;
   wire n10504;
   wire n10505;
   wire n10506;
   wire n10507;
   wire n10508;
   wire n10509;
   wire n10510;
   wire n10511;
   wire n10512;
   wire n10513;
   wire n10514;
   wire n10515;
   wire n10516;
   wire n10517;
   wire n10518;
   wire n10519;
   wire n10520;
   wire n10521;
   wire n10522;
   wire n10523;
   wire n10524;
   wire n10525;
   wire n10526;
   wire n10527;
   wire n10528;
   wire n10529;
   wire n10530;
   wire n10531;
   wire n10532;
   wire n10533;
   wire n10534;
   wire n10535;
   wire n10536;
   wire n10537;
   wire n10538;
   wire n10539;
   wire n10540;
   wire n10541;
   wire n10542;
   wire n10543;
   wire n10544;
   wire n10545;
   wire n10546;
   wire n10547;
   wire n10548;
   wire n10549;
   wire n10550;
   wire n10551;
   wire n10552;
   wire n10553;
   wire n10554;
   wire n10555;
   wire n10556;
   wire n10557;
   wire n10558;
   wire n10559;
   wire n10560;
   wire n10561;
   wire n10562;
   wire n10563;
   wire n10564;
   wire n10565;
   wire n10566;
   wire n10567;
   wire n10568;
   wire n10569;
   wire n10570;
   wire n10571;
   wire n10572;
   wire n10573;
   wire n10574;
   wire n10575;
   wire n10576;
   wire n10577;
   wire n10578;
   wire n10579;
   wire n10580;
   wire n10581;
   wire n10582;
   wire n10583;
   wire n10584;
   wire n10585;
   wire n10586;
   wire n10587;
   wire n10588;
   wire n10589;
   wire n10590;
   wire n10591;
   wire n10592;
   wire n10593;
   wire n10594;
   wire n10595;
   wire n10596;
   wire n10597;
   wire n10598;
   wire n10599;
   wire n10600;
   wire n10601;
   wire n10602;
   wire n10603;
   wire n10604;
   wire n10605;
   wire n10606;
   wire n10607;
   wire n10608;
   wire n10609;
   wire n10610;
   wire n10611;
   wire n10612;
   wire n10613;
   wire n10614;
   wire n10615;
   wire n10616;
   wire n10617;
   wire n10618;
   wire n10619;
   wire n10620;
   wire n10621;
   wire n10622;
   wire n10623;
   wire n10624;
   wire n10625;
   wire n10626;
   wire n10627;
   wire n10628;
   wire n10629;
   wire n10630;
   wire n10631;
   wire n10632;
   wire n10633;
   wire n10634;
   wire n10635;
   wire n10636;
   wire n10637;
   wire n10638;
   wire n10639;
   wire n10640;
   wire n10641;
   wire n10642;
   wire n10643;
   wire n10644;
   wire n10645;
   wire n10646;
   wire n10647;
   wire n10648;
   wire n10649;
   wire n10650;
   wire n10651;
   wire n10652;
   wire n10653;
   wire n10654;
   wire n10655;
   wire n10656;
   wire n10657;
   wire n10658;
   wire n10659;
   wire n10660;
   wire n10661;
   wire n10662;
   wire n10663;
   wire n10664;
   wire n10665;
   wire n10666;
   wire n10667;
   wire n10668;
   wire n10669;
   wire n10670;
   wire n10671;
   wire n10672;
   wire n10673;
   wire n10674;
   wire n10675;
   wire n10676;
   wire n10677;
   wire n10678;
   wire n10679;
   wire n10680;
   wire n10681;
   wire n10682;
   wire n10683;
   wire n10684;
   wire n10685;
   wire n10686;
   wire n10687;
   wire n10688;
   wire n10689;
   wire n10690;
   wire n10691;
   wire n10692;
   wire n10693;
   wire n10694;
   wire n10695;
   wire n10696;
   wire n10697;
   wire n10698;
   wire n10699;
   wire n10700;
   wire n10701;
   wire n10702;
   wire n10703;
   wire n10704;
   wire n10705;
   wire n10706;
   wire n10707;
   wire n10708;
   wire n10709;
   wire n10710;
   wire n10711;
   wire n10712;
   wire n10713;
   wire n10714;
   wire n10715;
   wire n10716;
   wire n10717;
   wire n10718;
   wire n10719;
   wire n10720;
   wire n10721;
   wire n10722;
   wire n10723;
   wire n10724;
   wire n10725;
   wire n10726;
   wire n10727;
   wire n10728;
   wire n10729;
   wire n10730;
   wire n10731;
   wire n10732;
   wire n10733;
   wire n10734;
   wire n10735;
   wire n10736;
   wire n10737;
   wire n10738;
   wire n10739;
   wire n10740;
   wire n10741;
   wire n10742;
   wire n10743;
   wire n10744;
   wire n10745;
   wire n10746;
   wire n10747;
   wire n10748;
   wire n10749;
   wire n10750;
   wire n10751;
   wire n10752;
   wire n10753;
   wire n10754;
   wire n10755;
   wire n10756;
   wire n10757;
   wire n10758;
   wire n10759;
   wire n10760;
   wire n10761;
   wire n10762;
   wire n10763;
   wire n10764;
   wire n10765;
   wire n10766;
   wire n10767;
   wire n10768;
   wire n10769;
   wire n10770;
   wire n10771;
   wire n10772;
   wire n10773;
   wire n10774;
   wire n10775;
   wire n10776;
   wire n10777;
   wire n10778;
   wire n10779;
   wire n10780;
   wire n10781;
   wire n10782;
   wire n10783;
   wire n10784;
   wire n10785;
   wire n10786;
   wire n10787;
   wire n10788;
   wire n10789;
   wire n10790;
   wire n10791;
   wire n10792;
   wire n10793;
   wire n10794;
   wire n10795;
   wire n10796;
   wire n10797;
   wire n10798;
   wire n10799;
   wire n10800;
   wire n10801;
   wire n10802;
   wire n10803;
   wire n10804;
   wire n10805;
   wire n10806;
   wire n10807;
   wire n10808;
   wire n10809;
   wire n10810;
   wire n10811;
   wire n10812;
   wire n10813;
   wire n10814;
   wire n10815;
   wire n10816;
   wire n10817;
   wire n10818;
   wire n10819;
   wire n10820;
   wire n10821;
   wire n10822;
   wire n10823;
   wire n10824;
   wire n10825;
   wire n10826;
   wire n10827;
   wire n10828;
   wire n10829;
   wire n10830;
   wire n10831;
   wire n10832;
   wire n10833;
   wire n10834;
   wire n10835;
   wire n10836;
   wire n10837;
   wire n10838;
   wire n10839;
   wire n10840;
   wire n10841;
   wire n10842;
   wire n10843;
   wire n10844;
   wire n10845;
   wire n10846;
   wire n10847;
   wire n10848;
   wire n10849;
   wire n10850;
   wire n10851;
   wire n10852;
   wire n10853;
   wire n10854;
   wire n10855;
   wire n10856;
   wire n10857;
   wire n10858;
   wire n10859;
   wire n10860;
   wire n10861;
   wire n10862;
   wire n10863;
   wire n10864;
   wire n10865;
   wire n10866;
   wire n10867;
   wire n10868;
   wire n10869;
   wire n10870;
   wire n10871;
   wire n10872;
   wire n10873;
   wire n10874;
   wire n10875;
   wire n10876;
   wire n10877;
   wire n10878;
   wire n10879;
   wire n10880;
   wire n10881;
   wire n10882;
   wire n10883;
   wire n10884;
   wire n10885;
   wire n10886;
   wire n10887;
   wire n10888;
   wire n10889;
   wire n10890;
   wire n10891;
   wire n10892;
   wire n10893;
   wire n10894;
   wire n10895;
   wire n10896;
   wire n10897;
   wire n10898;
   wire n10899;
   wire n10900;
   wire n10901;
   wire n10902;
   wire n10903;
   wire n10904;
   wire n10905;
   wire n10906;
   wire n10907;
   wire n10908;
   wire n10909;
   wire n10910;
   wire n10911;
   wire n10912;
   wire n10913;
   wire n10914;
   wire n10915;
   wire n10916;
   wire n10917;
   wire n10918;
   wire n10919;
   wire n10920;
   wire n10921;
   wire n10922;
   wire n10923;
   wire n10924;
   wire n10925;
   wire n10926;
   wire n10927;
   wire n10928;
   wire n10929;
   wire n10930;
   wire n10931;
   wire n10932;
   wire n10933;
   wire n10934;
   wire n10935;
   wire n10936;
   wire n10937;
   wire n10938;
   wire n10939;
   wire n10940;
   wire n10941;
   wire n10942;
   wire n10943;
   wire n10944;
   wire n10945;
   wire n10946;
   wire n10947;
   wire n10948;
   wire n10949;
   wire n10950;
   wire n10951;
   wire n10952;
   wire n10953;
   wire n10954;
   wire n10955;
   wire n10956;
   wire n10957;
   wire n10958;
   wire n10959;
   wire n10960;
   wire n10961;
   wire n10962;
   wire n10963;
   wire n10964;
   wire n10965;
   wire n10966;
   wire n10967;
   wire n10968;
   wire n10969;
   wire n10970;
   wire n10971;
   wire n10972;
   wire n10973;
   wire n10974;
   wire n10975;
   wire n10976;
   wire n10977;
   wire n10978;
   wire n10979;
   wire n10980;
   wire n10981;
   wire n10982;
   wire n10983;
   wire n10984;
   wire n10985;
   wire n10986;
   wire n10987;
   wire n10988;
   wire n10989;
   wire n10990;
   wire n10991;
   wire n10992;
   wire n10993;
   wire n10994;
   wire n10995;
   wire n10996;
   wire n10997;
   wire n10998;
   wire n10999;
   wire n11000;
   wire n11001;
   wire n11002;
   wire n11003;
   wire n11004;
   wire n11005;
   wire n11006;
   wire n11007;
   wire n11008;
   wire n11009;
   wire n11010;
   wire n11011;
   wire n11012;
   wire n11013;
   wire n11014;
   wire n11015;
   wire n11016;
   wire n11017;
   wire n11018;
   wire n11019;
   wire n11020;
   wire n11021;
   wire n11022;
   wire n11023;
   wire n11024;
   wire n11025;
   wire n11026;
   wire n11027;
   wire n11028;
   wire n11029;
   wire n11030;
   wire n11031;
   wire n11032;
   wire n11033;
   wire n11034;
   wire n11035;
   wire n11036;
   wire n11037;
   wire n11038;
   wire n11039;
   wire n11040;
   wire n11041;
   wire n11042;
   wire n11043;
   wire n11044;
   wire n11045;
   wire n11046;
   wire n11047;
   wire n11048;
   wire n11049;
   wire n11050;
   wire n11051;
   wire n11052;
   wire n11053;
   wire n11054;
   wire n11055;
   wire n11056;
   wire n11057;
   wire n11058;
   wire n11059;
   wire n11060;
   wire n11061;
   wire n11062;
   wire n11063;
   wire n11064;
   wire n11065;
   wire n11066;
   wire n11067;
   wire n11068;
   wire n11069;
   wire n11070;
   wire n11071;
   wire n11072;
   wire n11073;
   wire n11074;
   wire n11075;
   wire n11076;
   wire n11077;
   wire n11078;
   wire n11079;
   wire n11080;
   wire n11081;
   wire n11082;
   wire n11083;
   wire n11084;
   wire n11085;
   wire n11086;
   wire n11087;
   wire n11088;
   wire n11089;
   wire n11090;
   wire n11091;
   wire n11092;
   wire n11093;
   wire n11094;
   wire n11095;
   wire n11096;
   wire n11097;
   wire n11098;
   wire n11099;
   wire n11100;
   wire n11101;
   wire n11102;
   wire n11103;
   wire n11104;
   wire n11105;
   wire n11106;
   wire n11107;
   wire n11108;
   wire n11109;
   wire n11110;
   wire n11111;
   wire n11112;
   wire n11113;
   wire n11114;
   wire n11115;
   wire n11116;
   wire n11117;
   wire n11118;
   wire n11119;
   wire n11120;
   wire n11121;
   wire n11122;
   wire n11123;
   wire n11124;
   wire n11125;
   wire n11126;
   wire n11127;
   wire n11128;
   wire n11129;
   wire n11130;
   wire n11131;
   wire n11132;
   wire n11133;
   wire n11134;
   wire n11135;
   wire n11136;
   wire n11137;
   wire n11138;
   wire n11139;
   wire n11140;
   wire n11141;
   wire n11142;
   wire n11143;
   wire n11144;
   wire n11145;
   wire n11146;
   wire n11147;
   wire n11148;
   wire n11149;
   wire n11150;
   wire n11151;
   wire n11152;
   wire n11153;
   wire n11154;
   wire n11155;
   wire n11156;
   wire n11157;
   wire n11158;
   wire n11159;
   wire n11160;
   wire n11161;
   wire n11162;
   wire n11163;
   wire n11164;
   wire n11165;
   wire n11166;
   wire n11167;
   wire n11168;
   wire n11169;
   wire n11170;
   wire n11171;
   wire n11172;
   wire n11173;
   wire n11174;
   wire n11175;
   wire n11176;
   wire n11177;
   wire n11178;
   wire n11179;
   wire n11180;
   wire n11181;
   wire n11182;
   wire n11183;
   wire n11184;
   wire n11185;
   wire n11186;
   wire n11187;
   wire n11188;
   wire n11189;
   wire n11190;
   wire n11191;
   wire n11192;
   wire n11193;
   wire n11194;
   wire n11195;
   wire n11196;
   wire n11197;
   wire n11198;
   wire n11199;
   wire n11200;
   wire n11201;
   wire n11202;
   wire n11203;
   wire n11204;
   wire n11205;
   wire n11206;
   wire n11207;
   wire n11208;
   wire n11209;
   wire n11210;
   wire n11211;
   wire n11212;
   wire n11213;
   wire n11214;
   wire n11215;
   wire n11216;
   wire n11217;
   wire n11218;
   wire n11219;
   wire n11220;
   wire n11221;
   wire n11222;
   wire n11223;
   wire n11224;
   wire n11225;
   wire n11226;
   wire n11227;
   wire n11228;
   wire n11229;
   wire n11230;
   wire n11231;
   wire n11232;
   wire n11233;
   wire n11234;
   wire n11235;
   wire n11236;
   wire n11237;
   wire n11238;
   wire n11239;
   wire n11240;
   wire n11241;
   wire n11242;
   wire n11243;
   wire n11244;
   wire n11245;
   wire n11246;
   wire n11247;
   wire n11248;
   wire n11249;
   wire n11250;
   wire n11251;
   wire n11252;
   wire n11253;
   wire n11254;
   wire n11255;
   wire n11256;
   wire n11257;
   wire n11258;
   wire n11259;
   wire n11260;
   wire n11261;
   wire n11262;
   wire n11263;
   wire n11264;
   wire n11265;
   wire n11266;
   wire n11267;
   wire n11268;
   wire n11269;
   wire n11270;
   wire n11271;
   wire n11272;
   wire n11273;
   wire n11274;
   wire n11275;
   wire n11276;
   wire n11277;
   wire n11278;
   wire n11279;
   wire n11280;
   wire n11281;
   wire n11282;
   wire n11283;
   wire n11284;
   wire n11285;
   wire n11286;
   wire n11287;
   wire n11288;
   wire n11289;
   wire n11290;
   wire n11291;
   wire n11292;
   wire n11293;
   wire n11294;
   wire n11295;
   wire n11296;
   wire n11297;
   wire n11298;
   wire n11299;
   wire n11300;
   wire n11301;
   wire n11302;
   wire n11303;
   wire n11304;
   wire n11305;
   wire n11306;
   wire n11307;
   wire n11308;
   wire n11309;
   wire n11310;
   wire n11311;
   wire n11312;
   wire n11313;
   wire n11314;
   wire n11315;
   wire n11316;
   wire n11317;
   wire n11318;
   wire n11319;
   wire n11320;
   wire n11321;
   wire n11322;
   wire n11323;
   wire n11324;
   wire n11325;
   wire n11326;
   wire n11327;
   wire n11328;
   wire n11329;
   wire n11330;
   wire n11331;
   wire n11332;
   wire n11333;
   wire n11334;
   wire n11335;
   wire n11336;
   wire n11337;
   wire n11338;
   wire n11339;
   wire n11340;
   wire n11341;
   wire n11342;
   wire n11343;
   wire n11344;
   wire n11345;
   wire n11346;
   wire n11347;
   wire n11348;
   wire n11349;
   wire n11350;
   wire n11351;
   wire n11352;
   wire n11353;
   wire n11354;
   wire n11355;
   wire n11356;
   wire n11357;
   wire n11358;
   wire n11359;
   wire n11360;
   wire n11361;
   wire n11362;
   wire n11363;
   wire n11364;
   wire n11365;
   wire n11366;
   wire n11367;
   wire n11368;
   wire n11369;
   wire n11370;
   wire n11371;
   wire n11372;
   wire n11373;
   wire n11374;
   wire n11375;
   wire n11376;
   wire n11377;
   wire n11378;
   wire n11379;
   wire n11380;
   wire n11381;
   wire n11382;
   wire n11383;
   wire n11384;
   wire n11385;
   wire n11386;
   wire n11387;
   wire n11388;
   wire n11389;
   wire n11390;
   wire n11391;
   wire n11392;
   wire n11393;
   wire n11394;
   wire n11395;
   wire n11396;
   wire n11397;
   wire n11398;
   wire n11399;
   wire n11400;
   wire n11401;
   wire n11402;
   wire n11403;
   wire n11404;
   wire n11405;
   wire n11406;
   wire n11407;
   wire n11408;
   wire n11409;
   wire n11410;
   wire n11411;
   wire n11412;
   wire n11413;
   wire n11414;
   wire n11415;
   wire n11416;
   wire n11417;
   wire n11418;
   wire n11419;
   wire n11420;
   wire n11421;
   wire n11422;
   wire n11423;
   wire n11424;
   wire n11425;
   wire n11426;
   wire n11427;
   wire n11428;
   wire n11429;
   wire n11430;
   wire n11431;
   wire n11432;
   wire n11433;
   wire n11434;
   wire n11435;
   wire n11436;
   wire n11437;
   wire n11438;
   wire n11439;
   wire n11440;
   wire n11441;
   wire n11442;
   wire n11443;
   wire n11444;
   wire n11445;
   wire n11446;
   wire n11447;
   wire n11448;
   wire n11449;
   wire n11450;
   wire n11451;
   wire n11452;
   wire n11453;
   wire n11454;
   wire n11455;
   wire n11456;
   wire n11457;
   wire n11458;
   wire n11459;
   wire n11460;
   wire n11461;
   wire n11462;
   wire n11463;
   wire n11464;
   wire n11465;
   wire n11466;
   wire n11467;
   wire n11468;
   wire n11469;
   wire n11470;
   wire n11471;
   wire n11472;
   wire n11473;
   wire n11474;
   wire n11475;
   wire n11476;
   wire n11477;
   wire n11478;
   wire n11479;
   wire n11480;
   wire n11481;
   wire n11482;
   wire n11483;
   wire n11484;
   wire n11485;
   wire n11486;
   wire n11487;
   wire n11488;
   wire n11489;
   wire n11490;
   wire n11491;
   wire n11492;
   wire n11493;
   wire n11494;
   wire n11495;
   wire n11496;
   wire n11497;
   wire n11498;
   wire n11499;
   wire n11500;
   wire n11501;
   wire n11502;
   wire n11503;
   wire n11504;
   wire n11505;
   wire n11506;
   wire n11507;
   wire n11508;
   wire n11509;
   wire n11510;
   wire n11511;
   wire n11512;
   wire n11513;
   wire n11514;
   wire n11515;
   wire n11516;
   wire n11517;
   wire n11518;
   wire n11519;
   wire n11520;
   wire n11521;
   wire n11522;
   wire n11523;
   wire n11524;
   wire n11525;
   wire n11526;
   wire n11527;
   wire n11528;
   wire n11529;
   wire n11530;
   wire n11531;
   wire n11532;
   wire n11533;
   wire n11534;
   wire n11535;
   wire n11536;
   wire n11537;
   wire n11538;
   wire n11539;
   wire n11540;
   wire n11541;
   wire n11542;
   wire n11543;
   wire n11544;
   wire n11545;
   wire n11546;
   wire n11547;
   wire n11548;
   wire n11549;
   wire n11550;
   wire n11551;
   wire n11552;
   wire n11553;
   wire n11554;
   wire n11555;
   wire n11556;
   wire n11557;
   wire n11558;
   wire n11559;
   wire n11560;
   wire n11561;
   wire n11562;
   wire n11563;
   wire n11564;
   wire n11565;
   wire n11566;
   wire n11567;
   wire n11568;
   wire n11569;
   wire n11570;
   wire n11571;
   wire n11572;
   wire n11573;
   wire n11574;
   wire n11575;
   wire n11576;
   wire n11577;
   wire n11578;
   wire n11579;
   wire n11580;
   wire n11581;
   wire n11582;
   wire n11583;
   wire n11584;
   wire n11585;
   wire n11586;
   wire n11587;
   wire n11588;
   wire n11589;
   wire n11590;
   wire n11591;
   wire n11592;
   wire n11593;
   wire n11594;
   wire n11595;
   wire n11596;
   wire n11597;
   wire n11598;
   wire n11599;
   wire n11600;
   wire n11601;
   wire n11602;
   wire n11603;
   wire n11604;
   wire n11605;
   wire n11606;
   wire n11607;
   wire n11608;
   wire n11609;
   wire n11610;
   wire n11611;
   wire n11612;
   wire n11613;
   wire n11614;
   wire n11615;
   wire n11616;
   wire n11617;
   wire n11618;
   wire n11619;
   wire n11620;
   wire n11621;
   wire n11622;
   wire n11623;
   wire n11624;
   wire n11625;
   wire n11626;
   wire n11627;
   wire n11628;
   wire n11629;
   wire n11630;
   wire n11631;
   wire n11632;
   wire n11633;
   wire n11634;
   wire n11635;
   wire n11636;
   wire n11637;
   wire n11638;
   wire n11639;
   wire n11640;
   wire n11641;
   wire n11642;
   wire n11643;
   wire n11644;
   wire n11645;
   wire n11646;
   wire n11647;
   wire n11648;
   wire n11649;
   wire n11650;
   wire n11651;
   wire n11652;
   wire n11653;
   wire n11654;
   wire n11655;
   wire n11656;
   wire n11657;
   wire n11658;
   wire n11659;
   wire n11660;
   wire n11661;
   wire n11662;
   wire n11663;
   wire n11664;
   wire n11665;
   wire n11666;
   wire n11667;
   wire n11668;
   wire n11669;
   wire n11670;
   wire n11671;
   wire n11672;
   wire n11673;
   wire n11674;
   wire n11675;
   wire n11676;
   wire n11677;
   wire n11678;
   wire n11679;
   wire n11680;
   wire n11681;
   wire n11682;
   wire n11683;
   wire n11684;
   wire n11685;
   wire n11686;
   wire n11687;
   wire n11688;
   wire n11689;
   wire n11690;
   wire n11691;
   wire n11692;
   wire n11693;
   wire n11694;
   wire n11695;
   wire n11696;
   wire n11697;
   wire n11698;
   wire n11699;
   wire n11700;
   wire n11701;
   wire n11702;
   wire n11703;
   wire n11704;
   wire n11705;
   wire n11706;
   wire n11707;
   wire n11708;
   wire n11709;
   wire n11710;
   wire n11711;
   wire n11712;
   wire n11713;
   wire n11714;
   wire n11715;
   wire n11716;
   wire n11717;
   wire n11718;
   wire n11719;
   wire n11720;
   wire n11721;
   wire n11722;
   wire n11723;
   wire n11724;
   wire n11725;
   wire n11726;
   wire n11727;
   wire n11728;
   wire n11729;
   wire n11730;
   wire n11731;
   wire n11732;
   wire n11733;
   wire n11734;
   wire n11735;
   wire n11736;
   wire n11737;
   wire n11738;
   wire n11739;
   wire n11740;
   wire n11741;
   wire n11742;
   wire n11743;
   wire n11744;
   wire n11745;
   wire n11746;
   wire n11747;
   wire n11748;
   wire n11749;
   wire n11750;
   wire n11751;
   wire n11752;
   wire n11753;
   wire n11754;
   wire n11755;
   wire n11756;
   wire n11757;
   wire n11758;
   wire n11759;
   wire n11760;
   wire n11761;
   wire n11762;
   wire n11763;
   wire n11764;
   wire n11765;
   wire n11766;
   wire n11767;
   wire n11768;
   wire n11769;
   wire n11770;
   wire n11771;
   wire n11772;
   wire n11773;
   wire n11774;
   wire n11775;
   wire n11776;
   wire n11777;
   wire n11778;
   wire n11779;
   wire n11780;
   wire n11781;
   wire n11782;
   wire n11783;
   wire n11784;
   wire n11785;
   wire n11786;
   wire n11787;
   wire n11788;
   wire n11789;
   wire n11790;
   wire n11791;
   wire n11792;
   wire n11793;
   wire n11794;
   wire n11795;
   wire n11796;
   wire n11797;
   wire n11798;
   wire n11799;
   wire n11800;
   wire n11801;
   wire n11802;
   wire n11803;
   wire n11804;
   wire n11805;
   wire n11806;
   wire n11807;
   wire n11808;
   wire n11809;
   wire n11810;
   wire n11811;
   wire n11812;
   wire n11813;
   wire n11814;
   wire n11815;
   wire n11816;
   wire n11817;
   wire n11818;
   wire n11819;
   wire n11820;
   wire n11821;
   wire n11822;
   wire n11823;
   wire n11824;
   wire n11825;
   wire n11826;
   wire n11827;
   wire n11828;
   wire n11829;
   wire n11830;
   wire n11831;
   wire n11832;
   wire n11833;
   wire n11834;
   wire n11835;
   wire n11836;
   wire n11837;
   wire n11838;
   wire n11839;
   wire n11840;
   wire n11841;
   wire n11842;
   wire n11843;
   wire n11844;
   wire n11845;
   wire n11846;
   wire n11847;
   wire n11848;
   wire n11849;
   wire n11850;
   wire n11851;
   wire n11852;
   wire n11853;
   wire n11854;
   wire n11855;
   wire n11856;
   wire n11857;
   wire n11858;
   wire n11859;
   wire n11860;
   wire n11861;
   wire n11862;
   wire n11863;
   wire n11864;
   wire n11865;
   wire n11866;
   wire n11867;
   wire n11868;
   wire n11869;
   wire n11870;
   wire n11871;
   wire n11872;
   wire n11873;
   wire n11874;
   wire n11875;
   wire n11876;
   wire n11877;
   wire n11878;
   wire n11879;
   wire n11880;
   wire n11881;
   wire n11882;
   wire n11883;
   wire n11884;
   wire n11885;
   wire n11886;
   wire n11887;
   wire n11888;
   wire n11889;
   wire n11890;
   wire n11891;
   wire n11892;
   wire n11893;
   wire n11894;
   wire n11895;
   wire n11896;
   wire n11897;
   wire n11898;
   wire n11899;
   wire n11900;
   wire n11901;
   wire n11902;
   wire n11903;
   wire n11904;
   wire n11905;
   wire n11906;
   wire n11907;
   wire n11908;
   wire n11909;
   wire n11910;
   wire n11911;
   wire n11912;
   wire n11913;
   wire n11914;
   wire n11915;
   wire n11916;
   wire n11917;
   wire n11918;
   wire n11919;
   wire n11920;
   wire n11921;
   wire n11922;
   wire n11923;
   wire n11924;
   wire n11925;
   wire n11926;
   wire n11927;
   wire n11928;
   wire n11929;
   wire n11930;
   wire n11931;
   wire n11932;
   wire n11933;
   wire n11934;
   wire n11935;
   wire n11936;
   wire n11937;
   wire n11938;
   wire n11939;
   wire n11940;
   wire n11941;
   wire n11942;
   wire n11943;
   wire n11944;
   wire n11945;
   wire n11946;
   wire n11947;
   wire n11948;
   wire n11949;
   wire n11950;
   wire n11951;
   wire n11952;
   wire n11953;
   wire n11954;
   wire n11955;
   wire n11956;
   wire n11957;
   wire n11958;
   wire n11959;
   wire n11960;
   wire n11961;
   wire n11962;
   wire n11963;
   wire n11964;
   wire n11965;
   wire n11966;
   wire n11967;
   wire n11968;
   wire n11969;
   wire n11970;
   wire n11971;
   wire n11972;
   wire n11973;
   wire n11974;
   wire n11975;
   wire n11976;
   wire n11977;
   wire n11978;
   wire n11979;
   wire n11980;
   wire n11981;
   wire n11982;
   wire n11983;
   wire n11984;
   wire n11985;
   wire n11986;
   wire n11987;
   wire n11988;
   wire n11989;
   wire n11990;
   wire n11991;
   wire n11992;
   wire n11993;
   wire n11994;
   wire n11995;
   wire n11996;
   wire n11997;
   wire n11998;
   wire n11999;
   wire n12000;
   wire n12001;
   wire n12002;
   wire n12003;
   wire n12004;
   wire n12005;
   wire n12006;
   wire n12007;
   wire n12008;
   wire n12009;
   wire n12010;
   wire n12011;
   wire n12012;
   wire n12013;
   wire n12014;
   wire n12015;
   wire n12016;
   wire n12017;
   wire n12018;
   wire n12019;
   wire n12020;
   wire n12021;
   wire n12022;
   wire n12023;
   wire n12024;
   wire n12025;
   wire n12026;
   wire n12027;
   wire n12028;
   wire n12029;
   wire n12030;
   wire n12031;
   wire n12032;
   wire n12033;
   wire n12034;
   wire n12035;
   wire n12036;
   wire n12037;
   wire n12038;
   wire n12039;
   wire n12040;
   wire n12041;
   wire n12042;
   wire n12043;
   wire n12044;
   wire n12045;
   wire n12046;
   wire n12047;
   wire n12048;
   wire n12049;
   wire n12050;
   wire n12051;
   wire n12052;
   wire n12053;
   wire n12054;
   wire n12055;
   wire n12056;
   wire n12057;
   wire n12058;
   wire n12059;
   wire n12060;
   wire n12061;
   wire n12062;
   wire n12063;
   wire n12064;
   wire n12065;
   wire n12066;
   wire n12067;
   wire n12068;
   wire n12069;
   wire n12070;
   wire n12071;
   wire n12072;
   wire n12073;
   wire n12074;
   wire n12075;
   wire n12076;
   wire n12077;
   wire n12078;
   wire n12079;
   wire n12080;
   wire n12081;
   wire n12082;
   wire n12083;
   wire n12084;
   wire n12085;
   wire n12086;
   wire n12087;
   wire n12088;
   wire n12089;
   wire n12090;
   wire n12091;
   wire n12092;
   wire n12093;
   wire n12094;
   wire n12095;
   wire n12096;
   wire n12097;
   wire n12098;
   wire n12099;
   wire n12100;
   wire n12101;
   wire n12102;
   wire n12103;
   wire n12104;
   wire n12105;
   wire n12106;
   wire n12107;
   wire n12108;
   wire n12109;
   wire n12110;
   wire n12111;
   wire n12112;
   wire n12113;
   wire n12114;
   wire n12115;
   wire n12116;
   wire n12117;
   wire n12118;
   wire n12119;
   wire n12120;
   wire n12121;
   wire n12122;
   wire n12123;
   wire n12124;
   wire n12125;
   wire n12126;
   wire n12127;
   wire n12128;
   wire n12129;
   wire n12130;
   wire n12131;
   wire n12132;
   wire n12133;
   wire n12134;
   wire n12135;
   wire n12136;
   wire n12137;
   wire n12138;
   wire n12139;
   wire n12140;
   wire n12141;
   wire n12142;
   wire n12143;
   wire n12144;
   wire n12145;
   wire n12146;
   wire n12147;
   wire n12148;
   wire n12149;
   wire n12150;
   wire n12151;
   wire n12152;
   wire n12153;
   wire n12154;
   wire n12155;
   wire n12156;
   wire n12157;
   wire n12158;
   wire n12159;
   wire n12160;
   wire n12161;
   wire n12162;
   wire n12163;
   wire n12164;
   wire n12165;
   wire n12166;
   wire n12167;
   wire n12168;
   wire n12169;
   wire n12170;
   wire n12171;
   wire n12172;
   wire n12173;
   wire n12174;
   wire n12175;
   wire n12176;
   wire n12177;
   wire n12178;
   wire n12179;
   wire n12180;
   wire n12181;
   wire n12182;
   wire n12183;
   wire n12184;
   wire n12185;
   wire n12186;
   wire n12187;
   wire n12188;
   wire n12189;
   wire n12190;
   wire n12191;
   wire n12192;
   wire n12193;
   wire n12194;
   wire n12195;
   wire n12196;
   wire n12197;
   wire n12198;
   wire n12199;
   wire n12200;
   wire n12201;
   wire n12202;
   wire n12203;
   wire n12204;
   wire n12205;
   wire n12206;
   wire n12207;
   wire n12208;
   wire n12209;
   wire n12210;
   wire n12211;
   wire n12212;
   wire n12213;
   wire n12214;
   wire n12215;
   wire n12216;
   wire n12217;
   wire n12218;
   wire n12219;
   wire n12220;
   wire n12221;
   wire n12222;
   wire n12223;
   wire n12224;
   wire n12225;
   wire n12226;
   wire n12227;
   wire n12228;
   wire n12229;
   wire n12230;
   wire n12231;
   wire n12232;
   wire n12233;
   wire n12234;
   wire n12235;
   wire n12236;
   wire n12237;
   wire n12238;
   wire n12239;
   wire n12240;
   wire n12241;
   wire n12242;
   wire n12243;
   wire n12244;
   wire n12245;
   wire n12246;
   wire n12247;
   wire n12248;
   wire n12249;
   wire n12250;
   wire n12251;
   wire n12252;
   wire n12253;
   wire n12254;
   wire n12255;
   wire n12256;
   wire n12257;
   wire n12258;
   wire n12259;
   wire n12260;
   wire n12261;
   wire n12262;
   wire n12263;
   wire n12264;
   wire n12265;
   wire n12266;
   wire n12267;
   wire n12268;
   wire n12269;
   wire n12270;
   wire n12271;
   wire n12272;
   wire n12273;
   wire n12274;
   wire n12275;
   wire n12276;
   wire n12277;
   wire n12278;
   wire n12279;
   wire n12280;
   wire n12281;
   wire n12282;
   wire n12283;
   wire n12284;
   wire n12285;
   wire n12286;
   wire n12287;
   wire n12288;
   wire n12289;
   wire n12290;
   wire n12291;
   wire n12292;
   wire n12293;
   wire n12294;
   wire n12295;
   wire n12296;
   wire n12297;
   wire n12298;
   wire n12299;
   wire n12300;
   wire n12301;
   wire n12302;
   wire n12303;
   wire n12304;
   wire n12305;
   wire n12306;
   wire n12307;
   wire n12308;
   wire n12309;
   wire n12310;
   wire n12311;
   wire n12312;
   wire n12313;
   wire n12314;
   wire n12315;
   wire n12316;
   wire n12317;
   wire n12318;
   wire n12319;
   wire n12320;
   wire n12321;
   wire n12322;
   wire n12323;
   wire n12324;
   wire n12325;
   wire n12326;
   wire n12327;
   wire n12328;
   wire n12329;
   wire n12330;
   wire n12331;
   wire n12332;
   wire n12333;
   wire n12334;
   wire n12335;
   wire n12336;
   wire n12337;
   wire n12338;
   wire n12339;
   wire n12340;
   wire n12341;
   wire n12342;
   wire n12343;
   wire n12344;
   wire n12345;
   wire n12346;
   wire n12347;
   wire n12348;
   wire n12349;
   wire n12350;
   wire n12351;
   wire n12352;
   wire n12353;
   wire n12354;
   wire n12355;
   wire n12356;
   wire n12357;
   wire n12358;
   wire n12359;
   wire n12360;
   wire n12361;
   wire n12362;
   wire n12363;
   wire n12364;
   wire n12365;
   wire n12366;
   wire n12367;
   wire n12368;
   wire n12369;
   wire n12370;
   wire n12371;
   wire n12372;
   wire n12373;
   wire n12374;
   wire n12375;
   wire n12376;
   wire n12377;
   wire n12378;
   wire n12379;
   wire n12380;
   wire n12381;
   wire n12382;
   wire n12383;
   wire n12384;
   wire n12385;
   wire n12386;
   wire n12387;
   wire n12388;
   wire n12389;
   wire n12390;
   wire n12391;
   wire n12392;
   wire n12393;
   wire n12394;
   wire n12395;
   wire n12396;
   wire n12397;
   wire n12398;
   wire n12399;
   wire n12400;
   wire n12401;
   wire n12402;
   wire n12403;
   wire n12404;
   wire n12405;
   wire n12406;
   wire n12407;
   wire n12408;
   wire n12409;
   wire n12410;
   wire n12411;
   wire n12412;
   wire n12413;
   wire n12414;
   wire n12415;
   wire n12416;
   wire n12417;
   wire n12418;
   wire n12419;
   wire n12420;
   wire n12421;
   wire n12422;
   wire n12423;
   wire n12424;
   wire n12425;
   wire n12426;
   wire n12427;
   wire n12428;
   wire n12429;
   wire n12430;
   wire n12431;
   wire n12432;
   wire n12433;
   wire n12434;
   wire n12435;
   wire n12436;
   wire n12437;
   wire n12438;
   wire n12439;
   wire n12440;
   wire n12441;
   wire n12442;
   wire n12443;
   wire n12444;
   wire n12445;
   wire n12446;
   wire n12447;
   wire n12448;
   wire n12449;
   wire n12450;
   wire n12451;
   wire n12452;
   wire n12453;
   wire n12454;
   wire n12455;
   wire n12456;
   wire n12457;
   wire n12458;
   wire n12459;
   wire n12460;
   wire n12461;
   wire n12462;
   wire n12463;
   wire n12464;
   wire n12465;
   wire n12466;
   wire n12467;
   wire n12468;
   wire n12469;
   wire n12470;
   wire n12471;
   wire n12472;
   wire n12473;
   wire n12474;
   wire n12475;
   wire n12476;
   wire n12477;
   wire n12478;
   wire n12479;
   wire n12480;
   wire n12481;
   wire n12482;
   wire n12483;
   wire n12484;
   wire n12485;
   wire n12486;
   wire n12487;
   wire n12488;
   wire n12489;
   wire n12490;
   wire n12491;
   wire n12492;
   wire n12493;
   wire n12494;
   wire n12495;
   wire n12496;
   wire n12497;
   wire n12498;
   wire n12499;
   wire n12500;
   wire n12501;
   wire n12502;
   wire n12503;
   wire n12504;
   wire n12505;
   wire n12506;
   wire n12507;
   wire n12508;
   wire n12509;
   wire n12510;
   wire n12511;
   wire n12512;
   wire n12513;
   wire n12514;
   wire n12515;
   wire n12516;
   wire n12517;
   wire n12518;
   wire n12519;
   wire n12520;
   wire n12521;
   wire n12522;
   wire n12523;
   wire n12524;
   wire n12525;
   wire n12526;
   wire n12527;
   wire n12528;
   wire n12529;
   wire n12530;
   wire n12531;
   wire n12532;
   wire n12533;
   wire n12534;
   wire n12535;
   wire n12536;
   wire n12537;
   wire n12538;
   wire n12539;
   wire n12540;
   wire n12541;
   wire n12542;
   wire n12543;
   wire n12544;
   wire n12545;
   wire n12546;
   wire n12547;
   wire n12548;
   wire n12549;
   wire n12550;
   wire n12551;
   wire n12552;
   wire n12553;
   wire n12554;
   wire n12555;
   wire n12556;
   wire n12557;
   wire n12558;
   wire n12559;
   wire n12560;
   wire n12561;
   wire n12562;
   wire n12563;
   wire n12564;
   wire n12565;
   wire n12566;
   wire n12567;
   wire n12568;
   wire n12569;
   wire n12570;
   wire n12571;
   wire n12572;
   wire n12573;
   wire n12574;
   wire n12575;
   wire n12576;
   wire n12577;
   wire n12578;
   wire n12579;
   wire n12580;
   wire n12581;
   wire n12582;
   wire n12583;
   wire n12584;
   wire n12585;
   wire n12586;
   wire n12587;
   wire n12588;
   wire n12589;
   wire n12590;
   wire n12591;
   wire n12592;
   wire n12593;
   wire n12594;
   wire n12595;
   wire n12596;
   wire n12597;
   wire n12598;
   wire n12599;
   wire n12600;
   wire n12601;
   wire n12602;
   wire n12603;
   wire n12604;
   wire n12605;
   wire n12606;
   wire n12607;
   wire n12608;
   wire n12609;
   wire n12610;
   wire n12611;
   wire n12612;
   wire n12613;
   wire n12614;
   wire n12615;
   wire n12616;
   wire n12617;
   wire n12618;
   wire n12619;
   wire n12620;
   wire n12621;
   wire n12622;
   wire n12623;
   wire n12624;
   wire n12625;
   wire n12626;
   wire n12627;
   wire n12628;
   wire n12629;
   wire n12630;
   wire n12631;
   wire n12632;
   wire n12633;
   wire n12634;
   wire n12635;
   wire n12636;
   wire n12637;
   wire n12638;
   wire n12639;
   wire n12640;
   wire n12641;
   wire n12642;
   wire n12643;
   wire n12644;
   wire n12645;
   wire n12646;
   wire n12647;
   wire n12648;
   wire n12649;
   wire n12650;
   wire n12651;
   wire n12652;
   wire n12653;
   wire n12654;
   wire n12655;
   wire n12656;
   wire n12657;
   wire n12658;
   wire n12659;
   wire n12660;
   wire n12661;
   wire n12662;
   wire n12663;
   wire n12664;
   wire n12665;
   wire n12666;
   wire n12667;
   wire n12668;
   wire n12669;
   wire n12670;
   wire n12671;
   wire n12672;
   wire n12673;
   wire n12674;
   wire n12675;
   wire n12676;
   wire n12677;
   wire n12678;
   wire n12679;
   wire n12680;
   wire n12681;
   wire n12682;
   wire n12683;
   wire n12684;
   wire n12685;
   wire n12686;
   wire n12687;
   wire n12688;
   wire n12689;
   wire n12690;
   wire n12691;
   wire n12692;
   wire n12693;
   wire n12694;
   wire n12695;
   wire n12696;
   wire n12697;
   wire n12698;
   wire n12699;
   wire n12700;
   wire n12701;
   wire n12702;
   wire n12703;
   wire n12704;
   wire n12705;
   wire n12706;
   wire n12707;
   wire n12708;
   wire n12709;
   wire n12710;
   wire n12711;
   wire n12712;
   wire n12713;
   wire n12714;
   wire n12715;
   wire n12716;
   wire n12717;
   wire n12718;
   wire n12719;
   wire n12720;
   wire n12721;
   wire n12722;
   wire n12723;
   wire n12724;
   wire n12725;
   wire n12726;
   wire n12727;
   wire n12728;
   wire n12729;
   wire n12730;
   wire n12731;
   wire n12732;
   wire n12733;
   wire n12734;
   wire n12735;
   wire n12736;
   wire n12737;
   wire n12738;
   wire n12739;
   wire n12740;
   wire n12741;
   wire n12742;
   wire n12743;
   wire n12744;
   wire n12745;
   wire n12746;
   wire n12747;
   wire n12748;
   wire n12749;
   wire n12750;
   wire n12751;
   wire n12752;
   wire n12753;
   wire n12754;
   wire n12755;
   wire n12756;
   wire n12757;
   wire n12758;
   wire n12759;
   wire n12760;
   wire n12761;
   wire n12762;
   wire n12763;
   wire n12764;
   wire n12765;
   wire n12766;
   wire n12767;
   wire n12768;
   wire n12769;
   wire n12770;
   wire n12771;
   wire n12772;
   wire n12773;
   wire n12774;
   wire n12775;
   wire n12776;
   wire n12777;
   wire n12778;
   wire n12779;
   wire n12780;
   wire n12781;
   wire n12782;
   wire n12783;
   wire n12784;
   wire n12785;
   wire n12786;
   wire n12787;
   wire n12788;
   wire n12789;
   wire n12790;
   wire n12791;
   wire n12792;
   wire n12793;
   wire n12794;
   wire n12795;
   wire n12796;
   wire n12797;
   wire n12798;
   wire n12799;
   wire n12800;
   wire n12801;
   wire n12802;
   wire n12803;
   wire n12804;
   wire n12805;
   wire n12806;
   wire n12807;
   wire n12808;
   wire n12809;
   wire n12810;
   wire n12811;
   wire n12812;
   wire n12813;
   wire n12814;
   wire n12815;
   wire n12816;
   wire n12817;
   wire n12818;
   wire n12819;
   wire n12820;
   wire n12821;
   wire n12822;
   wire n12823;
   wire n12824;
   wire n12825;
   wire n12826;
   wire n12827;
   wire n12828;
   wire n12829;
   wire n12830;
   wire n12831;
   wire n12832;
   wire n12833;
   wire n12834;
   wire n12835;
   wire n12836;
   wire n12837;
   wire n12838;
   wire n12839;
   wire n12840;
   wire n12841;
   wire n12842;
   wire n12843;
   wire n12844;
   wire n12845;
   wire n12846;
   wire n12847;
   wire n12848;
   wire n12849;
   wire n12850;
   wire n12851;
   wire n12852;
   wire n12853;
   wire n12854;
   wire n12855;
   wire n12856;
   wire n12857;
   wire n12858;
   wire n12859;
   wire n12860;
   wire n12861;
   wire n12862;
   wire n12863;
   wire n12864;
   wire n12865;
   wire n12866;
   wire n12867;
   wire n12868;
   wire n12869;
   wire n12870;
   wire n12871;
   wire n12872;
   wire n12873;
   wire n12874;
   wire n12875;
   wire n12876;
   wire n12877;
   wire n12878;
   wire n12879;
   wire n12880;
   wire n12881;
   wire n12882;
   wire n12883;
   wire n12884;
   wire n12885;
   wire n12886;
   wire n12887;
   wire n12888;
   wire n12889;
   wire n12890;
   wire n12891;
   wire n12892;
   wire n12893;
   wire n12894;
   wire n12895;
   wire n12896;
   wire n12897;
   wire n12898;
   wire n12899;
   wire n12900;
   wire n12901;
   wire n12902;
   wire n12903;
   wire n12904;
   wire n12905;
   wire n12906;
   wire n12907;
   wire n12908;
   wire n12909;
   wire n12910;
   wire n12911;
   wire n12912;
   wire n12913;
   wire n12914;
   wire n12915;
   wire n12916;
   wire n12917;
   wire n12918;
   wire n12919;
   wire n12920;
   wire n12921;
   wire n12922;
   wire n12923;
   wire n12924;
   wire n12925;
   wire n12926;
   wire n12927;
   wire n12928;
   wire n12929;
   wire n12930;
   wire n12931;
   wire n12932;
   wire n12933;
   wire n12934;
   wire n12935;
   wire n12936;
   wire n12937;
   wire n12938;
   wire n12939;
   wire n12940;
   wire n12941;
   wire n12942;
   wire n12943;
   wire n12944;
   wire n12945;
   wire n12946;
   wire n12947;
   wire n12948;
   wire n12949;
   wire n12950;
   wire n12951;
   wire n12952;
   wire n12953;
   wire n12954;
   wire n12955;
   wire n12956;
   wire n12957;
   wire n12958;
   wire n12959;
   wire n12960;
   wire n12961;
   wire n12962;
   wire n12963;
   wire n12964;
   wire n12965;
   wire n12966;
   wire n12967;
   wire n12968;
   wire n12969;
   wire n12970;
   wire n12971;
   wire n12972;
   wire n12973;
   wire n12974;
   wire n12975;
   wire n12976;
   wire n12977;
   wire n12978;
   wire n12979;
   wire n12980;
   wire n12981;
   wire n12982;
   wire n12983;
   wire n12984;
   wire n12985;
   wire n12986;
   wire n12987;
   wire n12988;
   wire n12989;
   wire n12990;
   wire n12991;
   wire n12992;
   wire n12993;
   wire n12994;
   wire n12995;
   wire n12996;
   wire n12997;
   wire n12998;
   wire n12999;
   wire n13000;
   wire n13001;
   wire n13002;
   wire n13003;
   wire n13004;
   wire n13005;
   wire n13006;
   wire n13007;
   wire n13008;
   wire n13009;
   wire n13010;
   wire n13011;
   wire n13012;
   wire n13013;
   wire n13014;
   wire n13015;
   wire n13016;
   wire n13017;
   wire n13018;
   wire n13019;
   wire n13020;
   wire n13021;
   wire n13022;
   wire n13023;
   wire n13024;
   wire n13025;
   wire n13026;
   wire n13027;
   wire n13028;
   wire n13029;
   wire n13030;
   wire n13031;
   wire n13032;
   wire n13033;
   wire n13034;
   wire n13035;
   wire n13036;
   wire n13037;
   wire n13038;
   wire n13039;
   wire n13040;
   wire n13041;
   wire n13042;
   wire n13043;
   wire n13044;
   wire n13045;
   wire n13046;
   wire n13047;
   wire n13048;
   wire n13049;
   wire n13050;
   wire n13051;
   wire n13052;
   wire n13053;
   wire n13054;
   wire n13055;
   wire n13056;
   wire n13057;
   wire n13058;
   wire n13059;
   wire n13060;
   wire n13061;
   wire n13062;
   wire n13063;
   wire n13064;
   wire n13065;
   wire n13066;
   wire n13067;
   wire n13068;
   wire n13069;
   wire n13070;
   wire n13071;
   wire n13072;
   wire n13073;
   wire n13074;
   wire n13075;
   wire n13076;
   wire n13077;
   wire n13078;
   wire n13079;
   wire n13080;
   wire n13081;
   wire n13082;
   wire n13083;
   wire n13084;
   wire n13085;
   wire n13086;
   wire n13087;
   wire n13088;
   wire n13089;
   wire n13090;
   wire n13091;
   wire n13092;
   wire n13093;
   wire n13094;
   wire n13095;
   wire n13096;
   wire n13097;
   wire n13098;
   wire n13099;
   wire n13100;
   wire n13101;
   wire n13102;
   wire n13103;
   wire n13104;
   wire n13105;
   wire n13106;
   wire n13107;
   wire n13108;
   wire n13109;
   wire n13110;
   wire n13111;
   wire n13112;
   wire n13113;
   wire n13114;
   wire n13115;
   wire n13116;
   wire n13117;
   wire n13118;
   wire n13119;
   wire n13120;
   wire n13121;
   wire n13122;
   wire n13123;
   wire n13124;
   wire n13125;
   wire n13126;
   wire n13127;
   wire n13128;
   wire n13129;
   wire n13130;
   wire n13131;
   wire n13132;
   wire n13133;
   wire n13134;
   wire n13135;
   wire n13136;
   wire n13137;
   wire n13138;
   wire n13139;
   wire n13140;
   wire n13141;
   wire n13142;
   wire n13143;
   wire n13144;
   wire n13145;
   wire n13146;
   wire n13147;
   wire n13148;
   wire n13149;
   wire n13150;
   wire n13151;
   wire n13152;
   wire n13153;
   wire n13154;
   wire n13155;
   wire n13156;
   wire n13157;
   wire n13158;
   wire n13159;
   wire n13160;
   wire n13161;
   wire n13162;
   wire n13163;
   wire n13164;
   wire n13165;
   wire n13166;
   wire n13167;
   wire n13168;
   wire n13169;
   wire n13170;
   wire n13171;
   wire n13172;
   wire n13173;
   wire n13174;
   wire n13175;
   wire n13176;
   wire n13177;
   wire n13178;
   wire n13179;
   wire n13180;
   wire n13181;
   wire n13182;
   wire n13183;
   wire n13184;
   wire n13185;
   wire n13186;
   wire n13187;
   wire n13188;
   wire n13189;
   wire n13190;
   wire n13191;
   wire n13192;
   wire n13193;
   wire n13194;
   wire n13195;
   wire n13196;
   wire n13197;
   wire n13198;
   wire n13199;
   wire n13200;
   wire n13201;
   wire n13202;
   wire n13203;
   wire n13204;
   wire n13205;
   wire n13206;
   wire n13207;
   wire n13208;
   wire n13209;
   wire n13210;
   wire n13211;
   wire n13212;
   wire n13213;
   wire n13214;
   wire n13215;
   wire n13216;
   wire n13217;
   wire n13218;
   wire n13219;
   wire n13220;
   wire n13221;
   wire n13222;
   wire n13223;
   wire n13224;
   wire n13225;
   wire n13226;
   wire n13227;
   wire n13228;
   wire n13229;
   wire n13230;
   wire n13231;
   wire n13232;
   wire n13233;
   wire n13234;
   wire n13235;
   wire n13236;
   wire n13237;
   wire n13238;
   wire n13239;
   wire n13240;
   wire n13241;
   wire n13242;
   wire n13243;
   wire n13244;
   wire n13245;
   wire n13246;
   wire n13247;
   wire n13248;
   wire n13249;
   wire n13250;
   wire n13251;
   wire n13252;
   wire n13253;
   wire n13254;
   wire n13255;
   wire n13256;
   wire n13257;
   wire n13258;
   wire n13259;
   wire n13260;
   wire n13261;
   wire n13262;
   wire n13263;
   wire n13264;
   wire n13265;
   wire n13266;
   wire n13267;
   wire n13268;
   wire n13269;
   wire n13270;
   wire n13271;
   wire n13272;
   wire n13273;
   wire n13274;
   wire n13275;
   wire n13276;
   wire n13277;
   wire n13278;
   wire n13279;
   wire n13280;
   wire n13281;
   wire n13282;
   wire n13283;
   wire n13284;
   wire n13285;
   wire n13286;
   wire n13287;
   wire n13288;
   wire n13289;
   wire n13290;
   wire n13291;
   wire n13292;
   wire n13293;
   wire n13294;
   wire n13295;
   wire n13296;
   wire n13297;
   wire n13298;
   wire n13299;
   wire n13300;
   wire n13301;
   wire n13302;
   wire n13303;
   wire n13304;
   wire n13305;
   wire n13306;
   wire n13307;
   wire n13308;
   wire n13309;
   wire n13310;
   wire n13311;
   wire n13312;
   wire n13313;
   wire n13314;
   wire n13315;
   wire n13316;
   wire n13317;
   wire n13318;
   wire n13319;
   wire n13320;
   wire n13321;
   wire n13322;
   wire n13323;
   wire n13324;
   wire n13325;
   wire n13326;
   wire n13327;
   wire n13328;
   wire n13329;
   wire n13330;
   wire n13331;
   wire n13332;
   wire n13333;
   wire n13334;
   wire n13335;
   wire n13336;
   wire n13337;
   wire n13338;
   wire n13339;
   wire n13340;
   wire n13341;
   wire n13342;
   wire n13343;
   wire n13344;
   wire n13345;
   wire n13346;
   wire n13347;
   wire n13348;
   wire n13349;
   wire n13350;
   wire n13351;
   wire n13352;
   wire n13353;
   wire n13354;
   wire n13355;
   wire n13356;
   wire n13357;
   wire n13358;
   wire n13359;
   wire n13360;
   wire n13361;
   wire n13362;
   wire n13363;
   wire n13364;
   wire n13365;
   wire n13366;
   wire n13367;
   wire n13368;
   wire n13369;
   wire n13370;
   wire n13371;
   wire n13372;
   wire n13373;
   wire n13374;
   wire n13375;
   wire n13376;
   wire n13377;
   wire n13378;
   wire n13379;
   wire n13380;
   wire n13381;
   wire n13382;
   wire n13383;
   wire n13384;
   wire n13385;
   wire n13386;
   wire n13387;
   wire n13388;
   wire n13389;
   wire n13390;
   wire n13391;
   wire n13392;
   wire n13393;
   wire n13394;
   wire n13395;
   wire n13396;
   wire n13397;
   wire n13398;
   wire n13399;
   wire n13400;
   wire n13401;
   wire n13402;
   wire n13403;
   wire n13404;
   wire n13405;
   wire n13406;
   wire n13407;
   wire n13408;
   wire n13409;
   wire n13410;
   wire n13411;
   wire n13412;
   wire n13413;
   wire n13414;
   wire n13415;
   wire n13416;
   wire n13417;
   wire n13418;
   wire n13419;
   wire n13420;
   wire n13421;
   wire n13422;
   wire n13423;
   wire n13424;
   wire n13425;
   wire n13426;
   wire n13427;
   wire n13428;
   wire n13429;
   wire n13430;
   wire n13431;
   wire n13432;
   wire n13433;
   wire n13434;
   wire n13435;
   wire n13436;
   wire n13437;
   wire n13438;
   wire n13439;
   wire n13440;
   wire n13441;
   wire n13442;
   wire n13443;
   wire n13444;
   wire n13445;
   wire n13446;
   wire n13447;
   wire n13448;
   wire n13449;
   wire n13450;
   wire n13451;
   wire n13452;
   wire n13453;
   wire n13454;
   wire n13455;
   wire n13456;
   wire n13457;
   wire n13458;
   wire n13459;
   wire n13460;
   wire n13461;
   wire n13462;
   wire n13463;
   wire n13464;
   wire n13465;
   wire n13466;
   wire n13467;
   wire n13468;
   wire n13469;
   wire n13470;
   wire n13471;
   wire n13472;
   wire n13473;
   wire n13474;
   wire n13475;
   wire n13476;
   wire n13477;
   wire n13478;
   wire n13479;
   wire n13480;
   wire n13481;
   wire n13482;
   wire n13483;
   wire n13484;
   wire n13485;
   wire n13486;
   wire n13487;
   wire n13488;
   wire n13489;
   wire n13490;
   wire n13491;
   wire n13492;
   wire n13493;
   wire n13494;
   wire n13495;
   wire n13496;
   wire n13497;
   wire n13498;
   wire n13499;
   wire n13500;
   wire n13501;
   wire n13502;
   wire n13503;
   wire n13504;
   wire n13505;
   wire n13506;
   wire n13507;
   wire n13508;
   wire n13509;
   wire n13510;
   wire n13511;
   wire n13512;
   wire n13513;
   wire n13514;
   wire n13515;
   wire n13516;
   wire n13517;
   wire n13518;
   wire n13519;
   wire n13520;
   wire n13521;
   wire n13522;
   wire n13523;
   wire n13524;
   wire n13525;
   wire n13526;
   wire n13527;
   wire n13528;
   wire n13529;
   wire n13530;
   wire n13531;
   wire n13532;
   wire n13533;
   wire n13534;
   wire n13535;
   wire n13536;
   wire n13537;
   wire n13538;
   wire n13539;
   wire n13540;
   wire n13541;
   wire n13542;
   wire n13543;
   wire n13544;
   wire n13545;
   wire n13546;
   wire n13547;
   wire n13548;
   wire n13549;
   wire n13550;
   wire n13551;
   wire n13552;
   wire n13553;
   wire n13554;
   wire n13555;
   wire n13556;
   wire n13557;
   wire n13558;
   wire n13559;
   wire n13560;
   wire n13561;
   wire n13562;
   wire n13563;
   wire n13564;
   wire n13565;
   wire n13566;
   wire n13567;
   wire n13568;
   wire n13569;
   wire n13570;
   wire n13571;
   wire n13572;
   wire n13573;
   wire n13574;
   wire n13575;
   wire n13576;
   wire n13577;
   wire n13578;
   wire n13579;
   wire n13580;
   wire n13581;
   wire n13582;
   wire n13583;
   wire n13584;
   wire n13585;
   wire n13586;
   wire n13587;
   wire n13588;
   wire n13589;
   wire n13590;
   wire n13591;
   wire n13592;
   wire n13593;
   wire n13594;
   wire n13595;
   wire n13596;
   wire n13597;
   wire n13598;
   wire n13599;
   wire n13600;
   wire n13601;
   wire n13602;
   wire n13603;
   wire n13604;
   wire n13605;
   wire n13606;
   wire n13607;
   wire n13608;
   wire n13609;
   wire n13610;
   wire n13611;
   wire n13612;
   wire n13613;
   wire n13614;
   wire n13615;
   wire n13616;
   wire n13617;
   wire n13618;
   wire n13619;
   wire n13620;
   wire n13621;
   wire n13622;
   wire n13623;
   wire n13624;
   wire n13625;
   wire n13626;
   wire n13627;
   wire n13628;
   wire n13629;
   wire n13630;
   wire n13631;
   wire n13632;
   wire n13633;
   wire n13634;
   wire n13635;
   wire n13636;
   wire n13637;
   wire n13638;
   wire n13639;
   wire n13640;
   wire n13641;
   wire n13642;
   wire n13643;
   wire n13644;
   wire n13645;
   wire n13646;
   wire n13647;
   wire n13648;
   wire n13649;
   wire n13650;
   wire n13651;
   wire n13652;
   wire n13653;
   wire n13654;
   wire n13655;
   wire n13656;
   wire n13657;
   wire n13658;
   wire n13659;
   wire n13660;
   wire n13661;
   wire n13662;
   wire n13663;
   wire n13664;
   wire n13665;
   wire n13666;
   wire n13667;
   wire n13668;
   wire n13669;
   wire n13670;
   wire n13671;
   wire n13672;
   wire n13673;
   wire n13674;
   wire n13675;
   wire n13676;
   wire n13677;
   wire n13678;
   wire n13679;
   wire n13680;
   wire n13681;
   wire n13682;
   wire n13683;
   wire n13684;
   wire n13685;
   wire n13686;
   wire n13687;
   wire n13688;
   wire n13689;
   wire n13690;
   wire n13691;
   wire n13692;
   wire n13693;
   wire n13694;
   wire n13695;
   wire n13696;
   wire n13697;
   wire n13698;
   wire n13699;
   wire n13700;
   wire n13701;
   wire n13702;
   wire n13703;
   wire n13704;
   wire n13705;
   wire n13706;
   wire n13707;
   wire n13708;
   wire n13709;
   wire n13710;
   wire n13711;
   wire n13712;
   wire n13713;
   wire n13714;
   wire n13715;
   wire n13716;
   wire n13717;
   wire n13718;
   wire n13719;
   wire n13720;
   wire n13721;
   wire n13722;
   wire n13723;
   wire n13724;
   wire n13725;
   wire n13726;
   wire n13727;
   wire n13728;
   wire n13729;
   wire n13730;
   wire n13731;
   wire n13732;
   wire n13733;
   wire n13734;
   wire n13735;
   wire n13736;
   wire n13737;
   wire n13738;
   wire n13739;
   wire n13740;
   wire n13741;
   wire n13742;
   wire n13743;
   wire n13744;
   wire n13745;
   wire n13746;
   wire n13747;
   wire n13748;
   wire n13749;
   wire n13750;
   wire n13751;
   wire n13752;
   wire n13753;
   wire n13754;
   wire n13755;
   wire n13756;
   wire n13757;
   wire n13758;
   wire n13759;
   wire n13760;
   wire n13761;
   wire n13762;
   wire n13763;
   wire n13764;
   wire n13765;
   wire n13766;
   wire n13767;
   wire n13768;
   wire n13769;
   wire n13770;
   wire n13771;
   wire n13772;
   wire n13773;
   wire n13774;
   wire n13775;
   wire n13776;
   wire n13777;
   wire n13778;
   wire n13779;
   wire n13780;
   wire n13781;
   wire n13782;
   wire n13783;
   wire n13784;
   wire n13785;
   wire n13786;
   wire n13787;
   wire n13788;
   wire n13789;
   wire n13790;
   wire n13791;
   wire n13792;
   wire n13793;
   wire n13794;
   wire n13795;
   wire n13796;
   wire n13797;
   wire n13798;
   wire n13799;
   wire n13800;
   wire n13801;
   wire n13802;
   wire n13803;
   wire n13804;
   wire n13805;
   wire n13806;
   wire n13807;
   wire n13808;
   wire n13809;
   wire n13810;
   wire n13811;
   wire n13812;
   wire n13813;
   wire n13814;
   wire n13815;
   wire n13816;
   wire n13817;
   wire n13818;
   wire n13819;
   wire n13820;
   wire n13821;
   wire n13822;
   wire n13823;
   wire n13824;
   wire n13825;
   wire n13826;
   wire n13827;
   wire n13828;
   wire n13829;
   wire n13830;
   wire n13831;
   wire n13832;
   wire n13833;
   wire n13834;
   wire n13835;
   wire n13836;
   wire n13837;
   wire n13838;
   wire n13839;
   wire n13840;
   wire n13841;
   wire n13842;
   wire n13843;
   wire n13844;
   wire n13845;
   wire n13846;
   wire n13847;
   wire n13848;
   wire n13849;
   wire n13850;
   wire n13851;
   wire n13852;
   wire n13853;
   wire n13854;
   wire n13855;
   wire n13856;
   wire n13857;
   wire n13858;
   wire n13859;
   wire n13860;
   wire n13861;
   wire n13862;

   assign N18 = mem_access_addr[0] ;
   assign N19 = mem_access_addr[1] ;
   assign N20 = mem_access_addr[2] ;
   assign N21 = mem_access_addr[3] ;
   assign N22 = mem_access_addr[4] ;
   assign N23 = mem_access_addr[5] ;
   assign N24 = mem_access_addr[6] ;
   assign N25 = mem_access_addr[7] ;

   DFFHQX1 \ram_reg[253][15]  (.Q(\ram[253][15] ), 
	.D(n4645), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][14]  (.Q(\ram[253][14] ), 
	.D(n4644), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][13]  (.Q(\ram[253][13] ), 
	.D(n4643), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][12]  (.Q(\ram[253][12] ), 
	.D(n4642), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][11]  (.Q(\ram[253][11] ), 
	.D(n4641), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][10]  (.Q(\ram[253][10] ), 
	.D(n4640), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][9]  (.Q(\ram[253][9] ), 
	.D(n4639), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][8]  (.Q(\ram[253][8] ), 
	.D(n4638), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][7]  (.Q(\ram[253][7] ), 
	.D(n4637), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][6]  (.Q(\ram[253][6] ), 
	.D(n4636), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][5]  (.Q(\ram[253][5] ), 
	.D(n4635), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][4]  (.Q(\ram[253][4] ), 
	.D(n4634), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][3]  (.Q(\ram[253][3] ), 
	.D(n4633), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][2]  (.Q(\ram[253][2] ), 
	.D(n4632), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][1]  (.Q(\ram[253][1] ), 
	.D(n4631), 
	.CK(clk));
   DFFHQX1 \ram_reg[253][0]  (.Q(\ram[253][0] ), 
	.D(n4630), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][15]  (.Q(\ram[249][15] ), 
	.D(n4581), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][14]  (.Q(\ram[249][14] ), 
	.D(n4580), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][13]  (.Q(\ram[249][13] ), 
	.D(n4579), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][12]  (.Q(\ram[249][12] ), 
	.D(n4578), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][11]  (.Q(\ram[249][11] ), 
	.D(n4577), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][10]  (.Q(\ram[249][10] ), 
	.D(n4576), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][9]  (.Q(\ram[249][9] ), 
	.D(n4575), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][8]  (.Q(\ram[249][8] ), 
	.D(n4574), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][7]  (.Q(\ram[249][7] ), 
	.D(n4573), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][6]  (.Q(\ram[249][6] ), 
	.D(n4572), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][5]  (.Q(\ram[249][5] ), 
	.D(n4571), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][4]  (.Q(\ram[249][4] ), 
	.D(n4570), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][3]  (.Q(\ram[249][3] ), 
	.D(n4569), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][2]  (.Q(\ram[249][2] ), 
	.D(n4568), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][1]  (.Q(\ram[249][1] ), 
	.D(n4567), 
	.CK(clk));
   DFFHQX1 \ram_reg[249][0]  (.Q(\ram[249][0] ), 
	.D(n4566), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][15]  (.Q(\ram[245][15] ), 
	.D(n4517), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][14]  (.Q(\ram[245][14] ), 
	.D(n4516), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][13]  (.Q(\ram[245][13] ), 
	.D(n4515), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][12]  (.Q(\ram[245][12] ), 
	.D(n4514), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][11]  (.Q(\ram[245][11] ), 
	.D(n4513), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][10]  (.Q(\ram[245][10] ), 
	.D(n4512), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][9]  (.Q(\ram[245][9] ), 
	.D(n4511), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][8]  (.Q(\ram[245][8] ), 
	.D(n4510), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][7]  (.Q(\ram[245][7] ), 
	.D(n4509), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][6]  (.Q(\ram[245][6] ), 
	.D(n4508), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][5]  (.Q(\ram[245][5] ), 
	.D(n4507), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][4]  (.Q(\ram[245][4] ), 
	.D(n4506), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][3]  (.Q(\ram[245][3] ), 
	.D(n4505), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][2]  (.Q(\ram[245][2] ), 
	.D(n4504), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][1]  (.Q(\ram[245][1] ), 
	.D(n4503), 
	.CK(clk));
   DFFHQX1 \ram_reg[245][0]  (.Q(\ram[245][0] ), 
	.D(n4502), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][15]  (.Q(\ram[241][15] ), 
	.D(n4453), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][14]  (.Q(\ram[241][14] ), 
	.D(n4452), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][13]  (.Q(\ram[241][13] ), 
	.D(n4451), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][12]  (.Q(\ram[241][12] ), 
	.D(n4450), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][11]  (.Q(\ram[241][11] ), 
	.D(n4449), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][10]  (.Q(\ram[241][10] ), 
	.D(n4448), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][9]  (.Q(\ram[241][9] ), 
	.D(n4447), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][8]  (.Q(\ram[241][8] ), 
	.D(n4446), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][7]  (.Q(\ram[241][7] ), 
	.D(n4445), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][6]  (.Q(\ram[241][6] ), 
	.D(n4444), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][5]  (.Q(\ram[241][5] ), 
	.D(n4443), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][4]  (.Q(\ram[241][4] ), 
	.D(n4442), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][3]  (.Q(\ram[241][3] ), 
	.D(n4441), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][2]  (.Q(\ram[241][2] ), 
	.D(n4440), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][1]  (.Q(\ram[241][1] ), 
	.D(n4439), 
	.CK(clk));
   DFFHQX1 \ram_reg[241][0]  (.Q(\ram[241][0] ), 
	.D(n4438), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][15]  (.Q(\ram[237][15] ), 
	.D(n4389), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][14]  (.Q(\ram[237][14] ), 
	.D(n4388), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][13]  (.Q(\ram[237][13] ), 
	.D(n4387), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][12]  (.Q(\ram[237][12] ), 
	.D(n4386), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][11]  (.Q(\ram[237][11] ), 
	.D(n4385), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][10]  (.Q(\ram[237][10] ), 
	.D(n4384), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][9]  (.Q(\ram[237][9] ), 
	.D(n4383), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][8]  (.Q(\ram[237][8] ), 
	.D(n4382), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][7]  (.Q(\ram[237][7] ), 
	.D(n4381), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][6]  (.Q(\ram[237][6] ), 
	.D(n4380), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][5]  (.Q(\ram[237][5] ), 
	.D(n4379), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][4]  (.Q(\ram[237][4] ), 
	.D(n4378), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][3]  (.Q(\ram[237][3] ), 
	.D(n4377), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][2]  (.Q(\ram[237][2] ), 
	.D(n4376), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][1]  (.Q(\ram[237][1] ), 
	.D(n4375), 
	.CK(clk));
   DFFHQX1 \ram_reg[237][0]  (.Q(\ram[237][0] ), 
	.D(n4374), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][15]  (.Q(\ram[233][15] ), 
	.D(n4325), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][14]  (.Q(\ram[233][14] ), 
	.D(n4324), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][13]  (.Q(\ram[233][13] ), 
	.D(n4323), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][12]  (.Q(\ram[233][12] ), 
	.D(n4322), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][11]  (.Q(\ram[233][11] ), 
	.D(n4321), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][10]  (.Q(\ram[233][10] ), 
	.D(n4320), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][9]  (.Q(\ram[233][9] ), 
	.D(n4319), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][8]  (.Q(\ram[233][8] ), 
	.D(n4318), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][7]  (.Q(\ram[233][7] ), 
	.D(n4317), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][6]  (.Q(\ram[233][6] ), 
	.D(n4316), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][5]  (.Q(\ram[233][5] ), 
	.D(n4315), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][4]  (.Q(\ram[233][4] ), 
	.D(n4314), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][3]  (.Q(\ram[233][3] ), 
	.D(n4313), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][2]  (.Q(\ram[233][2] ), 
	.D(n4312), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][1]  (.Q(\ram[233][1] ), 
	.D(n4311), 
	.CK(clk));
   DFFHQX1 \ram_reg[233][0]  (.Q(\ram[233][0] ), 
	.D(n4310), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][15]  (.Q(\ram[229][15] ), 
	.D(n4261), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][14]  (.Q(\ram[229][14] ), 
	.D(n4260), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][13]  (.Q(\ram[229][13] ), 
	.D(n4259), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][12]  (.Q(\ram[229][12] ), 
	.D(n4258), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][11]  (.Q(\ram[229][11] ), 
	.D(n4257), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][10]  (.Q(\ram[229][10] ), 
	.D(n4256), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][9]  (.Q(\ram[229][9] ), 
	.D(n4255), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][8]  (.Q(\ram[229][8] ), 
	.D(n4254), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][7]  (.Q(\ram[229][7] ), 
	.D(n4253), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][6]  (.Q(\ram[229][6] ), 
	.D(n4252), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][5]  (.Q(\ram[229][5] ), 
	.D(n4251), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][4]  (.Q(\ram[229][4] ), 
	.D(n4250), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][3]  (.Q(\ram[229][3] ), 
	.D(n4249), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][2]  (.Q(\ram[229][2] ), 
	.D(n4248), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][1]  (.Q(\ram[229][1] ), 
	.D(n4247), 
	.CK(clk));
   DFFHQX1 \ram_reg[229][0]  (.Q(\ram[229][0] ), 
	.D(n4246), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][15]  (.Q(\ram[225][15] ), 
	.D(n4197), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][14]  (.Q(\ram[225][14] ), 
	.D(n4196), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][13]  (.Q(\ram[225][13] ), 
	.D(n4195), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][12]  (.Q(\ram[225][12] ), 
	.D(n4194), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][11]  (.Q(\ram[225][11] ), 
	.D(n4193), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][10]  (.Q(\ram[225][10] ), 
	.D(n4192), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][9]  (.Q(\ram[225][9] ), 
	.D(n4191), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][8]  (.Q(\ram[225][8] ), 
	.D(n4190), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][7]  (.Q(\ram[225][7] ), 
	.D(n4189), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][6]  (.Q(\ram[225][6] ), 
	.D(n4188), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][5]  (.Q(\ram[225][5] ), 
	.D(n4187), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][4]  (.Q(\ram[225][4] ), 
	.D(n4186), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][3]  (.Q(\ram[225][3] ), 
	.D(n4185), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][2]  (.Q(\ram[225][2] ), 
	.D(n4184), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][1]  (.Q(\ram[225][1] ), 
	.D(n4183), 
	.CK(clk));
   DFFHQX1 \ram_reg[225][0]  (.Q(\ram[225][0] ), 
	.D(n4182), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][15]  (.Q(\ram[221][15] ), 
	.D(n4133), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][14]  (.Q(\ram[221][14] ), 
	.D(n4132), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][13]  (.Q(\ram[221][13] ), 
	.D(n4131), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][12]  (.Q(\ram[221][12] ), 
	.D(n4130), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][11]  (.Q(\ram[221][11] ), 
	.D(n4129), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][10]  (.Q(\ram[221][10] ), 
	.D(n4128), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][9]  (.Q(\ram[221][9] ), 
	.D(n4127), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][8]  (.Q(\ram[221][8] ), 
	.D(n4126), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][7]  (.Q(\ram[221][7] ), 
	.D(n4125), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][6]  (.Q(\ram[221][6] ), 
	.D(n4124), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][5]  (.Q(\ram[221][5] ), 
	.D(n4123), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][4]  (.Q(\ram[221][4] ), 
	.D(n4122), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][3]  (.Q(\ram[221][3] ), 
	.D(n4121), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][2]  (.Q(\ram[221][2] ), 
	.D(n4120), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][1]  (.Q(\ram[221][1] ), 
	.D(n4119), 
	.CK(clk));
   DFFHQX1 \ram_reg[221][0]  (.Q(\ram[221][0] ), 
	.D(n4118), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][15]  (.Q(\ram[217][15] ), 
	.D(n4069), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][14]  (.Q(\ram[217][14] ), 
	.D(n4068), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][13]  (.Q(\ram[217][13] ), 
	.D(n4067), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][12]  (.Q(\ram[217][12] ), 
	.D(n4066), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][11]  (.Q(\ram[217][11] ), 
	.D(n4065), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][10]  (.Q(\ram[217][10] ), 
	.D(n4064), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][9]  (.Q(\ram[217][9] ), 
	.D(n4063), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][8]  (.Q(\ram[217][8] ), 
	.D(n4062), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][7]  (.Q(\ram[217][7] ), 
	.D(n4061), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][6]  (.Q(\ram[217][6] ), 
	.D(n4060), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][5]  (.Q(\ram[217][5] ), 
	.D(n4059), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][4]  (.Q(\ram[217][4] ), 
	.D(n4058), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][3]  (.Q(\ram[217][3] ), 
	.D(n4057), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][2]  (.Q(\ram[217][2] ), 
	.D(n4056), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][1]  (.Q(\ram[217][1] ), 
	.D(n4055), 
	.CK(clk));
   DFFHQX1 \ram_reg[217][0]  (.Q(\ram[217][0] ), 
	.D(n4054), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][15]  (.Q(\ram[213][15] ), 
	.D(n4005), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][14]  (.Q(\ram[213][14] ), 
	.D(n4004), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][13]  (.Q(\ram[213][13] ), 
	.D(n4003), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][12]  (.Q(\ram[213][12] ), 
	.D(n4002), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][11]  (.Q(\ram[213][11] ), 
	.D(n4001), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][10]  (.Q(\ram[213][10] ), 
	.D(n4000), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][9]  (.Q(\ram[213][9] ), 
	.D(n3999), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][8]  (.Q(\ram[213][8] ), 
	.D(n3998), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][7]  (.Q(\ram[213][7] ), 
	.D(n3997), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][6]  (.Q(\ram[213][6] ), 
	.D(n3996), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][5]  (.Q(\ram[213][5] ), 
	.D(n3995), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][4]  (.Q(\ram[213][4] ), 
	.D(n3994), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][3]  (.Q(\ram[213][3] ), 
	.D(n3993), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][2]  (.Q(\ram[213][2] ), 
	.D(n3992), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][1]  (.Q(\ram[213][1] ), 
	.D(n3991), 
	.CK(clk));
   DFFHQX1 \ram_reg[213][0]  (.Q(\ram[213][0] ), 
	.D(n3990), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][15]  (.Q(\ram[209][15] ), 
	.D(n3941), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][14]  (.Q(\ram[209][14] ), 
	.D(n3940), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][13]  (.Q(\ram[209][13] ), 
	.D(n3939), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][12]  (.Q(\ram[209][12] ), 
	.D(n3938), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][11]  (.Q(\ram[209][11] ), 
	.D(n3937), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][10]  (.Q(\ram[209][10] ), 
	.D(n3936), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][9]  (.Q(\ram[209][9] ), 
	.D(n3935), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][8]  (.Q(\ram[209][8] ), 
	.D(n3934), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][7]  (.Q(\ram[209][7] ), 
	.D(n3933), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][6]  (.Q(\ram[209][6] ), 
	.D(n3932), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][5]  (.Q(\ram[209][5] ), 
	.D(n3931), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][4]  (.Q(\ram[209][4] ), 
	.D(n3930), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][3]  (.Q(\ram[209][3] ), 
	.D(n3929), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][2]  (.Q(\ram[209][2] ), 
	.D(n3928), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][1]  (.Q(\ram[209][1] ), 
	.D(n3927), 
	.CK(clk));
   DFFHQX1 \ram_reg[209][0]  (.Q(\ram[209][0] ), 
	.D(n3926), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][15]  (.Q(\ram[205][15] ), 
	.D(n3877), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][14]  (.Q(\ram[205][14] ), 
	.D(n3876), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][13]  (.Q(\ram[205][13] ), 
	.D(n3875), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][12]  (.Q(\ram[205][12] ), 
	.D(n3874), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][11]  (.Q(\ram[205][11] ), 
	.D(n3873), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][10]  (.Q(\ram[205][10] ), 
	.D(n3872), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][9]  (.Q(\ram[205][9] ), 
	.D(n3871), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][8]  (.Q(\ram[205][8] ), 
	.D(n3870), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][7]  (.Q(\ram[205][7] ), 
	.D(n3869), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][6]  (.Q(\ram[205][6] ), 
	.D(n3868), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][5]  (.Q(\ram[205][5] ), 
	.D(n3867), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][4]  (.Q(\ram[205][4] ), 
	.D(n3866), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][3]  (.Q(\ram[205][3] ), 
	.D(n3865), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][2]  (.Q(\ram[205][2] ), 
	.D(n3864), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][1]  (.Q(\ram[205][1] ), 
	.D(n3863), 
	.CK(clk));
   DFFHQX1 \ram_reg[205][0]  (.Q(\ram[205][0] ), 
	.D(n3862), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][15]  (.Q(\ram[201][15] ), 
	.D(n3813), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][14]  (.Q(\ram[201][14] ), 
	.D(n3812), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][13]  (.Q(\ram[201][13] ), 
	.D(n3811), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][12]  (.Q(\ram[201][12] ), 
	.D(n3810), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][11]  (.Q(\ram[201][11] ), 
	.D(n3809), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][10]  (.Q(\ram[201][10] ), 
	.D(n3808), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][9]  (.Q(\ram[201][9] ), 
	.D(n3807), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][8]  (.Q(\ram[201][8] ), 
	.D(n3806), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][7]  (.Q(\ram[201][7] ), 
	.D(n3805), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][6]  (.Q(\ram[201][6] ), 
	.D(n3804), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][5]  (.Q(\ram[201][5] ), 
	.D(n3803), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][4]  (.Q(\ram[201][4] ), 
	.D(n3802), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][3]  (.Q(\ram[201][3] ), 
	.D(n3801), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][2]  (.Q(\ram[201][2] ), 
	.D(n3800), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][1]  (.Q(\ram[201][1] ), 
	.D(n3799), 
	.CK(clk));
   DFFHQX1 \ram_reg[201][0]  (.Q(\ram[201][0] ), 
	.D(n3798), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][15]  (.Q(\ram[197][15] ), 
	.D(n3749), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][14]  (.Q(\ram[197][14] ), 
	.D(n3748), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][13]  (.Q(\ram[197][13] ), 
	.D(n3747), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][12]  (.Q(\ram[197][12] ), 
	.D(n3746), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][11]  (.Q(\ram[197][11] ), 
	.D(n3745), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][10]  (.Q(\ram[197][10] ), 
	.D(n3744), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][9]  (.Q(\ram[197][9] ), 
	.D(n3743), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][8]  (.Q(\ram[197][8] ), 
	.D(n3742), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][7]  (.Q(\ram[197][7] ), 
	.D(n3741), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][6]  (.Q(\ram[197][6] ), 
	.D(n3740), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][5]  (.Q(\ram[197][5] ), 
	.D(n3739), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][4]  (.Q(\ram[197][4] ), 
	.D(n3738), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][3]  (.Q(\ram[197][3] ), 
	.D(n3737), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][2]  (.Q(\ram[197][2] ), 
	.D(n3736), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][1]  (.Q(\ram[197][1] ), 
	.D(n3735), 
	.CK(clk));
   DFFHQX1 \ram_reg[197][0]  (.Q(\ram[197][0] ), 
	.D(n3734), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][15]  (.Q(\ram[193][15] ), 
	.D(n3685), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][14]  (.Q(\ram[193][14] ), 
	.D(n3684), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][13]  (.Q(\ram[193][13] ), 
	.D(n3683), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][12]  (.Q(\ram[193][12] ), 
	.D(n3682), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][11]  (.Q(\ram[193][11] ), 
	.D(n3681), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][10]  (.Q(\ram[193][10] ), 
	.D(n3680), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][9]  (.Q(\ram[193][9] ), 
	.D(n3679), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][8]  (.Q(\ram[193][8] ), 
	.D(n3678), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][7]  (.Q(\ram[193][7] ), 
	.D(n3677), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][6]  (.Q(\ram[193][6] ), 
	.D(n3676), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][5]  (.Q(\ram[193][5] ), 
	.D(n3675), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][4]  (.Q(\ram[193][4] ), 
	.D(n3674), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][3]  (.Q(\ram[193][3] ), 
	.D(n3673), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][2]  (.Q(\ram[193][2] ), 
	.D(n3672), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][1]  (.Q(\ram[193][1] ), 
	.D(n3671), 
	.CK(clk));
   DFFHQX1 \ram_reg[193][0]  (.Q(\ram[193][0] ), 
	.D(n3670), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][15]  (.Q(\ram[189][15] ), 
	.D(n3621), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][14]  (.Q(\ram[189][14] ), 
	.D(n3620), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][13]  (.Q(\ram[189][13] ), 
	.D(n3619), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][12]  (.Q(\ram[189][12] ), 
	.D(n3618), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][11]  (.Q(\ram[189][11] ), 
	.D(n3617), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][10]  (.Q(\ram[189][10] ), 
	.D(n3616), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][9]  (.Q(\ram[189][9] ), 
	.D(n3615), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][8]  (.Q(\ram[189][8] ), 
	.D(n3614), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][7]  (.Q(\ram[189][7] ), 
	.D(n3613), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][6]  (.Q(\ram[189][6] ), 
	.D(n3612), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][5]  (.Q(\ram[189][5] ), 
	.D(n3611), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][4]  (.Q(\ram[189][4] ), 
	.D(n3610), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][3]  (.Q(\ram[189][3] ), 
	.D(n3609), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][2]  (.Q(\ram[189][2] ), 
	.D(n3608), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][1]  (.Q(\ram[189][1] ), 
	.D(n3607), 
	.CK(clk));
   DFFHQX1 \ram_reg[189][0]  (.Q(\ram[189][0] ), 
	.D(n3606), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][15]  (.Q(\ram[185][15] ), 
	.D(n3557), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][14]  (.Q(\ram[185][14] ), 
	.D(n3556), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][13]  (.Q(\ram[185][13] ), 
	.D(n3555), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][12]  (.Q(\ram[185][12] ), 
	.D(n3554), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][11]  (.Q(\ram[185][11] ), 
	.D(n3553), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][10]  (.Q(\ram[185][10] ), 
	.D(n3552), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][9]  (.Q(\ram[185][9] ), 
	.D(n3551), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][8]  (.Q(\ram[185][8] ), 
	.D(n3550), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][7]  (.Q(\ram[185][7] ), 
	.D(n3549), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][6]  (.Q(\ram[185][6] ), 
	.D(n3548), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][5]  (.Q(\ram[185][5] ), 
	.D(n3547), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][4]  (.Q(\ram[185][4] ), 
	.D(n3546), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][3]  (.Q(\ram[185][3] ), 
	.D(n3545), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][2]  (.Q(\ram[185][2] ), 
	.D(n3544), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][1]  (.Q(\ram[185][1] ), 
	.D(n3543), 
	.CK(clk));
   DFFHQX1 \ram_reg[185][0]  (.Q(\ram[185][0] ), 
	.D(n3542), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][15]  (.Q(\ram[181][15] ), 
	.D(n3493), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][14]  (.Q(\ram[181][14] ), 
	.D(n3492), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][13]  (.Q(\ram[181][13] ), 
	.D(n3491), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][12]  (.Q(\ram[181][12] ), 
	.D(n3490), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][11]  (.Q(\ram[181][11] ), 
	.D(n3489), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][10]  (.Q(\ram[181][10] ), 
	.D(n3488), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][9]  (.Q(\ram[181][9] ), 
	.D(n3487), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][8]  (.Q(\ram[181][8] ), 
	.D(n3486), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][7]  (.Q(\ram[181][7] ), 
	.D(n3485), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][6]  (.Q(\ram[181][6] ), 
	.D(n3484), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][5]  (.Q(\ram[181][5] ), 
	.D(n3483), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][4]  (.Q(\ram[181][4] ), 
	.D(n3482), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][3]  (.Q(\ram[181][3] ), 
	.D(n3481), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][2]  (.Q(\ram[181][2] ), 
	.D(n3480), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][1]  (.Q(\ram[181][1] ), 
	.D(n3479), 
	.CK(clk));
   DFFHQX1 \ram_reg[181][0]  (.Q(\ram[181][0] ), 
	.D(n3478), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][15]  (.Q(\ram[177][15] ), 
	.D(n3429), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][14]  (.Q(\ram[177][14] ), 
	.D(n3428), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][13]  (.Q(\ram[177][13] ), 
	.D(n3427), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][12]  (.Q(\ram[177][12] ), 
	.D(n3426), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][11]  (.Q(\ram[177][11] ), 
	.D(n3425), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][10]  (.Q(\ram[177][10] ), 
	.D(n3424), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][9]  (.Q(\ram[177][9] ), 
	.D(n3423), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][8]  (.Q(\ram[177][8] ), 
	.D(n3422), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][7]  (.Q(\ram[177][7] ), 
	.D(n3421), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][6]  (.Q(\ram[177][6] ), 
	.D(n3420), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][5]  (.Q(\ram[177][5] ), 
	.D(n3419), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][4]  (.Q(\ram[177][4] ), 
	.D(n3418), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][3]  (.Q(\ram[177][3] ), 
	.D(n3417), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][2]  (.Q(\ram[177][2] ), 
	.D(n3416), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][1]  (.Q(\ram[177][1] ), 
	.D(n3415), 
	.CK(clk));
   DFFHQX1 \ram_reg[177][0]  (.Q(\ram[177][0] ), 
	.D(n3414), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][15]  (.Q(\ram[173][15] ), 
	.D(n3365), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][14]  (.Q(\ram[173][14] ), 
	.D(n3364), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][13]  (.Q(\ram[173][13] ), 
	.D(n3363), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][12]  (.Q(\ram[173][12] ), 
	.D(n3362), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][11]  (.Q(\ram[173][11] ), 
	.D(n3361), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][10]  (.Q(\ram[173][10] ), 
	.D(n3360), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][9]  (.Q(\ram[173][9] ), 
	.D(n3359), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][8]  (.Q(\ram[173][8] ), 
	.D(n3358), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][7]  (.Q(\ram[173][7] ), 
	.D(n3357), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][6]  (.Q(\ram[173][6] ), 
	.D(n3356), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][5]  (.Q(\ram[173][5] ), 
	.D(n3355), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][4]  (.Q(\ram[173][4] ), 
	.D(n3354), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][3]  (.Q(\ram[173][3] ), 
	.D(n3353), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][2]  (.Q(\ram[173][2] ), 
	.D(n3352), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][1]  (.Q(\ram[173][1] ), 
	.D(n3351), 
	.CK(clk));
   DFFHQX1 \ram_reg[173][0]  (.Q(\ram[173][0] ), 
	.D(n3350), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][15]  (.Q(\ram[169][15] ), 
	.D(n3301), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][14]  (.Q(\ram[169][14] ), 
	.D(n3300), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][13]  (.Q(\ram[169][13] ), 
	.D(n3299), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][12]  (.Q(\ram[169][12] ), 
	.D(n3298), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][11]  (.Q(\ram[169][11] ), 
	.D(n3297), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][10]  (.Q(\ram[169][10] ), 
	.D(n3296), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][9]  (.Q(\ram[169][9] ), 
	.D(n3295), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][8]  (.Q(\ram[169][8] ), 
	.D(n3294), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][7]  (.Q(\ram[169][7] ), 
	.D(n3293), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][6]  (.Q(\ram[169][6] ), 
	.D(n3292), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][5]  (.Q(\ram[169][5] ), 
	.D(n3291), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][4]  (.Q(\ram[169][4] ), 
	.D(n3290), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][3]  (.Q(\ram[169][3] ), 
	.D(n3289), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][2]  (.Q(\ram[169][2] ), 
	.D(n3288), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][1]  (.Q(\ram[169][1] ), 
	.D(n3287), 
	.CK(clk));
   DFFHQX1 \ram_reg[169][0]  (.Q(\ram[169][0] ), 
	.D(n3286), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][15]  (.Q(\ram[165][15] ), 
	.D(n3237), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][14]  (.Q(\ram[165][14] ), 
	.D(n3236), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][13]  (.Q(\ram[165][13] ), 
	.D(n3235), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][12]  (.Q(\ram[165][12] ), 
	.D(n3234), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][11]  (.Q(\ram[165][11] ), 
	.D(n3233), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][10]  (.Q(\ram[165][10] ), 
	.D(n3232), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][9]  (.Q(\ram[165][9] ), 
	.D(n3231), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][8]  (.Q(\ram[165][8] ), 
	.D(n3230), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][7]  (.Q(\ram[165][7] ), 
	.D(n3229), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][6]  (.Q(\ram[165][6] ), 
	.D(n3228), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][5]  (.Q(\ram[165][5] ), 
	.D(n3227), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][4]  (.Q(\ram[165][4] ), 
	.D(n3226), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][3]  (.Q(\ram[165][3] ), 
	.D(n3225), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][2]  (.Q(\ram[165][2] ), 
	.D(n3224), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][1]  (.Q(\ram[165][1] ), 
	.D(n3223), 
	.CK(clk));
   DFFHQX1 \ram_reg[165][0]  (.Q(\ram[165][0] ), 
	.D(n3222), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][15]  (.Q(\ram[161][15] ), 
	.D(n3173), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][14]  (.Q(\ram[161][14] ), 
	.D(n3172), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][13]  (.Q(\ram[161][13] ), 
	.D(n3171), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][12]  (.Q(\ram[161][12] ), 
	.D(n3170), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][11]  (.Q(\ram[161][11] ), 
	.D(n3169), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][10]  (.Q(\ram[161][10] ), 
	.D(n3168), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][9]  (.Q(\ram[161][9] ), 
	.D(n3167), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][8]  (.Q(\ram[161][8] ), 
	.D(n3166), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][7]  (.Q(\ram[161][7] ), 
	.D(n3165), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][6]  (.Q(\ram[161][6] ), 
	.D(n3164), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][5]  (.Q(\ram[161][5] ), 
	.D(n3163), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][4]  (.Q(\ram[161][4] ), 
	.D(n3162), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][3]  (.Q(\ram[161][3] ), 
	.D(n3161), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][2]  (.Q(\ram[161][2] ), 
	.D(n3160), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][1]  (.Q(\ram[161][1] ), 
	.D(n3159), 
	.CK(clk));
   DFFHQX1 \ram_reg[161][0]  (.Q(\ram[161][0] ), 
	.D(n3158), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][15]  (.Q(\ram[157][15] ), 
	.D(n3109), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][14]  (.Q(\ram[157][14] ), 
	.D(n3108), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][13]  (.Q(\ram[157][13] ), 
	.D(n3107), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][12]  (.Q(\ram[157][12] ), 
	.D(n3106), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][11]  (.Q(\ram[157][11] ), 
	.D(n3105), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][10]  (.Q(\ram[157][10] ), 
	.D(n3104), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][9]  (.Q(\ram[157][9] ), 
	.D(n3103), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][8]  (.Q(\ram[157][8] ), 
	.D(n3102), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][7]  (.Q(\ram[157][7] ), 
	.D(n3101), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][6]  (.Q(\ram[157][6] ), 
	.D(n3100), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][5]  (.Q(\ram[157][5] ), 
	.D(n3099), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][4]  (.Q(\ram[157][4] ), 
	.D(n3098), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][3]  (.Q(\ram[157][3] ), 
	.D(n3097), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][2]  (.Q(\ram[157][2] ), 
	.D(n3096), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][1]  (.Q(\ram[157][1] ), 
	.D(n3095), 
	.CK(clk));
   DFFHQX1 \ram_reg[157][0]  (.Q(\ram[157][0] ), 
	.D(n3094), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][15]  (.Q(\ram[153][15] ), 
	.D(n3045), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][14]  (.Q(\ram[153][14] ), 
	.D(n3044), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][13]  (.Q(\ram[153][13] ), 
	.D(n3043), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][12]  (.Q(\ram[153][12] ), 
	.D(n3042), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][11]  (.Q(\ram[153][11] ), 
	.D(n3041), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][10]  (.Q(\ram[153][10] ), 
	.D(n3040), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][9]  (.Q(\ram[153][9] ), 
	.D(n3039), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][8]  (.Q(\ram[153][8] ), 
	.D(n3038), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][7]  (.Q(\ram[153][7] ), 
	.D(n3037), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][6]  (.Q(\ram[153][6] ), 
	.D(n3036), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][5]  (.Q(\ram[153][5] ), 
	.D(n3035), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][4]  (.Q(\ram[153][4] ), 
	.D(n3034), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][3]  (.Q(\ram[153][3] ), 
	.D(n3033), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][2]  (.Q(\ram[153][2] ), 
	.D(n3032), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][1]  (.Q(\ram[153][1] ), 
	.D(n3031), 
	.CK(clk));
   DFFHQX1 \ram_reg[153][0]  (.Q(\ram[153][0] ), 
	.D(n3030), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][15]  (.Q(\ram[149][15] ), 
	.D(n2981), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][14]  (.Q(\ram[149][14] ), 
	.D(n2980), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][13]  (.Q(\ram[149][13] ), 
	.D(n2979), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][12]  (.Q(\ram[149][12] ), 
	.D(n2978), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][11]  (.Q(\ram[149][11] ), 
	.D(n2977), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][10]  (.Q(\ram[149][10] ), 
	.D(n2976), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][9]  (.Q(\ram[149][9] ), 
	.D(n2975), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][8]  (.Q(\ram[149][8] ), 
	.D(n2974), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][7]  (.Q(\ram[149][7] ), 
	.D(n2973), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][6]  (.Q(\ram[149][6] ), 
	.D(n2972), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][5]  (.Q(\ram[149][5] ), 
	.D(n2971), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][4]  (.Q(\ram[149][4] ), 
	.D(n2970), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][3]  (.Q(\ram[149][3] ), 
	.D(n2969), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][2]  (.Q(\ram[149][2] ), 
	.D(n2968), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][1]  (.Q(\ram[149][1] ), 
	.D(n2967), 
	.CK(clk));
   DFFHQX1 \ram_reg[149][0]  (.Q(\ram[149][0] ), 
	.D(n2966), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][15]  (.Q(\ram[145][15] ), 
	.D(n2917), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][14]  (.Q(\ram[145][14] ), 
	.D(n2916), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][13]  (.Q(\ram[145][13] ), 
	.D(n2915), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][12]  (.Q(\ram[145][12] ), 
	.D(n2914), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][11]  (.Q(\ram[145][11] ), 
	.D(n2913), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][10]  (.Q(\ram[145][10] ), 
	.D(n2912), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][9]  (.Q(\ram[145][9] ), 
	.D(n2911), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][8]  (.Q(\ram[145][8] ), 
	.D(n2910), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][7]  (.Q(\ram[145][7] ), 
	.D(n2909), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][6]  (.Q(\ram[145][6] ), 
	.D(n2908), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][5]  (.Q(\ram[145][5] ), 
	.D(n2907), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][4]  (.Q(\ram[145][4] ), 
	.D(n2906), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][3]  (.Q(\ram[145][3] ), 
	.D(n2905), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][2]  (.Q(\ram[145][2] ), 
	.D(n2904), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][1]  (.Q(\ram[145][1] ), 
	.D(n2903), 
	.CK(clk));
   DFFHQX1 \ram_reg[145][0]  (.Q(\ram[145][0] ), 
	.D(n2902), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][15]  (.Q(\ram[141][15] ), 
	.D(n2853), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][14]  (.Q(\ram[141][14] ), 
	.D(n2852), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][13]  (.Q(\ram[141][13] ), 
	.D(n2851), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][12]  (.Q(\ram[141][12] ), 
	.D(n2850), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][11]  (.Q(\ram[141][11] ), 
	.D(n2849), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][10]  (.Q(\ram[141][10] ), 
	.D(n2848), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][9]  (.Q(\ram[141][9] ), 
	.D(n2847), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][8]  (.Q(\ram[141][8] ), 
	.D(n2846), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][7]  (.Q(\ram[141][7] ), 
	.D(n2845), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][6]  (.Q(\ram[141][6] ), 
	.D(n2844), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][5]  (.Q(\ram[141][5] ), 
	.D(n2843), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][4]  (.Q(\ram[141][4] ), 
	.D(n2842), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][3]  (.Q(\ram[141][3] ), 
	.D(n2841), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][2]  (.Q(\ram[141][2] ), 
	.D(n2840), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][1]  (.Q(\ram[141][1] ), 
	.D(n2839), 
	.CK(clk));
   DFFHQX1 \ram_reg[141][0]  (.Q(\ram[141][0] ), 
	.D(n2838), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][15]  (.Q(\ram[137][15] ), 
	.D(n2789), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][14]  (.Q(\ram[137][14] ), 
	.D(n2788), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][13]  (.Q(\ram[137][13] ), 
	.D(n2787), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][12]  (.Q(\ram[137][12] ), 
	.D(n2786), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][11]  (.Q(\ram[137][11] ), 
	.D(n2785), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][10]  (.Q(\ram[137][10] ), 
	.D(n2784), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][9]  (.Q(\ram[137][9] ), 
	.D(n2783), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][8]  (.Q(\ram[137][8] ), 
	.D(n2782), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][7]  (.Q(\ram[137][7] ), 
	.D(n2781), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][6]  (.Q(\ram[137][6] ), 
	.D(n2780), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][5]  (.Q(\ram[137][5] ), 
	.D(n2779), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][4]  (.Q(\ram[137][4] ), 
	.D(n2778), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][3]  (.Q(\ram[137][3] ), 
	.D(n2777), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][2]  (.Q(\ram[137][2] ), 
	.D(n2776), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][1]  (.Q(\ram[137][1] ), 
	.D(n2775), 
	.CK(clk));
   DFFHQX1 \ram_reg[137][0]  (.Q(\ram[137][0] ), 
	.D(n2774), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][15]  (.Q(\ram[133][15] ), 
	.D(n2725), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][14]  (.Q(\ram[133][14] ), 
	.D(n2724), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][13]  (.Q(\ram[133][13] ), 
	.D(n2723), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][12]  (.Q(\ram[133][12] ), 
	.D(n2722), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][11]  (.Q(\ram[133][11] ), 
	.D(n2721), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][10]  (.Q(\ram[133][10] ), 
	.D(n2720), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][9]  (.Q(\ram[133][9] ), 
	.D(n2719), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][8]  (.Q(\ram[133][8] ), 
	.D(n2718), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][7]  (.Q(\ram[133][7] ), 
	.D(n2717), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][6]  (.Q(\ram[133][6] ), 
	.D(n2716), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][5]  (.Q(\ram[133][5] ), 
	.D(n2715), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][4]  (.Q(\ram[133][4] ), 
	.D(n2714), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][3]  (.Q(\ram[133][3] ), 
	.D(n2713), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][2]  (.Q(\ram[133][2] ), 
	.D(n2712), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][1]  (.Q(\ram[133][1] ), 
	.D(n2711), 
	.CK(clk));
   DFFHQX1 \ram_reg[133][0]  (.Q(\ram[133][0] ), 
	.D(n2710), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][15]  (.Q(\ram[129][15] ), 
	.D(n2661), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][14]  (.Q(\ram[129][14] ), 
	.D(n2660), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][13]  (.Q(\ram[129][13] ), 
	.D(n2659), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][12]  (.Q(\ram[129][12] ), 
	.D(n2658), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][11]  (.Q(\ram[129][11] ), 
	.D(n2657), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][10]  (.Q(\ram[129][10] ), 
	.D(n2656), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][9]  (.Q(\ram[129][9] ), 
	.D(n2655), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][8]  (.Q(\ram[129][8] ), 
	.D(n2654), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][7]  (.Q(\ram[129][7] ), 
	.D(n2653), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][6]  (.Q(\ram[129][6] ), 
	.D(n2652), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][5]  (.Q(\ram[129][5] ), 
	.D(n2651), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][4]  (.Q(\ram[129][4] ), 
	.D(n2650), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][3]  (.Q(\ram[129][3] ), 
	.D(n2649), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][2]  (.Q(\ram[129][2] ), 
	.D(n2648), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][1]  (.Q(\ram[129][1] ), 
	.D(n2647), 
	.CK(clk));
   DFFHQX1 \ram_reg[129][0]  (.Q(\ram[129][0] ), 
	.D(n2646), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][15]  (.Q(\ram[125][15] ), 
	.D(n2597), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][14]  (.Q(\ram[125][14] ), 
	.D(n2596), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][13]  (.Q(\ram[125][13] ), 
	.D(n2595), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][12]  (.Q(\ram[125][12] ), 
	.D(n2594), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][11]  (.Q(\ram[125][11] ), 
	.D(n2593), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][10]  (.Q(\ram[125][10] ), 
	.D(n2592), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][9]  (.Q(\ram[125][9] ), 
	.D(n2591), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][8]  (.Q(\ram[125][8] ), 
	.D(n2590), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][7]  (.Q(\ram[125][7] ), 
	.D(n2589), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][6]  (.Q(\ram[125][6] ), 
	.D(n2588), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][5]  (.Q(\ram[125][5] ), 
	.D(n2587), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][4]  (.Q(\ram[125][4] ), 
	.D(n2586), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][3]  (.Q(\ram[125][3] ), 
	.D(n2585), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][2]  (.Q(\ram[125][2] ), 
	.D(n2584), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][1]  (.Q(\ram[125][1] ), 
	.D(n2583), 
	.CK(clk));
   DFFHQX1 \ram_reg[125][0]  (.Q(\ram[125][0] ), 
	.D(n2582), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][15]  (.Q(\ram[121][15] ), 
	.D(n2533), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][14]  (.Q(\ram[121][14] ), 
	.D(n2532), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][13]  (.Q(\ram[121][13] ), 
	.D(n2531), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][12]  (.Q(\ram[121][12] ), 
	.D(n2530), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][11]  (.Q(\ram[121][11] ), 
	.D(n2529), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][10]  (.Q(\ram[121][10] ), 
	.D(n2528), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][9]  (.Q(\ram[121][9] ), 
	.D(n2527), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][8]  (.Q(\ram[121][8] ), 
	.D(n2526), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][7]  (.Q(\ram[121][7] ), 
	.D(n2525), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][6]  (.Q(\ram[121][6] ), 
	.D(n2524), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][5]  (.Q(\ram[121][5] ), 
	.D(n2523), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][4]  (.Q(\ram[121][4] ), 
	.D(n2522), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][3]  (.Q(\ram[121][3] ), 
	.D(n2521), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][2]  (.Q(\ram[121][2] ), 
	.D(n2520), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][1]  (.Q(\ram[121][1] ), 
	.D(n2519), 
	.CK(clk));
   DFFHQX1 \ram_reg[121][0]  (.Q(\ram[121][0] ), 
	.D(n2518), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][15]  (.Q(\ram[117][15] ), 
	.D(n2469), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][14]  (.Q(\ram[117][14] ), 
	.D(n2468), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][13]  (.Q(\ram[117][13] ), 
	.D(n2467), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][12]  (.Q(\ram[117][12] ), 
	.D(n2466), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][11]  (.Q(\ram[117][11] ), 
	.D(n2465), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][10]  (.Q(\ram[117][10] ), 
	.D(n2464), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][9]  (.Q(\ram[117][9] ), 
	.D(n2463), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][8]  (.Q(\ram[117][8] ), 
	.D(n2462), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][7]  (.Q(\ram[117][7] ), 
	.D(n2461), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][6]  (.Q(\ram[117][6] ), 
	.D(n2460), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][5]  (.Q(\ram[117][5] ), 
	.D(n2459), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][4]  (.Q(\ram[117][4] ), 
	.D(n2458), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][3]  (.Q(\ram[117][3] ), 
	.D(n2457), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][2]  (.Q(\ram[117][2] ), 
	.D(n2456), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][1]  (.Q(\ram[117][1] ), 
	.D(n2455), 
	.CK(clk));
   DFFHQX1 \ram_reg[117][0]  (.Q(\ram[117][0] ), 
	.D(n2454), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][15]  (.Q(\ram[113][15] ), 
	.D(n2405), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][14]  (.Q(\ram[113][14] ), 
	.D(n2404), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][13]  (.Q(\ram[113][13] ), 
	.D(n2403), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][12]  (.Q(\ram[113][12] ), 
	.D(n2402), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][11]  (.Q(\ram[113][11] ), 
	.D(n2401), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][10]  (.Q(\ram[113][10] ), 
	.D(n2400), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][9]  (.Q(\ram[113][9] ), 
	.D(n2399), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][8]  (.Q(\ram[113][8] ), 
	.D(n2398), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][7]  (.Q(\ram[113][7] ), 
	.D(n2397), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][6]  (.Q(\ram[113][6] ), 
	.D(n2396), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][5]  (.Q(\ram[113][5] ), 
	.D(n2395), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][4]  (.Q(\ram[113][4] ), 
	.D(n2394), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][3]  (.Q(\ram[113][3] ), 
	.D(n2393), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][2]  (.Q(\ram[113][2] ), 
	.D(n2392), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][1]  (.Q(\ram[113][1] ), 
	.D(n2391), 
	.CK(clk));
   DFFHQX1 \ram_reg[113][0]  (.Q(\ram[113][0] ), 
	.D(n2390), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][15]  (.Q(\ram[109][15] ), 
	.D(n2341), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][14]  (.Q(\ram[109][14] ), 
	.D(n2340), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][13]  (.Q(\ram[109][13] ), 
	.D(n2339), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][12]  (.Q(\ram[109][12] ), 
	.D(n2338), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][11]  (.Q(\ram[109][11] ), 
	.D(n2337), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][10]  (.Q(\ram[109][10] ), 
	.D(n2336), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][9]  (.Q(\ram[109][9] ), 
	.D(n2335), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][8]  (.Q(\ram[109][8] ), 
	.D(n2334), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][7]  (.Q(\ram[109][7] ), 
	.D(n2333), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][6]  (.Q(\ram[109][6] ), 
	.D(n2332), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][5]  (.Q(\ram[109][5] ), 
	.D(n2331), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][4]  (.Q(\ram[109][4] ), 
	.D(n2330), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][3]  (.Q(\ram[109][3] ), 
	.D(n2329), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][2]  (.Q(\ram[109][2] ), 
	.D(n2328), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][1]  (.Q(\ram[109][1] ), 
	.D(n2327), 
	.CK(clk));
   DFFHQX1 \ram_reg[109][0]  (.Q(\ram[109][0] ), 
	.D(n2326), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][15]  (.Q(\ram[105][15] ), 
	.D(n2277), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][14]  (.Q(\ram[105][14] ), 
	.D(n2276), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][13]  (.Q(\ram[105][13] ), 
	.D(n2275), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][12]  (.Q(\ram[105][12] ), 
	.D(n2274), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][11]  (.Q(\ram[105][11] ), 
	.D(n2273), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][10]  (.Q(\ram[105][10] ), 
	.D(n2272), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][9]  (.Q(\ram[105][9] ), 
	.D(n2271), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][8]  (.Q(\ram[105][8] ), 
	.D(n2270), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][7]  (.Q(\ram[105][7] ), 
	.D(n2269), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][6]  (.Q(\ram[105][6] ), 
	.D(n2268), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][5]  (.Q(\ram[105][5] ), 
	.D(n2267), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][4]  (.Q(\ram[105][4] ), 
	.D(n2266), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][3]  (.Q(\ram[105][3] ), 
	.D(n2265), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][2]  (.Q(\ram[105][2] ), 
	.D(n2264), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][1]  (.Q(\ram[105][1] ), 
	.D(n2263), 
	.CK(clk));
   DFFHQX1 \ram_reg[105][0]  (.Q(\ram[105][0] ), 
	.D(n2262), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][15]  (.Q(\ram[101][15] ), 
	.D(n2213), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][14]  (.Q(\ram[101][14] ), 
	.D(n2212), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][13]  (.Q(\ram[101][13] ), 
	.D(n2211), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][12]  (.Q(\ram[101][12] ), 
	.D(n2210), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][11]  (.Q(\ram[101][11] ), 
	.D(n2209), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][10]  (.Q(\ram[101][10] ), 
	.D(n2208), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][9]  (.Q(\ram[101][9] ), 
	.D(n2207), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][8]  (.Q(\ram[101][8] ), 
	.D(n2206), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][7]  (.Q(\ram[101][7] ), 
	.D(n2205), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][6]  (.Q(\ram[101][6] ), 
	.D(n2204), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][5]  (.Q(\ram[101][5] ), 
	.D(n2203), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][4]  (.Q(\ram[101][4] ), 
	.D(n2202), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][3]  (.Q(\ram[101][3] ), 
	.D(n2201), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][2]  (.Q(\ram[101][2] ), 
	.D(n2200), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][1]  (.Q(\ram[101][1] ), 
	.D(n2199), 
	.CK(clk));
   DFFHQX1 \ram_reg[101][0]  (.Q(\ram[101][0] ), 
	.D(n2198), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][15]  (.Q(\ram[97][15] ), 
	.D(n2149), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][14]  (.Q(\ram[97][14] ), 
	.D(n2148), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][13]  (.Q(\ram[97][13] ), 
	.D(n2147), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][12]  (.Q(\ram[97][12] ), 
	.D(n2146), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][11]  (.Q(\ram[97][11] ), 
	.D(n2145), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][10]  (.Q(\ram[97][10] ), 
	.D(n2144), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][9]  (.Q(\ram[97][9] ), 
	.D(n2143), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][8]  (.Q(\ram[97][8] ), 
	.D(n2142), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][7]  (.Q(\ram[97][7] ), 
	.D(n2141), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][6]  (.Q(\ram[97][6] ), 
	.D(n2140), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][5]  (.Q(\ram[97][5] ), 
	.D(n2139), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][4]  (.Q(\ram[97][4] ), 
	.D(n2138), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][3]  (.Q(\ram[97][3] ), 
	.D(n2137), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][2]  (.Q(\ram[97][2] ), 
	.D(n2136), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][1]  (.Q(\ram[97][1] ), 
	.D(n2135), 
	.CK(clk));
   DFFHQX1 \ram_reg[97][0]  (.Q(\ram[97][0] ), 
	.D(n2134), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][15]  (.Q(\ram[93][15] ), 
	.D(n2085), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][14]  (.Q(\ram[93][14] ), 
	.D(n2084), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][13]  (.Q(\ram[93][13] ), 
	.D(n2083), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][12]  (.Q(\ram[93][12] ), 
	.D(n2082), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][11]  (.Q(\ram[93][11] ), 
	.D(n2081), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][10]  (.Q(\ram[93][10] ), 
	.D(n2080), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][9]  (.Q(\ram[93][9] ), 
	.D(n2079), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][8]  (.Q(\ram[93][8] ), 
	.D(n2078), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][7]  (.Q(\ram[93][7] ), 
	.D(n2077), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][6]  (.Q(\ram[93][6] ), 
	.D(n2076), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][5]  (.Q(\ram[93][5] ), 
	.D(n2075), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][4]  (.Q(\ram[93][4] ), 
	.D(n2074), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][3]  (.Q(\ram[93][3] ), 
	.D(n2073), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][2]  (.Q(\ram[93][2] ), 
	.D(n2072), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][1]  (.Q(\ram[93][1] ), 
	.D(n2071), 
	.CK(clk));
   DFFHQX1 \ram_reg[93][0]  (.Q(\ram[93][0] ), 
	.D(n2070), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][15]  (.Q(\ram[89][15] ), 
	.D(n2021), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][14]  (.Q(\ram[89][14] ), 
	.D(n2020), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][13]  (.Q(\ram[89][13] ), 
	.D(n2019), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][12]  (.Q(\ram[89][12] ), 
	.D(n2018), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][11]  (.Q(\ram[89][11] ), 
	.D(n2017), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][10]  (.Q(\ram[89][10] ), 
	.D(n2016), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][9]  (.Q(\ram[89][9] ), 
	.D(n2015), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][8]  (.Q(\ram[89][8] ), 
	.D(n2014), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][7]  (.Q(\ram[89][7] ), 
	.D(n2013), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][6]  (.Q(\ram[89][6] ), 
	.D(n2012), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][5]  (.Q(\ram[89][5] ), 
	.D(n2011), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][4]  (.Q(\ram[89][4] ), 
	.D(n2010), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][3]  (.Q(\ram[89][3] ), 
	.D(n2009), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][2]  (.Q(\ram[89][2] ), 
	.D(n2008), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][1]  (.Q(\ram[89][1] ), 
	.D(n2007), 
	.CK(clk));
   DFFHQX1 \ram_reg[89][0]  (.Q(\ram[89][0] ), 
	.D(n2006), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][15]  (.Q(\ram[85][15] ), 
	.D(n1957), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][14]  (.Q(\ram[85][14] ), 
	.D(n1956), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][13]  (.Q(\ram[85][13] ), 
	.D(n1955), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][12]  (.Q(\ram[85][12] ), 
	.D(n1954), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][11]  (.Q(\ram[85][11] ), 
	.D(n1953), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][10]  (.Q(\ram[85][10] ), 
	.D(n1952), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][9]  (.Q(\ram[85][9] ), 
	.D(n1951), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][8]  (.Q(\ram[85][8] ), 
	.D(n1950), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][7]  (.Q(\ram[85][7] ), 
	.D(n1949), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][6]  (.Q(\ram[85][6] ), 
	.D(n1948), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][5]  (.Q(\ram[85][5] ), 
	.D(n1947), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][4]  (.Q(\ram[85][4] ), 
	.D(n1946), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][3]  (.Q(\ram[85][3] ), 
	.D(n1945), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][2]  (.Q(\ram[85][2] ), 
	.D(n1944), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][1]  (.Q(\ram[85][1] ), 
	.D(n1943), 
	.CK(clk));
   DFFHQX1 \ram_reg[85][0]  (.Q(\ram[85][0] ), 
	.D(n1942), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][15]  (.Q(\ram[81][15] ), 
	.D(n1893), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][14]  (.Q(\ram[81][14] ), 
	.D(n1892), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][13]  (.Q(\ram[81][13] ), 
	.D(n1891), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][12]  (.Q(\ram[81][12] ), 
	.D(n1890), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][11]  (.Q(\ram[81][11] ), 
	.D(n1889), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][10]  (.Q(\ram[81][10] ), 
	.D(n1888), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][9]  (.Q(\ram[81][9] ), 
	.D(n1887), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][8]  (.Q(\ram[81][8] ), 
	.D(n1886), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][7]  (.Q(\ram[81][7] ), 
	.D(n1885), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][6]  (.Q(\ram[81][6] ), 
	.D(n1884), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][5]  (.Q(\ram[81][5] ), 
	.D(n1883), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][4]  (.Q(\ram[81][4] ), 
	.D(n1882), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][3]  (.Q(\ram[81][3] ), 
	.D(n1881), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][2]  (.Q(\ram[81][2] ), 
	.D(n1880), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][1]  (.Q(\ram[81][1] ), 
	.D(n1879), 
	.CK(clk));
   DFFHQX1 \ram_reg[81][0]  (.Q(\ram[81][0] ), 
	.D(n1878), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][15]  (.Q(\ram[77][15] ), 
	.D(n1829), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][14]  (.Q(\ram[77][14] ), 
	.D(n1828), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][13]  (.Q(\ram[77][13] ), 
	.D(n1827), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][12]  (.Q(\ram[77][12] ), 
	.D(n1826), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][11]  (.Q(\ram[77][11] ), 
	.D(n1825), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][10]  (.Q(\ram[77][10] ), 
	.D(n1824), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][9]  (.Q(\ram[77][9] ), 
	.D(n1823), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][8]  (.Q(\ram[77][8] ), 
	.D(n1822), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][7]  (.Q(\ram[77][7] ), 
	.D(n1821), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][6]  (.Q(\ram[77][6] ), 
	.D(n1820), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][5]  (.Q(\ram[77][5] ), 
	.D(n1819), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][4]  (.Q(\ram[77][4] ), 
	.D(n1818), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][3]  (.Q(\ram[77][3] ), 
	.D(n1817), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][2]  (.Q(\ram[77][2] ), 
	.D(n1816), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][1]  (.Q(\ram[77][1] ), 
	.D(n1815), 
	.CK(clk));
   DFFHQX1 \ram_reg[77][0]  (.Q(\ram[77][0] ), 
	.D(n1814), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][15]  (.Q(\ram[73][15] ), 
	.D(n1765), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][14]  (.Q(\ram[73][14] ), 
	.D(n1764), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][13]  (.Q(\ram[73][13] ), 
	.D(n1763), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][12]  (.Q(\ram[73][12] ), 
	.D(n1762), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][11]  (.Q(\ram[73][11] ), 
	.D(n1761), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][10]  (.Q(\ram[73][10] ), 
	.D(n1760), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][9]  (.Q(\ram[73][9] ), 
	.D(n1759), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][8]  (.Q(\ram[73][8] ), 
	.D(n1758), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][7]  (.Q(\ram[73][7] ), 
	.D(n1757), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][6]  (.Q(\ram[73][6] ), 
	.D(n1756), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][5]  (.Q(\ram[73][5] ), 
	.D(n1755), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][4]  (.Q(\ram[73][4] ), 
	.D(n1754), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][3]  (.Q(\ram[73][3] ), 
	.D(n1753), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][2]  (.Q(\ram[73][2] ), 
	.D(n1752), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][1]  (.Q(\ram[73][1] ), 
	.D(n1751), 
	.CK(clk));
   DFFHQX1 \ram_reg[73][0]  (.Q(\ram[73][0] ), 
	.D(n1750), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][15]  (.Q(\ram[69][15] ), 
	.D(n1701), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][14]  (.Q(\ram[69][14] ), 
	.D(n1700), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][13]  (.Q(\ram[69][13] ), 
	.D(n1699), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][12]  (.Q(\ram[69][12] ), 
	.D(n1698), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][11]  (.Q(\ram[69][11] ), 
	.D(n1697), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][10]  (.Q(\ram[69][10] ), 
	.D(n1696), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][9]  (.Q(\ram[69][9] ), 
	.D(n1695), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][8]  (.Q(\ram[69][8] ), 
	.D(n1694), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][7]  (.Q(\ram[69][7] ), 
	.D(n1693), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][6]  (.Q(\ram[69][6] ), 
	.D(n1692), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][5]  (.Q(\ram[69][5] ), 
	.D(n1691), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][4]  (.Q(\ram[69][4] ), 
	.D(n1690), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][3]  (.Q(\ram[69][3] ), 
	.D(n1689), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][2]  (.Q(\ram[69][2] ), 
	.D(n1688), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][1]  (.Q(\ram[69][1] ), 
	.D(n1687), 
	.CK(clk));
   DFFHQX1 \ram_reg[69][0]  (.Q(\ram[69][0] ), 
	.D(n1686), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][15]  (.Q(\ram[65][15] ), 
	.D(n1637), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][14]  (.Q(\ram[65][14] ), 
	.D(n1636), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][13]  (.Q(\ram[65][13] ), 
	.D(n1635), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][12]  (.Q(\ram[65][12] ), 
	.D(n1634), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][11]  (.Q(\ram[65][11] ), 
	.D(n1633), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][10]  (.Q(\ram[65][10] ), 
	.D(n1632), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][9]  (.Q(\ram[65][9] ), 
	.D(n1631), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][8]  (.Q(\ram[65][8] ), 
	.D(n1630), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][7]  (.Q(\ram[65][7] ), 
	.D(n1629), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][6]  (.Q(\ram[65][6] ), 
	.D(n1628), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][5]  (.Q(\ram[65][5] ), 
	.D(n1627), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][4]  (.Q(\ram[65][4] ), 
	.D(n1626), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][3]  (.Q(\ram[65][3] ), 
	.D(n1625), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][2]  (.Q(\ram[65][2] ), 
	.D(n1624), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][1]  (.Q(\ram[65][1] ), 
	.D(n1623), 
	.CK(clk));
   DFFHQX1 \ram_reg[65][0]  (.Q(\ram[65][0] ), 
	.D(n1622), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][15]  (.Q(\ram[61][15] ), 
	.D(n1573), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][14]  (.Q(\ram[61][14] ), 
	.D(n1572), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][13]  (.Q(\ram[61][13] ), 
	.D(n1571), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][12]  (.Q(\ram[61][12] ), 
	.D(n1570), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][11]  (.Q(\ram[61][11] ), 
	.D(n1569), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][10]  (.Q(\ram[61][10] ), 
	.D(n1568), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][9]  (.Q(\ram[61][9] ), 
	.D(n1567), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][8]  (.Q(\ram[61][8] ), 
	.D(n1566), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][7]  (.Q(\ram[61][7] ), 
	.D(n1565), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][6]  (.Q(\ram[61][6] ), 
	.D(n1564), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][5]  (.Q(\ram[61][5] ), 
	.D(n1563), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][4]  (.Q(\ram[61][4] ), 
	.D(n1562), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][3]  (.Q(\ram[61][3] ), 
	.D(n1561), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][2]  (.Q(\ram[61][2] ), 
	.D(n1560), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][1]  (.Q(\ram[61][1] ), 
	.D(n1559), 
	.CK(clk));
   DFFHQX1 \ram_reg[61][0]  (.Q(\ram[61][0] ), 
	.D(n1558), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][15]  (.Q(\ram[57][15] ), 
	.D(n1509), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][14]  (.Q(\ram[57][14] ), 
	.D(n1508), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][13]  (.Q(\ram[57][13] ), 
	.D(n1507), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][12]  (.Q(\ram[57][12] ), 
	.D(n1506), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][11]  (.Q(\ram[57][11] ), 
	.D(n1505), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][10]  (.Q(\ram[57][10] ), 
	.D(n1504), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][9]  (.Q(\ram[57][9] ), 
	.D(n1503), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][8]  (.Q(\ram[57][8] ), 
	.D(n1502), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][7]  (.Q(\ram[57][7] ), 
	.D(n1501), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][6]  (.Q(\ram[57][6] ), 
	.D(n1500), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][5]  (.Q(\ram[57][5] ), 
	.D(n1499), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][4]  (.Q(\ram[57][4] ), 
	.D(n1498), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][3]  (.Q(\ram[57][3] ), 
	.D(n1497), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][2]  (.Q(\ram[57][2] ), 
	.D(n1496), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][1]  (.Q(\ram[57][1] ), 
	.D(n1495), 
	.CK(clk));
   DFFHQX1 \ram_reg[57][0]  (.Q(\ram[57][0] ), 
	.D(n1494), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][15]  (.Q(\ram[53][15] ), 
	.D(n1445), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][14]  (.Q(\ram[53][14] ), 
	.D(n1444), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][13]  (.Q(\ram[53][13] ), 
	.D(n1443), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][12]  (.Q(\ram[53][12] ), 
	.D(n1442), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][11]  (.Q(\ram[53][11] ), 
	.D(n1441), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][10]  (.Q(\ram[53][10] ), 
	.D(n1440), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][9]  (.Q(\ram[53][9] ), 
	.D(n1439), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][8]  (.Q(\ram[53][8] ), 
	.D(n1438), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][7]  (.Q(\ram[53][7] ), 
	.D(n1437), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][6]  (.Q(\ram[53][6] ), 
	.D(n1436), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][5]  (.Q(\ram[53][5] ), 
	.D(n1435), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][4]  (.Q(\ram[53][4] ), 
	.D(n1434), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][3]  (.Q(\ram[53][3] ), 
	.D(n1433), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][2]  (.Q(\ram[53][2] ), 
	.D(n1432), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][1]  (.Q(\ram[53][1] ), 
	.D(n1431), 
	.CK(clk));
   DFFHQX1 \ram_reg[53][0]  (.Q(\ram[53][0] ), 
	.D(n1430), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][15]  (.Q(\ram[49][15] ), 
	.D(n1381), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][14]  (.Q(\ram[49][14] ), 
	.D(n1380), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][13]  (.Q(\ram[49][13] ), 
	.D(n1379), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][12]  (.Q(\ram[49][12] ), 
	.D(n1378), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][11]  (.Q(\ram[49][11] ), 
	.D(n1377), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][10]  (.Q(\ram[49][10] ), 
	.D(n1376), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][9]  (.Q(\ram[49][9] ), 
	.D(n1375), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][8]  (.Q(\ram[49][8] ), 
	.D(n1374), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][7]  (.Q(\ram[49][7] ), 
	.D(n1373), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][6]  (.Q(\ram[49][6] ), 
	.D(n1372), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][5]  (.Q(\ram[49][5] ), 
	.D(n1371), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][4]  (.Q(\ram[49][4] ), 
	.D(n1370), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][3]  (.Q(\ram[49][3] ), 
	.D(n1369), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][2]  (.Q(\ram[49][2] ), 
	.D(n1368), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][1]  (.Q(\ram[49][1] ), 
	.D(n1367), 
	.CK(clk));
   DFFHQX1 \ram_reg[49][0]  (.Q(\ram[49][0] ), 
	.D(n1366), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][15]  (.Q(\ram[45][15] ), 
	.D(n1317), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][14]  (.Q(\ram[45][14] ), 
	.D(n1316), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][13]  (.Q(\ram[45][13] ), 
	.D(n1315), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][12]  (.Q(\ram[45][12] ), 
	.D(n1314), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][11]  (.Q(\ram[45][11] ), 
	.D(n1313), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][10]  (.Q(\ram[45][10] ), 
	.D(n1312), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][9]  (.Q(\ram[45][9] ), 
	.D(n1311), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][8]  (.Q(\ram[45][8] ), 
	.D(n1310), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][7]  (.Q(\ram[45][7] ), 
	.D(n1309), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][6]  (.Q(\ram[45][6] ), 
	.D(n1308), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][5]  (.Q(\ram[45][5] ), 
	.D(n1307), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][4]  (.Q(\ram[45][4] ), 
	.D(n1306), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][3]  (.Q(\ram[45][3] ), 
	.D(n1305), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][2]  (.Q(\ram[45][2] ), 
	.D(n1304), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][1]  (.Q(\ram[45][1] ), 
	.D(n1303), 
	.CK(clk));
   DFFHQX1 \ram_reg[45][0]  (.Q(\ram[45][0] ), 
	.D(n1302), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][15]  (.Q(\ram[41][15] ), 
	.D(n1253), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][14]  (.Q(\ram[41][14] ), 
	.D(n1252), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][13]  (.Q(\ram[41][13] ), 
	.D(n1251), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][12]  (.Q(\ram[41][12] ), 
	.D(n1250), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][11]  (.Q(\ram[41][11] ), 
	.D(n1249), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][10]  (.Q(\ram[41][10] ), 
	.D(n1248), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][9]  (.Q(\ram[41][9] ), 
	.D(n1247), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][8]  (.Q(\ram[41][8] ), 
	.D(n1246), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][7]  (.Q(\ram[41][7] ), 
	.D(n1245), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][6]  (.Q(\ram[41][6] ), 
	.D(n1244), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][5]  (.Q(\ram[41][5] ), 
	.D(n1243), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][4]  (.Q(\ram[41][4] ), 
	.D(n1242), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][3]  (.Q(\ram[41][3] ), 
	.D(n1241), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][2]  (.Q(\ram[41][2] ), 
	.D(n1240), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][1]  (.Q(\ram[41][1] ), 
	.D(n1239), 
	.CK(clk));
   DFFHQX1 \ram_reg[41][0]  (.Q(\ram[41][0] ), 
	.D(n1238), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][15]  (.Q(\ram[37][15] ), 
	.D(n1189), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][14]  (.Q(\ram[37][14] ), 
	.D(n1188), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][13]  (.Q(\ram[37][13] ), 
	.D(n1187), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][12]  (.Q(\ram[37][12] ), 
	.D(n1186), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][11]  (.Q(\ram[37][11] ), 
	.D(n1185), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][10]  (.Q(\ram[37][10] ), 
	.D(n1184), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][9]  (.Q(\ram[37][9] ), 
	.D(n1183), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][8]  (.Q(\ram[37][8] ), 
	.D(n1182), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][7]  (.Q(\ram[37][7] ), 
	.D(n1181), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][6]  (.Q(\ram[37][6] ), 
	.D(n1180), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][5]  (.Q(\ram[37][5] ), 
	.D(n1179), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][4]  (.Q(\ram[37][4] ), 
	.D(n1178), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][3]  (.Q(\ram[37][3] ), 
	.D(n1177), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][2]  (.Q(\ram[37][2] ), 
	.D(n1176), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][1]  (.Q(\ram[37][1] ), 
	.D(n1175), 
	.CK(clk));
   DFFHQX1 \ram_reg[37][0]  (.Q(\ram[37][0] ), 
	.D(n1174), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][15]  (.Q(\ram[33][15] ), 
	.D(n1125), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][14]  (.Q(\ram[33][14] ), 
	.D(n1124), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][13]  (.Q(\ram[33][13] ), 
	.D(n1123), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][12]  (.Q(\ram[33][12] ), 
	.D(n1122), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][11]  (.Q(\ram[33][11] ), 
	.D(n1121), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][10]  (.Q(\ram[33][10] ), 
	.D(n1120), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][9]  (.Q(\ram[33][9] ), 
	.D(n1119), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][8]  (.Q(\ram[33][8] ), 
	.D(n1118), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][7]  (.Q(\ram[33][7] ), 
	.D(n1117), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][6]  (.Q(\ram[33][6] ), 
	.D(n1116), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][5]  (.Q(\ram[33][5] ), 
	.D(n1115), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][4]  (.Q(\ram[33][4] ), 
	.D(n1114), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][3]  (.Q(\ram[33][3] ), 
	.D(n1113), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][2]  (.Q(\ram[33][2] ), 
	.D(n1112), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][1]  (.Q(\ram[33][1] ), 
	.D(n1111), 
	.CK(clk));
   DFFHQX1 \ram_reg[33][0]  (.Q(\ram[33][0] ), 
	.D(n1110), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][15]  (.Q(\ram[29][15] ), 
	.D(n1061), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][14]  (.Q(\ram[29][14] ), 
	.D(n1060), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][13]  (.Q(\ram[29][13] ), 
	.D(n1059), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][12]  (.Q(\ram[29][12] ), 
	.D(n1058), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][11]  (.Q(\ram[29][11] ), 
	.D(n1057), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][10]  (.Q(\ram[29][10] ), 
	.D(n1056), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][9]  (.Q(\ram[29][9] ), 
	.D(n1055), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][8]  (.Q(\ram[29][8] ), 
	.D(n1054), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][7]  (.Q(\ram[29][7] ), 
	.D(n1053), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][6]  (.Q(\ram[29][6] ), 
	.D(n1052), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][5]  (.Q(\ram[29][5] ), 
	.D(n1051), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][4]  (.Q(\ram[29][4] ), 
	.D(n1050), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][3]  (.Q(\ram[29][3] ), 
	.D(n1049), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][2]  (.Q(\ram[29][2] ), 
	.D(n1048), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][1]  (.Q(\ram[29][1] ), 
	.D(n1047), 
	.CK(clk));
   DFFHQX1 \ram_reg[29][0]  (.Q(\ram[29][0] ), 
	.D(n1046), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][15]  (.Q(\ram[25][15] ), 
	.D(n997), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][14]  (.Q(\ram[25][14] ), 
	.D(n996), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][13]  (.Q(\ram[25][13] ), 
	.D(n995), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][12]  (.Q(\ram[25][12] ), 
	.D(n994), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][11]  (.Q(\ram[25][11] ), 
	.D(n993), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][10]  (.Q(\ram[25][10] ), 
	.D(n992), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][9]  (.Q(\ram[25][9] ), 
	.D(n991), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][8]  (.Q(\ram[25][8] ), 
	.D(n990), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][7]  (.Q(\ram[25][7] ), 
	.D(n989), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][6]  (.Q(\ram[25][6] ), 
	.D(n988), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][5]  (.Q(\ram[25][5] ), 
	.D(n987), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][4]  (.Q(\ram[25][4] ), 
	.D(n986), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][3]  (.Q(\ram[25][3] ), 
	.D(n985), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][2]  (.Q(\ram[25][2] ), 
	.D(n984), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][1]  (.Q(\ram[25][1] ), 
	.D(n983), 
	.CK(clk));
   DFFHQX1 \ram_reg[25][0]  (.Q(\ram[25][0] ), 
	.D(n982), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][15]  (.Q(\ram[21][15] ), 
	.D(n933), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][14]  (.Q(\ram[21][14] ), 
	.D(n932), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][13]  (.Q(\ram[21][13] ), 
	.D(n931), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][12]  (.Q(\ram[21][12] ), 
	.D(n930), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][11]  (.Q(\ram[21][11] ), 
	.D(n929), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][10]  (.Q(\ram[21][10] ), 
	.D(n928), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][9]  (.Q(\ram[21][9] ), 
	.D(n927), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][8]  (.Q(\ram[21][8] ), 
	.D(n926), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][7]  (.Q(\ram[21][7] ), 
	.D(n925), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][6]  (.Q(\ram[21][6] ), 
	.D(n924), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][5]  (.Q(\ram[21][5] ), 
	.D(n923), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][4]  (.Q(\ram[21][4] ), 
	.D(n922), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][3]  (.Q(\ram[21][3] ), 
	.D(n921), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][2]  (.Q(\ram[21][2] ), 
	.D(n920), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][1]  (.Q(\ram[21][1] ), 
	.D(n919), 
	.CK(clk));
   DFFHQX1 \ram_reg[21][0]  (.Q(\ram[21][0] ), 
	.D(n918), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][15]  (.Q(\ram[17][15] ), 
	.D(n869), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][14]  (.Q(\ram[17][14] ), 
	.D(n868), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][13]  (.Q(\ram[17][13] ), 
	.D(n867), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][12]  (.Q(\ram[17][12] ), 
	.D(n866), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][11]  (.Q(\ram[17][11] ), 
	.D(n865), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][10]  (.Q(\ram[17][10] ), 
	.D(n864), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][9]  (.Q(\ram[17][9] ), 
	.D(n863), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][8]  (.Q(\ram[17][8] ), 
	.D(n862), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][7]  (.Q(\ram[17][7] ), 
	.D(n861), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][6]  (.Q(\ram[17][6] ), 
	.D(n860), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][5]  (.Q(\ram[17][5] ), 
	.D(n859), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][4]  (.Q(\ram[17][4] ), 
	.D(n858), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][3]  (.Q(\ram[17][3] ), 
	.D(n857), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][2]  (.Q(\ram[17][2] ), 
	.D(n856), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][1]  (.Q(\ram[17][1] ), 
	.D(n855), 
	.CK(clk));
   DFFHQX1 \ram_reg[17][0]  (.Q(\ram[17][0] ), 
	.D(n854), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][15]  (.Q(\ram[13][15] ), 
	.D(n805), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][14]  (.Q(\ram[13][14] ), 
	.D(n804), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][13]  (.Q(\ram[13][13] ), 
	.D(n803), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][12]  (.Q(\ram[13][12] ), 
	.D(n802), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][11]  (.Q(\ram[13][11] ), 
	.D(n801), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][10]  (.Q(\ram[13][10] ), 
	.D(n800), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][9]  (.Q(\ram[13][9] ), 
	.D(n799), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][8]  (.Q(\ram[13][8] ), 
	.D(n798), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][7]  (.Q(\ram[13][7] ), 
	.D(n797), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][6]  (.Q(\ram[13][6] ), 
	.D(n796), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][5]  (.Q(\ram[13][5] ), 
	.D(n795), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][4]  (.Q(\ram[13][4] ), 
	.D(n794), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][3]  (.Q(\ram[13][3] ), 
	.D(n793), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][2]  (.Q(\ram[13][2] ), 
	.D(n792), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][1]  (.Q(\ram[13][1] ), 
	.D(n791), 
	.CK(clk));
   DFFHQX1 \ram_reg[13][0]  (.Q(\ram[13][0] ), 
	.D(n790), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][15]  (.Q(\ram[9][15] ), 
	.D(n741), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][14]  (.Q(\ram[9][14] ), 
	.D(n740), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][13]  (.Q(\ram[9][13] ), 
	.D(n739), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][12]  (.Q(\ram[9][12] ), 
	.D(n738), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][11]  (.Q(\ram[9][11] ), 
	.D(n737), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][10]  (.Q(\ram[9][10] ), 
	.D(n736), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][9]  (.Q(\ram[9][9] ), 
	.D(n735), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][8]  (.Q(\ram[9][8] ), 
	.D(n734), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][7]  (.Q(\ram[9][7] ), 
	.D(n733), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][6]  (.Q(\ram[9][6] ), 
	.D(n732), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][5]  (.Q(\ram[9][5] ), 
	.D(n731), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][4]  (.Q(\ram[9][4] ), 
	.D(n730), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][3]  (.Q(\ram[9][3] ), 
	.D(n729), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][2]  (.Q(\ram[9][2] ), 
	.D(n728), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][1]  (.Q(\ram[9][1] ), 
	.D(n727), 
	.CK(clk));
   DFFHQX1 \ram_reg[9][0]  (.Q(\ram[9][0] ), 
	.D(n726), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][15]  (.Q(\ram[5][15] ), 
	.D(n677), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][14]  (.Q(\ram[5][14] ), 
	.D(n676), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][13]  (.Q(\ram[5][13] ), 
	.D(n675), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][12]  (.Q(\ram[5][12] ), 
	.D(n674), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][11]  (.Q(\ram[5][11] ), 
	.D(n673), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][10]  (.Q(\ram[5][10] ), 
	.D(n672), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][9]  (.Q(\ram[5][9] ), 
	.D(n671), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][8]  (.Q(\ram[5][8] ), 
	.D(n670), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][7]  (.Q(\ram[5][7] ), 
	.D(n669), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][6]  (.Q(\ram[5][6] ), 
	.D(n668), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][5]  (.Q(\ram[5][5] ), 
	.D(n667), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][4]  (.Q(\ram[5][4] ), 
	.D(n666), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][3]  (.Q(\ram[5][3] ), 
	.D(n665), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][2]  (.Q(\ram[5][2] ), 
	.D(n664), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][1]  (.Q(\ram[5][1] ), 
	.D(n663), 
	.CK(clk));
   DFFHQX1 \ram_reg[5][0]  (.Q(\ram[5][0] ), 
	.D(n662), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][15]  (.Q(\ram[1][15] ), 
	.D(n613), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][14]  (.Q(\ram[1][14] ), 
	.D(n612), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][13]  (.Q(\ram[1][13] ), 
	.D(n611), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][12]  (.Q(\ram[1][12] ), 
	.D(n610), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][11]  (.Q(\ram[1][11] ), 
	.D(n609), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][10]  (.Q(\ram[1][10] ), 
	.D(n608), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][9]  (.Q(\ram[1][9] ), 
	.D(n607), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][8]  (.Q(\ram[1][8] ), 
	.D(n606), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][7]  (.Q(\ram[1][7] ), 
	.D(n605), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][6]  (.Q(\ram[1][6] ), 
	.D(n604), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][5]  (.Q(\ram[1][5] ), 
	.D(n603), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][4]  (.Q(\ram[1][4] ), 
	.D(n602), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][3]  (.Q(\ram[1][3] ), 
	.D(n601), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][2]  (.Q(\ram[1][2] ), 
	.D(n600), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][1]  (.Q(\ram[1][1] ), 
	.D(n599), 
	.CK(clk));
   DFFHQX1 \ram_reg[1][0]  (.Q(\ram[1][0] ), 
	.D(n598), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][15]  (.Q(\ram[255][15] ), 
	.D(n4677), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][14]  (.Q(\ram[255][14] ), 
	.D(n4676), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][13]  (.Q(\ram[255][13] ), 
	.D(n4675), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][12]  (.Q(\ram[255][12] ), 
	.D(n4674), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][11]  (.Q(\ram[255][11] ), 
	.D(n4673), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][10]  (.Q(\ram[255][10] ), 
	.D(n4672), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][9]  (.Q(\ram[255][9] ), 
	.D(n4671), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][8]  (.Q(\ram[255][8] ), 
	.D(n4670), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][7]  (.Q(\ram[255][7] ), 
	.D(n4669), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][6]  (.Q(\ram[255][6] ), 
	.D(n4668), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][5]  (.Q(\ram[255][5] ), 
	.D(n4667), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][4]  (.Q(\ram[255][4] ), 
	.D(n4666), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][3]  (.Q(\ram[255][3] ), 
	.D(n4665), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][2]  (.Q(\ram[255][2] ), 
	.D(n4664), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][1]  (.Q(\ram[255][1] ), 
	.D(n4663), 
	.CK(clk));
   DFFHQX1 \ram_reg[255][0]  (.Q(\ram[255][0] ), 
	.D(n4662), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][15]  (.Q(\ram[251][15] ), 
	.D(n4613), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][14]  (.Q(\ram[251][14] ), 
	.D(n4612), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][13]  (.Q(\ram[251][13] ), 
	.D(n4611), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][12]  (.Q(\ram[251][12] ), 
	.D(n4610), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][11]  (.Q(\ram[251][11] ), 
	.D(n4609), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][10]  (.Q(\ram[251][10] ), 
	.D(n4608), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][9]  (.Q(\ram[251][9] ), 
	.D(n4607), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][8]  (.Q(\ram[251][8] ), 
	.D(n4606), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][7]  (.Q(\ram[251][7] ), 
	.D(n4605), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][6]  (.Q(\ram[251][6] ), 
	.D(n4604), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][5]  (.Q(\ram[251][5] ), 
	.D(n4603), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][4]  (.Q(\ram[251][4] ), 
	.D(n4602), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][3]  (.Q(\ram[251][3] ), 
	.D(n4601), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][2]  (.Q(\ram[251][2] ), 
	.D(n4600), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][1]  (.Q(\ram[251][1] ), 
	.D(n4599), 
	.CK(clk));
   DFFHQX1 \ram_reg[251][0]  (.Q(\ram[251][0] ), 
	.D(n4598), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][15]  (.Q(\ram[247][15] ), 
	.D(n4549), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][14]  (.Q(\ram[247][14] ), 
	.D(n4548), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][13]  (.Q(\ram[247][13] ), 
	.D(n4547), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][12]  (.Q(\ram[247][12] ), 
	.D(n4546), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][11]  (.Q(\ram[247][11] ), 
	.D(n4545), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][10]  (.Q(\ram[247][10] ), 
	.D(n4544), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][9]  (.Q(\ram[247][9] ), 
	.D(n4543), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][8]  (.Q(\ram[247][8] ), 
	.D(n4542), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][7]  (.Q(\ram[247][7] ), 
	.D(n4541), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][6]  (.Q(\ram[247][6] ), 
	.D(n4540), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][5]  (.Q(\ram[247][5] ), 
	.D(n4539), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][4]  (.Q(\ram[247][4] ), 
	.D(n4538), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][3]  (.Q(\ram[247][3] ), 
	.D(n4537), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][2]  (.Q(\ram[247][2] ), 
	.D(n4536), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][1]  (.Q(\ram[247][1] ), 
	.D(n4535), 
	.CK(clk));
   DFFHQX1 \ram_reg[247][0]  (.Q(\ram[247][0] ), 
	.D(n4534), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][15]  (.Q(\ram[243][15] ), 
	.D(n4485), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][14]  (.Q(\ram[243][14] ), 
	.D(n4484), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][13]  (.Q(\ram[243][13] ), 
	.D(n4483), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][12]  (.Q(\ram[243][12] ), 
	.D(n4482), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][11]  (.Q(\ram[243][11] ), 
	.D(n4481), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][10]  (.Q(\ram[243][10] ), 
	.D(n4480), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][9]  (.Q(\ram[243][9] ), 
	.D(n4479), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][8]  (.Q(\ram[243][8] ), 
	.D(n4478), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][7]  (.Q(\ram[243][7] ), 
	.D(n4477), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][6]  (.Q(\ram[243][6] ), 
	.D(n4476), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][5]  (.Q(\ram[243][5] ), 
	.D(n4475), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][4]  (.Q(\ram[243][4] ), 
	.D(n4474), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][3]  (.Q(\ram[243][3] ), 
	.D(n4473), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][2]  (.Q(\ram[243][2] ), 
	.D(n4472), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][1]  (.Q(\ram[243][1] ), 
	.D(n4471), 
	.CK(clk));
   DFFHQX1 \ram_reg[243][0]  (.Q(\ram[243][0] ), 
	.D(n4470), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][15]  (.Q(\ram[239][15] ), 
	.D(n4421), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][14]  (.Q(\ram[239][14] ), 
	.D(n4420), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][13]  (.Q(\ram[239][13] ), 
	.D(n4419), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][12]  (.Q(\ram[239][12] ), 
	.D(n4418), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][11]  (.Q(\ram[239][11] ), 
	.D(n4417), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][10]  (.Q(\ram[239][10] ), 
	.D(n4416), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][9]  (.Q(\ram[239][9] ), 
	.D(n4415), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][8]  (.Q(\ram[239][8] ), 
	.D(n4414), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][7]  (.Q(\ram[239][7] ), 
	.D(n4413), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][6]  (.Q(\ram[239][6] ), 
	.D(n4412), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][5]  (.Q(\ram[239][5] ), 
	.D(n4411), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][4]  (.Q(\ram[239][4] ), 
	.D(n4410), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][3]  (.Q(\ram[239][3] ), 
	.D(n4409), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][2]  (.Q(\ram[239][2] ), 
	.D(n4408), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][1]  (.Q(\ram[239][1] ), 
	.D(n4407), 
	.CK(clk));
   DFFHQX1 \ram_reg[239][0]  (.Q(\ram[239][0] ), 
	.D(n4406), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][15]  (.Q(\ram[235][15] ), 
	.D(n4357), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][14]  (.Q(\ram[235][14] ), 
	.D(n4356), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][13]  (.Q(\ram[235][13] ), 
	.D(n4355), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][12]  (.Q(\ram[235][12] ), 
	.D(n4354), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][11]  (.Q(\ram[235][11] ), 
	.D(n4353), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][10]  (.Q(\ram[235][10] ), 
	.D(n4352), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][9]  (.Q(\ram[235][9] ), 
	.D(n4351), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][8]  (.Q(\ram[235][8] ), 
	.D(n4350), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][7]  (.Q(\ram[235][7] ), 
	.D(n4349), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][6]  (.Q(\ram[235][6] ), 
	.D(n4348), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][5]  (.Q(\ram[235][5] ), 
	.D(n4347), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][4]  (.Q(\ram[235][4] ), 
	.D(n4346), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][3]  (.Q(\ram[235][3] ), 
	.D(n4345), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][2]  (.Q(\ram[235][2] ), 
	.D(n4344), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][1]  (.Q(\ram[235][1] ), 
	.D(n4343), 
	.CK(clk));
   DFFHQX1 \ram_reg[235][0]  (.Q(\ram[235][0] ), 
	.D(n4342), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][15]  (.Q(\ram[231][15] ), 
	.D(n4293), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][14]  (.Q(\ram[231][14] ), 
	.D(n4292), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][13]  (.Q(\ram[231][13] ), 
	.D(n4291), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][12]  (.Q(\ram[231][12] ), 
	.D(n4290), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][11]  (.Q(\ram[231][11] ), 
	.D(n4289), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][10]  (.Q(\ram[231][10] ), 
	.D(n4288), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][9]  (.Q(\ram[231][9] ), 
	.D(n4287), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][8]  (.Q(\ram[231][8] ), 
	.D(n4286), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][7]  (.Q(\ram[231][7] ), 
	.D(n4285), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][6]  (.Q(\ram[231][6] ), 
	.D(n4284), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][5]  (.Q(\ram[231][5] ), 
	.D(n4283), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][4]  (.Q(\ram[231][4] ), 
	.D(n4282), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][3]  (.Q(\ram[231][3] ), 
	.D(n4281), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][2]  (.Q(\ram[231][2] ), 
	.D(n4280), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][1]  (.Q(\ram[231][1] ), 
	.D(n4279), 
	.CK(clk));
   DFFHQX1 \ram_reg[231][0]  (.Q(\ram[231][0] ), 
	.D(n4278), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][15]  (.Q(\ram[227][15] ), 
	.D(n4229), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][14]  (.Q(\ram[227][14] ), 
	.D(n4228), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][13]  (.Q(\ram[227][13] ), 
	.D(n4227), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][12]  (.Q(\ram[227][12] ), 
	.D(n4226), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][11]  (.Q(\ram[227][11] ), 
	.D(n4225), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][10]  (.Q(\ram[227][10] ), 
	.D(n4224), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][9]  (.Q(\ram[227][9] ), 
	.D(n4223), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][8]  (.Q(\ram[227][8] ), 
	.D(n4222), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][7]  (.Q(\ram[227][7] ), 
	.D(n4221), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][6]  (.Q(\ram[227][6] ), 
	.D(n4220), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][5]  (.Q(\ram[227][5] ), 
	.D(n4219), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][4]  (.Q(\ram[227][4] ), 
	.D(n4218), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][3]  (.Q(\ram[227][3] ), 
	.D(n4217), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][2]  (.Q(\ram[227][2] ), 
	.D(n4216), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][1]  (.Q(\ram[227][1] ), 
	.D(n4215), 
	.CK(clk));
   DFFHQX1 \ram_reg[227][0]  (.Q(\ram[227][0] ), 
	.D(n4214), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][15]  (.Q(\ram[223][15] ), 
	.D(n4165), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][14]  (.Q(\ram[223][14] ), 
	.D(n4164), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][13]  (.Q(\ram[223][13] ), 
	.D(n4163), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][12]  (.Q(\ram[223][12] ), 
	.D(n4162), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][11]  (.Q(\ram[223][11] ), 
	.D(n4161), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][10]  (.Q(\ram[223][10] ), 
	.D(n4160), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][9]  (.Q(\ram[223][9] ), 
	.D(n4159), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][8]  (.Q(\ram[223][8] ), 
	.D(n4158), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][7]  (.Q(\ram[223][7] ), 
	.D(n4157), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][6]  (.Q(\ram[223][6] ), 
	.D(n4156), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][5]  (.Q(\ram[223][5] ), 
	.D(n4155), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][4]  (.Q(\ram[223][4] ), 
	.D(n4154), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][3]  (.Q(\ram[223][3] ), 
	.D(n4153), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][2]  (.Q(\ram[223][2] ), 
	.D(n4152), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][1]  (.Q(\ram[223][1] ), 
	.D(n4151), 
	.CK(clk));
   DFFHQX1 \ram_reg[223][0]  (.Q(\ram[223][0] ), 
	.D(n4150), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][15]  (.Q(\ram[219][15] ), 
	.D(n4101), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][14]  (.Q(\ram[219][14] ), 
	.D(n4100), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][13]  (.Q(\ram[219][13] ), 
	.D(n4099), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][12]  (.Q(\ram[219][12] ), 
	.D(n4098), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][11]  (.Q(\ram[219][11] ), 
	.D(n4097), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][10]  (.Q(\ram[219][10] ), 
	.D(n4096), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][9]  (.Q(\ram[219][9] ), 
	.D(n4095), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][8]  (.Q(\ram[219][8] ), 
	.D(n4094), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][7]  (.Q(\ram[219][7] ), 
	.D(n4093), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][6]  (.Q(\ram[219][6] ), 
	.D(n4092), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][5]  (.Q(\ram[219][5] ), 
	.D(n4091), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][4]  (.Q(\ram[219][4] ), 
	.D(n4090), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][3]  (.Q(\ram[219][3] ), 
	.D(n4089), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][2]  (.Q(\ram[219][2] ), 
	.D(n4088), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][1]  (.Q(\ram[219][1] ), 
	.D(n4087), 
	.CK(clk));
   DFFHQX1 \ram_reg[219][0]  (.Q(\ram[219][0] ), 
	.D(n4086), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][15]  (.Q(\ram[215][15] ), 
	.D(n4037), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][14]  (.Q(\ram[215][14] ), 
	.D(n4036), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][13]  (.Q(\ram[215][13] ), 
	.D(n4035), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][12]  (.Q(\ram[215][12] ), 
	.D(n4034), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][11]  (.Q(\ram[215][11] ), 
	.D(n4033), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][10]  (.Q(\ram[215][10] ), 
	.D(n4032), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][9]  (.Q(\ram[215][9] ), 
	.D(n4031), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][8]  (.Q(\ram[215][8] ), 
	.D(n4030), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][7]  (.Q(\ram[215][7] ), 
	.D(n4029), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][6]  (.Q(\ram[215][6] ), 
	.D(n4028), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][5]  (.Q(\ram[215][5] ), 
	.D(n4027), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][4]  (.Q(\ram[215][4] ), 
	.D(n4026), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][3]  (.Q(\ram[215][3] ), 
	.D(n4025), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][2]  (.Q(\ram[215][2] ), 
	.D(n4024), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][1]  (.Q(\ram[215][1] ), 
	.D(n4023), 
	.CK(clk));
   DFFHQX1 \ram_reg[215][0]  (.Q(\ram[215][0] ), 
	.D(n4022), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][15]  (.Q(\ram[211][15] ), 
	.D(n3973), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][14]  (.Q(\ram[211][14] ), 
	.D(n3972), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][13]  (.Q(\ram[211][13] ), 
	.D(n3971), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][12]  (.Q(\ram[211][12] ), 
	.D(n3970), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][11]  (.Q(\ram[211][11] ), 
	.D(n3969), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][10]  (.Q(\ram[211][10] ), 
	.D(n3968), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][9]  (.Q(\ram[211][9] ), 
	.D(n3967), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][8]  (.Q(\ram[211][8] ), 
	.D(n3966), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][7]  (.Q(\ram[211][7] ), 
	.D(n3965), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][6]  (.Q(\ram[211][6] ), 
	.D(n3964), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][5]  (.Q(\ram[211][5] ), 
	.D(n3963), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][4]  (.Q(\ram[211][4] ), 
	.D(n3962), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][3]  (.Q(\ram[211][3] ), 
	.D(n3961), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][2]  (.Q(\ram[211][2] ), 
	.D(n3960), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][1]  (.Q(\ram[211][1] ), 
	.D(n3959), 
	.CK(clk));
   DFFHQX1 \ram_reg[211][0]  (.Q(\ram[211][0] ), 
	.D(n3958), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][15]  (.Q(\ram[207][15] ), 
	.D(n3909), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][14]  (.Q(\ram[207][14] ), 
	.D(n3908), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][13]  (.Q(\ram[207][13] ), 
	.D(n3907), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][12]  (.Q(\ram[207][12] ), 
	.D(n3906), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][11]  (.Q(\ram[207][11] ), 
	.D(n3905), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][10]  (.Q(\ram[207][10] ), 
	.D(n3904), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][9]  (.Q(\ram[207][9] ), 
	.D(n3903), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][8]  (.Q(\ram[207][8] ), 
	.D(n3902), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][7]  (.Q(\ram[207][7] ), 
	.D(n3901), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][6]  (.Q(\ram[207][6] ), 
	.D(n3900), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][5]  (.Q(\ram[207][5] ), 
	.D(n3899), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][4]  (.Q(\ram[207][4] ), 
	.D(n3898), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][3]  (.Q(\ram[207][3] ), 
	.D(n3897), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][2]  (.Q(\ram[207][2] ), 
	.D(n3896), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][1]  (.Q(\ram[207][1] ), 
	.D(n3895), 
	.CK(clk));
   DFFHQX1 \ram_reg[207][0]  (.Q(\ram[207][0] ), 
	.D(n3894), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][15]  (.Q(\ram[203][15] ), 
	.D(n3845), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][14]  (.Q(\ram[203][14] ), 
	.D(n3844), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][13]  (.Q(\ram[203][13] ), 
	.D(n3843), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][12]  (.Q(\ram[203][12] ), 
	.D(n3842), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][11]  (.Q(\ram[203][11] ), 
	.D(n3841), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][10]  (.Q(\ram[203][10] ), 
	.D(n3840), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][9]  (.Q(\ram[203][9] ), 
	.D(n3839), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][8]  (.Q(\ram[203][8] ), 
	.D(n3838), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][7]  (.Q(\ram[203][7] ), 
	.D(n3837), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][6]  (.Q(\ram[203][6] ), 
	.D(n3836), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][5]  (.Q(\ram[203][5] ), 
	.D(n3835), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][4]  (.Q(\ram[203][4] ), 
	.D(n3834), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][3]  (.Q(\ram[203][3] ), 
	.D(n3833), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][2]  (.Q(\ram[203][2] ), 
	.D(n3832), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][1]  (.Q(\ram[203][1] ), 
	.D(n3831), 
	.CK(clk));
   DFFHQX1 \ram_reg[203][0]  (.Q(\ram[203][0] ), 
	.D(n3830), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][15]  (.Q(\ram[199][15] ), 
	.D(n3781), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][14]  (.Q(\ram[199][14] ), 
	.D(n3780), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][13]  (.Q(\ram[199][13] ), 
	.D(n3779), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][12]  (.Q(\ram[199][12] ), 
	.D(n3778), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][11]  (.Q(\ram[199][11] ), 
	.D(n3777), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][10]  (.Q(\ram[199][10] ), 
	.D(n3776), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][9]  (.Q(\ram[199][9] ), 
	.D(n3775), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][8]  (.Q(\ram[199][8] ), 
	.D(n3774), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][7]  (.Q(\ram[199][7] ), 
	.D(n3773), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][6]  (.Q(\ram[199][6] ), 
	.D(n3772), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][5]  (.Q(\ram[199][5] ), 
	.D(n3771), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][4]  (.Q(\ram[199][4] ), 
	.D(n3770), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][3]  (.Q(\ram[199][3] ), 
	.D(n3769), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][2]  (.Q(\ram[199][2] ), 
	.D(n3768), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][1]  (.Q(\ram[199][1] ), 
	.D(n3767), 
	.CK(clk));
   DFFHQX1 \ram_reg[199][0]  (.Q(\ram[199][0] ), 
	.D(n3766), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][15]  (.Q(\ram[195][15] ), 
	.D(n3717), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][14]  (.Q(\ram[195][14] ), 
	.D(n3716), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][13]  (.Q(\ram[195][13] ), 
	.D(n3715), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][12]  (.Q(\ram[195][12] ), 
	.D(n3714), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][11]  (.Q(\ram[195][11] ), 
	.D(n3713), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][10]  (.Q(\ram[195][10] ), 
	.D(n3712), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][9]  (.Q(\ram[195][9] ), 
	.D(n3711), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][8]  (.Q(\ram[195][8] ), 
	.D(n3710), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][7]  (.Q(\ram[195][7] ), 
	.D(n3709), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][6]  (.Q(\ram[195][6] ), 
	.D(n3708), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][5]  (.Q(\ram[195][5] ), 
	.D(n3707), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][4]  (.Q(\ram[195][4] ), 
	.D(n3706), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][3]  (.Q(\ram[195][3] ), 
	.D(n3705), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][2]  (.Q(\ram[195][2] ), 
	.D(n3704), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][1]  (.Q(\ram[195][1] ), 
	.D(n3703), 
	.CK(clk));
   DFFHQX1 \ram_reg[195][0]  (.Q(\ram[195][0] ), 
	.D(n3702), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][15]  (.Q(\ram[191][15] ), 
	.D(n3653), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][14]  (.Q(\ram[191][14] ), 
	.D(n3652), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][13]  (.Q(\ram[191][13] ), 
	.D(n3651), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][12]  (.Q(\ram[191][12] ), 
	.D(n3650), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][11]  (.Q(\ram[191][11] ), 
	.D(n3649), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][10]  (.Q(\ram[191][10] ), 
	.D(n3648), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][9]  (.Q(\ram[191][9] ), 
	.D(n3647), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][8]  (.Q(\ram[191][8] ), 
	.D(n3646), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][7]  (.Q(\ram[191][7] ), 
	.D(n3645), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][6]  (.Q(\ram[191][6] ), 
	.D(n3644), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][5]  (.Q(\ram[191][5] ), 
	.D(n3643), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][4]  (.Q(\ram[191][4] ), 
	.D(n3642), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][3]  (.Q(\ram[191][3] ), 
	.D(n3641), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][2]  (.Q(\ram[191][2] ), 
	.D(n3640), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][1]  (.Q(\ram[191][1] ), 
	.D(n3639), 
	.CK(clk));
   DFFHQX1 \ram_reg[191][0]  (.Q(\ram[191][0] ), 
	.D(n3638), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][15]  (.Q(\ram[187][15] ), 
	.D(n3589), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][14]  (.Q(\ram[187][14] ), 
	.D(n3588), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][13]  (.Q(\ram[187][13] ), 
	.D(n3587), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][12]  (.Q(\ram[187][12] ), 
	.D(n3586), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][11]  (.Q(\ram[187][11] ), 
	.D(n3585), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][10]  (.Q(\ram[187][10] ), 
	.D(n3584), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][9]  (.Q(\ram[187][9] ), 
	.D(n3583), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][8]  (.Q(\ram[187][8] ), 
	.D(n3582), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][7]  (.Q(\ram[187][7] ), 
	.D(n3581), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][6]  (.Q(\ram[187][6] ), 
	.D(n3580), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][5]  (.Q(\ram[187][5] ), 
	.D(n3579), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][4]  (.Q(\ram[187][4] ), 
	.D(n3578), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][3]  (.Q(\ram[187][3] ), 
	.D(n3577), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][2]  (.Q(\ram[187][2] ), 
	.D(n3576), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][1]  (.Q(\ram[187][1] ), 
	.D(n3575), 
	.CK(clk));
   DFFHQX1 \ram_reg[187][0]  (.Q(\ram[187][0] ), 
	.D(n3574), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][15]  (.Q(\ram[183][15] ), 
	.D(n3525), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][14]  (.Q(\ram[183][14] ), 
	.D(n3524), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][13]  (.Q(\ram[183][13] ), 
	.D(n3523), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][12]  (.Q(\ram[183][12] ), 
	.D(n3522), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][11]  (.Q(\ram[183][11] ), 
	.D(n3521), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][10]  (.Q(\ram[183][10] ), 
	.D(n3520), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][9]  (.Q(\ram[183][9] ), 
	.D(n3519), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][8]  (.Q(\ram[183][8] ), 
	.D(n3518), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][7]  (.Q(\ram[183][7] ), 
	.D(n3517), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][6]  (.Q(\ram[183][6] ), 
	.D(n3516), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][5]  (.Q(\ram[183][5] ), 
	.D(n3515), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][4]  (.Q(\ram[183][4] ), 
	.D(n3514), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][3]  (.Q(\ram[183][3] ), 
	.D(n3513), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][2]  (.Q(\ram[183][2] ), 
	.D(n3512), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][1]  (.Q(\ram[183][1] ), 
	.D(n3511), 
	.CK(clk));
   DFFHQX1 \ram_reg[183][0]  (.Q(\ram[183][0] ), 
	.D(n3510), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][15]  (.Q(\ram[179][15] ), 
	.D(n3461), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][14]  (.Q(\ram[179][14] ), 
	.D(n3460), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][13]  (.Q(\ram[179][13] ), 
	.D(n3459), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][12]  (.Q(\ram[179][12] ), 
	.D(n3458), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][11]  (.Q(\ram[179][11] ), 
	.D(n3457), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][10]  (.Q(\ram[179][10] ), 
	.D(n3456), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][9]  (.Q(\ram[179][9] ), 
	.D(n3455), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][8]  (.Q(\ram[179][8] ), 
	.D(n3454), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][7]  (.Q(\ram[179][7] ), 
	.D(n3453), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][6]  (.Q(\ram[179][6] ), 
	.D(n3452), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][5]  (.Q(\ram[179][5] ), 
	.D(n3451), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][4]  (.Q(\ram[179][4] ), 
	.D(n3450), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][3]  (.Q(\ram[179][3] ), 
	.D(n3449), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][2]  (.Q(\ram[179][2] ), 
	.D(n3448), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][1]  (.Q(\ram[179][1] ), 
	.D(n3447), 
	.CK(clk));
   DFFHQX1 \ram_reg[179][0]  (.Q(\ram[179][0] ), 
	.D(n3446), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][15]  (.Q(\ram[175][15] ), 
	.D(n3397), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][14]  (.Q(\ram[175][14] ), 
	.D(n3396), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][13]  (.Q(\ram[175][13] ), 
	.D(n3395), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][12]  (.Q(\ram[175][12] ), 
	.D(n3394), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][11]  (.Q(\ram[175][11] ), 
	.D(n3393), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][10]  (.Q(\ram[175][10] ), 
	.D(n3392), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][9]  (.Q(\ram[175][9] ), 
	.D(n3391), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][8]  (.Q(\ram[175][8] ), 
	.D(n3390), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][7]  (.Q(\ram[175][7] ), 
	.D(n3389), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][6]  (.Q(\ram[175][6] ), 
	.D(n3388), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][5]  (.Q(\ram[175][5] ), 
	.D(n3387), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][4]  (.Q(\ram[175][4] ), 
	.D(n3386), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][3]  (.Q(\ram[175][3] ), 
	.D(n3385), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][2]  (.Q(\ram[175][2] ), 
	.D(n3384), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][1]  (.Q(\ram[175][1] ), 
	.D(n3383), 
	.CK(clk));
   DFFHQX1 \ram_reg[175][0]  (.Q(\ram[175][0] ), 
	.D(n3382), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][15]  (.Q(\ram[171][15] ), 
	.D(n3333), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][14]  (.Q(\ram[171][14] ), 
	.D(n3332), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][13]  (.Q(\ram[171][13] ), 
	.D(n3331), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][12]  (.Q(\ram[171][12] ), 
	.D(n3330), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][11]  (.Q(\ram[171][11] ), 
	.D(n3329), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][10]  (.Q(\ram[171][10] ), 
	.D(n3328), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][9]  (.Q(\ram[171][9] ), 
	.D(n3327), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][8]  (.Q(\ram[171][8] ), 
	.D(n3326), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][7]  (.Q(\ram[171][7] ), 
	.D(n3325), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][6]  (.Q(\ram[171][6] ), 
	.D(n3324), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][5]  (.Q(\ram[171][5] ), 
	.D(n3323), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][4]  (.Q(\ram[171][4] ), 
	.D(n3322), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][3]  (.Q(\ram[171][3] ), 
	.D(n3321), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][2]  (.Q(\ram[171][2] ), 
	.D(n3320), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][1]  (.Q(\ram[171][1] ), 
	.D(n3319), 
	.CK(clk));
   DFFHQX1 \ram_reg[171][0]  (.Q(\ram[171][0] ), 
	.D(n3318), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][15]  (.Q(\ram[167][15] ), 
	.D(n3269), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][14]  (.Q(\ram[167][14] ), 
	.D(n3268), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][13]  (.Q(\ram[167][13] ), 
	.D(n3267), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][12]  (.Q(\ram[167][12] ), 
	.D(n3266), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][11]  (.Q(\ram[167][11] ), 
	.D(n3265), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][10]  (.Q(\ram[167][10] ), 
	.D(n3264), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][9]  (.Q(\ram[167][9] ), 
	.D(n3263), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][8]  (.Q(\ram[167][8] ), 
	.D(n3262), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][7]  (.Q(\ram[167][7] ), 
	.D(n3261), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][6]  (.Q(\ram[167][6] ), 
	.D(n3260), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][5]  (.Q(\ram[167][5] ), 
	.D(n3259), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][4]  (.Q(\ram[167][4] ), 
	.D(n3258), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][3]  (.Q(\ram[167][3] ), 
	.D(n3257), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][2]  (.Q(\ram[167][2] ), 
	.D(n3256), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][1]  (.Q(\ram[167][1] ), 
	.D(n3255), 
	.CK(clk));
   DFFHQX1 \ram_reg[167][0]  (.Q(\ram[167][0] ), 
	.D(n3254), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][15]  (.Q(\ram[163][15] ), 
	.D(n3205), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][14]  (.Q(\ram[163][14] ), 
	.D(n3204), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][13]  (.Q(\ram[163][13] ), 
	.D(n3203), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][12]  (.Q(\ram[163][12] ), 
	.D(n3202), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][11]  (.Q(\ram[163][11] ), 
	.D(n3201), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][10]  (.Q(\ram[163][10] ), 
	.D(n3200), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][9]  (.Q(\ram[163][9] ), 
	.D(n3199), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][8]  (.Q(\ram[163][8] ), 
	.D(n3198), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][7]  (.Q(\ram[163][7] ), 
	.D(n3197), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][6]  (.Q(\ram[163][6] ), 
	.D(n3196), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][5]  (.Q(\ram[163][5] ), 
	.D(n3195), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][4]  (.Q(\ram[163][4] ), 
	.D(n3194), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][3]  (.Q(\ram[163][3] ), 
	.D(n3193), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][2]  (.Q(\ram[163][2] ), 
	.D(n3192), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][1]  (.Q(\ram[163][1] ), 
	.D(n3191), 
	.CK(clk));
   DFFHQX1 \ram_reg[163][0]  (.Q(\ram[163][0] ), 
	.D(n3190), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][15]  (.Q(\ram[159][15] ), 
	.D(n3141), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][14]  (.Q(\ram[159][14] ), 
	.D(n3140), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][13]  (.Q(\ram[159][13] ), 
	.D(n3139), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][12]  (.Q(\ram[159][12] ), 
	.D(n3138), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][11]  (.Q(\ram[159][11] ), 
	.D(n3137), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][10]  (.Q(\ram[159][10] ), 
	.D(n3136), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][9]  (.Q(\ram[159][9] ), 
	.D(n3135), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][8]  (.Q(\ram[159][8] ), 
	.D(n3134), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][7]  (.Q(\ram[159][7] ), 
	.D(n3133), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][6]  (.Q(\ram[159][6] ), 
	.D(n3132), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][5]  (.Q(\ram[159][5] ), 
	.D(n3131), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][4]  (.Q(\ram[159][4] ), 
	.D(n3130), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][3]  (.Q(\ram[159][3] ), 
	.D(n3129), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][2]  (.Q(\ram[159][2] ), 
	.D(n3128), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][1]  (.Q(\ram[159][1] ), 
	.D(n3127), 
	.CK(clk));
   DFFHQX1 \ram_reg[159][0]  (.Q(\ram[159][0] ), 
	.D(n3126), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][15]  (.Q(\ram[155][15] ), 
	.D(n3077), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][14]  (.Q(\ram[155][14] ), 
	.D(n3076), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][13]  (.Q(\ram[155][13] ), 
	.D(n3075), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][12]  (.Q(\ram[155][12] ), 
	.D(n3074), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][11]  (.Q(\ram[155][11] ), 
	.D(n3073), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][10]  (.Q(\ram[155][10] ), 
	.D(n3072), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][9]  (.Q(\ram[155][9] ), 
	.D(n3071), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][8]  (.Q(\ram[155][8] ), 
	.D(n3070), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][7]  (.Q(\ram[155][7] ), 
	.D(n3069), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][6]  (.Q(\ram[155][6] ), 
	.D(n3068), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][5]  (.Q(\ram[155][5] ), 
	.D(n3067), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][4]  (.Q(\ram[155][4] ), 
	.D(n3066), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][3]  (.Q(\ram[155][3] ), 
	.D(n3065), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][2]  (.Q(\ram[155][2] ), 
	.D(n3064), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][1]  (.Q(\ram[155][1] ), 
	.D(n3063), 
	.CK(clk));
   DFFHQX1 \ram_reg[155][0]  (.Q(\ram[155][0] ), 
	.D(n3062), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][15]  (.Q(\ram[151][15] ), 
	.D(n3013), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][14]  (.Q(\ram[151][14] ), 
	.D(n3012), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][13]  (.Q(\ram[151][13] ), 
	.D(n3011), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][12]  (.Q(\ram[151][12] ), 
	.D(n3010), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][11]  (.Q(\ram[151][11] ), 
	.D(n3009), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][10]  (.Q(\ram[151][10] ), 
	.D(n3008), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][9]  (.Q(\ram[151][9] ), 
	.D(n3007), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][8]  (.Q(\ram[151][8] ), 
	.D(n3006), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][7]  (.Q(\ram[151][7] ), 
	.D(n3005), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][6]  (.Q(\ram[151][6] ), 
	.D(n3004), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][5]  (.Q(\ram[151][5] ), 
	.D(n3003), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][4]  (.Q(\ram[151][4] ), 
	.D(n3002), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][3]  (.Q(\ram[151][3] ), 
	.D(n3001), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][2]  (.Q(\ram[151][2] ), 
	.D(n3000), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][1]  (.Q(\ram[151][1] ), 
	.D(n2999), 
	.CK(clk));
   DFFHQX1 \ram_reg[151][0]  (.Q(\ram[151][0] ), 
	.D(n2998), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][15]  (.Q(\ram[147][15] ), 
	.D(n2949), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][14]  (.Q(\ram[147][14] ), 
	.D(n2948), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][13]  (.Q(\ram[147][13] ), 
	.D(n2947), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][12]  (.Q(\ram[147][12] ), 
	.D(n2946), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][11]  (.Q(\ram[147][11] ), 
	.D(n2945), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][10]  (.Q(\ram[147][10] ), 
	.D(n2944), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][9]  (.Q(\ram[147][9] ), 
	.D(n2943), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][8]  (.Q(\ram[147][8] ), 
	.D(n2942), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][7]  (.Q(\ram[147][7] ), 
	.D(n2941), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][6]  (.Q(\ram[147][6] ), 
	.D(n2940), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][5]  (.Q(\ram[147][5] ), 
	.D(n2939), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][4]  (.Q(\ram[147][4] ), 
	.D(n2938), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][3]  (.Q(\ram[147][3] ), 
	.D(n2937), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][2]  (.Q(\ram[147][2] ), 
	.D(n2936), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][1]  (.Q(\ram[147][1] ), 
	.D(n2935), 
	.CK(clk));
   DFFHQX1 \ram_reg[147][0]  (.Q(\ram[147][0] ), 
	.D(n2934), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][15]  (.Q(\ram[143][15] ), 
	.D(n2885), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][14]  (.Q(\ram[143][14] ), 
	.D(n2884), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][13]  (.Q(\ram[143][13] ), 
	.D(n2883), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][12]  (.Q(\ram[143][12] ), 
	.D(n2882), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][11]  (.Q(\ram[143][11] ), 
	.D(n2881), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][10]  (.Q(\ram[143][10] ), 
	.D(n2880), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][9]  (.Q(\ram[143][9] ), 
	.D(n2879), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][8]  (.Q(\ram[143][8] ), 
	.D(n2878), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][7]  (.Q(\ram[143][7] ), 
	.D(n2877), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][6]  (.Q(\ram[143][6] ), 
	.D(n2876), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][5]  (.Q(\ram[143][5] ), 
	.D(n2875), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][4]  (.Q(\ram[143][4] ), 
	.D(n2874), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][3]  (.Q(\ram[143][3] ), 
	.D(n2873), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][2]  (.Q(\ram[143][2] ), 
	.D(n2872), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][1]  (.Q(\ram[143][1] ), 
	.D(n2871), 
	.CK(clk));
   DFFHQX1 \ram_reg[143][0]  (.Q(\ram[143][0] ), 
	.D(n2870), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][15]  (.Q(\ram[139][15] ), 
	.D(n2821), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][14]  (.Q(\ram[139][14] ), 
	.D(n2820), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][13]  (.Q(\ram[139][13] ), 
	.D(n2819), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][12]  (.Q(\ram[139][12] ), 
	.D(n2818), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][11]  (.Q(\ram[139][11] ), 
	.D(n2817), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][10]  (.Q(\ram[139][10] ), 
	.D(n2816), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][9]  (.Q(\ram[139][9] ), 
	.D(n2815), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][8]  (.Q(\ram[139][8] ), 
	.D(n2814), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][7]  (.Q(\ram[139][7] ), 
	.D(n2813), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][6]  (.Q(\ram[139][6] ), 
	.D(n2812), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][5]  (.Q(\ram[139][5] ), 
	.D(n2811), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][4]  (.Q(\ram[139][4] ), 
	.D(n2810), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][3]  (.Q(\ram[139][3] ), 
	.D(n2809), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][2]  (.Q(\ram[139][2] ), 
	.D(n2808), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][1]  (.Q(\ram[139][1] ), 
	.D(n2807), 
	.CK(clk));
   DFFHQX1 \ram_reg[139][0]  (.Q(\ram[139][0] ), 
	.D(n2806), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][15]  (.Q(\ram[135][15] ), 
	.D(n2757), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][14]  (.Q(\ram[135][14] ), 
	.D(n2756), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][13]  (.Q(\ram[135][13] ), 
	.D(n2755), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][12]  (.Q(\ram[135][12] ), 
	.D(n2754), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][11]  (.Q(\ram[135][11] ), 
	.D(n2753), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][10]  (.Q(\ram[135][10] ), 
	.D(n2752), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][9]  (.Q(\ram[135][9] ), 
	.D(n2751), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][8]  (.Q(\ram[135][8] ), 
	.D(n2750), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][7]  (.Q(\ram[135][7] ), 
	.D(n2749), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][6]  (.Q(\ram[135][6] ), 
	.D(n2748), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][5]  (.Q(\ram[135][5] ), 
	.D(n2747), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][4]  (.Q(\ram[135][4] ), 
	.D(n2746), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][3]  (.Q(\ram[135][3] ), 
	.D(n2745), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][2]  (.Q(\ram[135][2] ), 
	.D(n2744), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][1]  (.Q(\ram[135][1] ), 
	.D(n2743), 
	.CK(clk));
   DFFHQX1 \ram_reg[135][0]  (.Q(\ram[135][0] ), 
	.D(n2742), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][15]  (.Q(\ram[131][15] ), 
	.D(n2693), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][14]  (.Q(\ram[131][14] ), 
	.D(n2692), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][13]  (.Q(\ram[131][13] ), 
	.D(n2691), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][12]  (.Q(\ram[131][12] ), 
	.D(n2690), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][11]  (.Q(\ram[131][11] ), 
	.D(n2689), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][10]  (.Q(\ram[131][10] ), 
	.D(n2688), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][9]  (.Q(\ram[131][9] ), 
	.D(n2687), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][8]  (.Q(\ram[131][8] ), 
	.D(n2686), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][7]  (.Q(\ram[131][7] ), 
	.D(n2685), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][6]  (.Q(\ram[131][6] ), 
	.D(n2684), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][5]  (.Q(\ram[131][5] ), 
	.D(n2683), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][4]  (.Q(\ram[131][4] ), 
	.D(n2682), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][3]  (.Q(\ram[131][3] ), 
	.D(n2681), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][2]  (.Q(\ram[131][2] ), 
	.D(n2680), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][1]  (.Q(\ram[131][1] ), 
	.D(n2679), 
	.CK(clk));
   DFFHQX1 \ram_reg[131][0]  (.Q(\ram[131][0] ), 
	.D(n2678), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][15]  (.Q(\ram[127][15] ), 
	.D(n2629), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][14]  (.Q(\ram[127][14] ), 
	.D(n2628), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][13]  (.Q(\ram[127][13] ), 
	.D(n2627), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][12]  (.Q(\ram[127][12] ), 
	.D(n2626), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][11]  (.Q(\ram[127][11] ), 
	.D(n2625), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][10]  (.Q(\ram[127][10] ), 
	.D(n2624), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][9]  (.Q(\ram[127][9] ), 
	.D(n2623), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][8]  (.Q(\ram[127][8] ), 
	.D(n2622), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][7]  (.Q(\ram[127][7] ), 
	.D(n2621), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][6]  (.Q(\ram[127][6] ), 
	.D(n2620), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][5]  (.Q(\ram[127][5] ), 
	.D(n2619), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][4]  (.Q(\ram[127][4] ), 
	.D(n2618), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][3]  (.Q(\ram[127][3] ), 
	.D(n2617), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][2]  (.Q(\ram[127][2] ), 
	.D(n2616), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][1]  (.Q(\ram[127][1] ), 
	.D(n2615), 
	.CK(clk));
   DFFHQX1 \ram_reg[127][0]  (.Q(\ram[127][0] ), 
	.D(n2614), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][15]  (.Q(\ram[123][15] ), 
	.D(n2565), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][14]  (.Q(\ram[123][14] ), 
	.D(n2564), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][13]  (.Q(\ram[123][13] ), 
	.D(n2563), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][12]  (.Q(\ram[123][12] ), 
	.D(n2562), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][11]  (.Q(\ram[123][11] ), 
	.D(n2561), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][10]  (.Q(\ram[123][10] ), 
	.D(n2560), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][9]  (.Q(\ram[123][9] ), 
	.D(n2559), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][8]  (.Q(\ram[123][8] ), 
	.D(n2558), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][7]  (.Q(\ram[123][7] ), 
	.D(n2557), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][6]  (.Q(\ram[123][6] ), 
	.D(n2556), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][5]  (.Q(\ram[123][5] ), 
	.D(n2555), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][4]  (.Q(\ram[123][4] ), 
	.D(n2554), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][3]  (.Q(\ram[123][3] ), 
	.D(n2553), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][2]  (.Q(\ram[123][2] ), 
	.D(n2552), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][1]  (.Q(\ram[123][1] ), 
	.D(n2551), 
	.CK(clk));
   DFFHQX1 \ram_reg[123][0]  (.Q(\ram[123][0] ), 
	.D(n2550), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][15]  (.Q(\ram[119][15] ), 
	.D(n2501), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][14]  (.Q(\ram[119][14] ), 
	.D(n2500), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][13]  (.Q(\ram[119][13] ), 
	.D(n2499), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][12]  (.Q(\ram[119][12] ), 
	.D(n2498), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][11]  (.Q(\ram[119][11] ), 
	.D(n2497), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][10]  (.Q(\ram[119][10] ), 
	.D(n2496), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][9]  (.Q(\ram[119][9] ), 
	.D(n2495), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][8]  (.Q(\ram[119][8] ), 
	.D(n2494), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][7]  (.Q(\ram[119][7] ), 
	.D(n2493), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][6]  (.Q(\ram[119][6] ), 
	.D(n2492), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][5]  (.Q(\ram[119][5] ), 
	.D(n2491), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][4]  (.Q(\ram[119][4] ), 
	.D(n2490), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][3]  (.Q(\ram[119][3] ), 
	.D(n2489), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][2]  (.Q(\ram[119][2] ), 
	.D(n2488), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][1]  (.Q(\ram[119][1] ), 
	.D(n2487), 
	.CK(clk));
   DFFHQX1 \ram_reg[119][0]  (.Q(\ram[119][0] ), 
	.D(n2486), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][15]  (.Q(\ram[115][15] ), 
	.D(n2437), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][14]  (.Q(\ram[115][14] ), 
	.D(n2436), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][13]  (.Q(\ram[115][13] ), 
	.D(n2435), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][12]  (.Q(\ram[115][12] ), 
	.D(n2434), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][11]  (.Q(\ram[115][11] ), 
	.D(n2433), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][10]  (.Q(\ram[115][10] ), 
	.D(n2432), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][9]  (.Q(\ram[115][9] ), 
	.D(n2431), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][8]  (.Q(\ram[115][8] ), 
	.D(n2430), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][7]  (.Q(\ram[115][7] ), 
	.D(n2429), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][6]  (.Q(\ram[115][6] ), 
	.D(n2428), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][5]  (.Q(\ram[115][5] ), 
	.D(n2427), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][4]  (.Q(\ram[115][4] ), 
	.D(n2426), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][3]  (.Q(\ram[115][3] ), 
	.D(n2425), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][2]  (.Q(\ram[115][2] ), 
	.D(n2424), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][1]  (.Q(\ram[115][1] ), 
	.D(n2423), 
	.CK(clk));
   DFFHQX1 \ram_reg[115][0]  (.Q(\ram[115][0] ), 
	.D(n2422), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][15]  (.Q(\ram[111][15] ), 
	.D(n2373), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][14]  (.Q(\ram[111][14] ), 
	.D(n2372), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][13]  (.Q(\ram[111][13] ), 
	.D(n2371), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][12]  (.Q(\ram[111][12] ), 
	.D(n2370), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][11]  (.Q(\ram[111][11] ), 
	.D(n2369), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][10]  (.Q(\ram[111][10] ), 
	.D(n2368), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][9]  (.Q(\ram[111][9] ), 
	.D(n2367), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][8]  (.Q(\ram[111][8] ), 
	.D(n2366), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][7]  (.Q(\ram[111][7] ), 
	.D(n2365), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][6]  (.Q(\ram[111][6] ), 
	.D(n2364), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][5]  (.Q(\ram[111][5] ), 
	.D(n2363), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][4]  (.Q(\ram[111][4] ), 
	.D(n2362), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][3]  (.Q(\ram[111][3] ), 
	.D(n2361), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][2]  (.Q(\ram[111][2] ), 
	.D(n2360), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][1]  (.Q(\ram[111][1] ), 
	.D(n2359), 
	.CK(clk));
   DFFHQX1 \ram_reg[111][0]  (.Q(\ram[111][0] ), 
	.D(n2358), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][15]  (.Q(\ram[107][15] ), 
	.D(n2309), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][14]  (.Q(\ram[107][14] ), 
	.D(n2308), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][13]  (.Q(\ram[107][13] ), 
	.D(n2307), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][12]  (.Q(\ram[107][12] ), 
	.D(n2306), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][11]  (.Q(\ram[107][11] ), 
	.D(n2305), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][10]  (.Q(\ram[107][10] ), 
	.D(n2304), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][9]  (.Q(\ram[107][9] ), 
	.D(n2303), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][8]  (.Q(\ram[107][8] ), 
	.D(n2302), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][7]  (.Q(\ram[107][7] ), 
	.D(n2301), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][6]  (.Q(\ram[107][6] ), 
	.D(n2300), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][5]  (.Q(\ram[107][5] ), 
	.D(n2299), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][4]  (.Q(\ram[107][4] ), 
	.D(n2298), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][3]  (.Q(\ram[107][3] ), 
	.D(n2297), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][2]  (.Q(\ram[107][2] ), 
	.D(n2296), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][1]  (.Q(\ram[107][1] ), 
	.D(n2295), 
	.CK(clk));
   DFFHQX1 \ram_reg[107][0]  (.Q(\ram[107][0] ), 
	.D(n2294), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][15]  (.Q(\ram[103][15] ), 
	.D(n2245), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][14]  (.Q(\ram[103][14] ), 
	.D(n2244), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][13]  (.Q(\ram[103][13] ), 
	.D(n2243), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][12]  (.Q(\ram[103][12] ), 
	.D(n2242), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][11]  (.Q(\ram[103][11] ), 
	.D(n2241), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][10]  (.Q(\ram[103][10] ), 
	.D(n2240), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][9]  (.Q(\ram[103][9] ), 
	.D(n2239), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][8]  (.Q(\ram[103][8] ), 
	.D(n2238), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][7]  (.Q(\ram[103][7] ), 
	.D(n2237), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][6]  (.Q(\ram[103][6] ), 
	.D(n2236), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][5]  (.Q(\ram[103][5] ), 
	.D(n2235), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][4]  (.Q(\ram[103][4] ), 
	.D(n2234), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][3]  (.Q(\ram[103][3] ), 
	.D(n2233), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][2]  (.Q(\ram[103][2] ), 
	.D(n2232), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][1]  (.Q(\ram[103][1] ), 
	.D(n2231), 
	.CK(clk));
   DFFHQX1 \ram_reg[103][0]  (.Q(\ram[103][0] ), 
	.D(n2230), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][15]  (.Q(\ram[99][15] ), 
	.D(n2181), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][14]  (.Q(\ram[99][14] ), 
	.D(n2180), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][13]  (.Q(\ram[99][13] ), 
	.D(n2179), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][12]  (.Q(\ram[99][12] ), 
	.D(n2178), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][11]  (.Q(\ram[99][11] ), 
	.D(n2177), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][10]  (.Q(\ram[99][10] ), 
	.D(n2176), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][9]  (.Q(\ram[99][9] ), 
	.D(n2175), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][8]  (.Q(\ram[99][8] ), 
	.D(n2174), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][7]  (.Q(\ram[99][7] ), 
	.D(n2173), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][6]  (.Q(\ram[99][6] ), 
	.D(n2172), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][5]  (.Q(\ram[99][5] ), 
	.D(n2171), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][4]  (.Q(\ram[99][4] ), 
	.D(n2170), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][3]  (.Q(\ram[99][3] ), 
	.D(n2169), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][2]  (.Q(\ram[99][2] ), 
	.D(n2168), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][1]  (.Q(\ram[99][1] ), 
	.D(n2167), 
	.CK(clk));
   DFFHQX1 \ram_reg[99][0]  (.Q(\ram[99][0] ), 
	.D(n2166), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][15]  (.Q(\ram[95][15] ), 
	.D(n2117), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][14]  (.Q(\ram[95][14] ), 
	.D(n2116), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][13]  (.Q(\ram[95][13] ), 
	.D(n2115), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][12]  (.Q(\ram[95][12] ), 
	.D(n2114), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][11]  (.Q(\ram[95][11] ), 
	.D(n2113), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][10]  (.Q(\ram[95][10] ), 
	.D(n2112), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][9]  (.Q(\ram[95][9] ), 
	.D(n2111), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][8]  (.Q(\ram[95][8] ), 
	.D(n2110), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][7]  (.Q(\ram[95][7] ), 
	.D(n2109), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][6]  (.Q(\ram[95][6] ), 
	.D(n2108), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][5]  (.Q(\ram[95][5] ), 
	.D(n2107), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][4]  (.Q(\ram[95][4] ), 
	.D(n2106), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][3]  (.Q(\ram[95][3] ), 
	.D(n2105), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][2]  (.Q(\ram[95][2] ), 
	.D(n2104), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][1]  (.Q(\ram[95][1] ), 
	.D(n2103), 
	.CK(clk));
   DFFHQX1 \ram_reg[95][0]  (.Q(\ram[95][0] ), 
	.D(n2102), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][15]  (.Q(\ram[91][15] ), 
	.D(n2053), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][14]  (.Q(\ram[91][14] ), 
	.D(n2052), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][13]  (.Q(\ram[91][13] ), 
	.D(n2051), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][12]  (.Q(\ram[91][12] ), 
	.D(n2050), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][11]  (.Q(\ram[91][11] ), 
	.D(n2049), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][10]  (.Q(\ram[91][10] ), 
	.D(n2048), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][9]  (.Q(\ram[91][9] ), 
	.D(n2047), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][8]  (.Q(\ram[91][8] ), 
	.D(n2046), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][7]  (.Q(\ram[91][7] ), 
	.D(n2045), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][6]  (.Q(\ram[91][6] ), 
	.D(n2044), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][5]  (.Q(\ram[91][5] ), 
	.D(n2043), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][4]  (.Q(\ram[91][4] ), 
	.D(n2042), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][3]  (.Q(\ram[91][3] ), 
	.D(n2041), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][2]  (.Q(\ram[91][2] ), 
	.D(n2040), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][1]  (.Q(\ram[91][1] ), 
	.D(n2039), 
	.CK(clk));
   DFFHQX1 \ram_reg[91][0]  (.Q(\ram[91][0] ), 
	.D(n2038), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][15]  (.Q(\ram[87][15] ), 
	.D(n1989), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][14]  (.Q(\ram[87][14] ), 
	.D(n1988), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][13]  (.Q(\ram[87][13] ), 
	.D(n1987), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][12]  (.Q(\ram[87][12] ), 
	.D(n1986), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][11]  (.Q(\ram[87][11] ), 
	.D(n1985), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][10]  (.Q(\ram[87][10] ), 
	.D(n1984), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][9]  (.Q(\ram[87][9] ), 
	.D(n1983), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][8]  (.Q(\ram[87][8] ), 
	.D(n1982), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][7]  (.Q(\ram[87][7] ), 
	.D(n1981), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][6]  (.Q(\ram[87][6] ), 
	.D(n1980), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][5]  (.Q(\ram[87][5] ), 
	.D(n1979), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][4]  (.Q(\ram[87][4] ), 
	.D(n1978), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][3]  (.Q(\ram[87][3] ), 
	.D(n1977), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][2]  (.Q(\ram[87][2] ), 
	.D(n1976), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][1]  (.Q(\ram[87][1] ), 
	.D(n1975), 
	.CK(clk));
   DFFHQX1 \ram_reg[87][0]  (.Q(\ram[87][0] ), 
	.D(n1974), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][15]  (.Q(\ram[83][15] ), 
	.D(n1925), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][14]  (.Q(\ram[83][14] ), 
	.D(n1924), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][13]  (.Q(\ram[83][13] ), 
	.D(n1923), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][12]  (.Q(\ram[83][12] ), 
	.D(n1922), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][11]  (.Q(\ram[83][11] ), 
	.D(n1921), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][10]  (.Q(\ram[83][10] ), 
	.D(n1920), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][9]  (.Q(\ram[83][9] ), 
	.D(n1919), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][8]  (.Q(\ram[83][8] ), 
	.D(n1918), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][7]  (.Q(\ram[83][7] ), 
	.D(n1917), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][6]  (.Q(\ram[83][6] ), 
	.D(n1916), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][5]  (.Q(\ram[83][5] ), 
	.D(n1915), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][4]  (.Q(\ram[83][4] ), 
	.D(n1914), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][3]  (.Q(\ram[83][3] ), 
	.D(n1913), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][2]  (.Q(\ram[83][2] ), 
	.D(n1912), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][1]  (.Q(\ram[83][1] ), 
	.D(n1911), 
	.CK(clk));
   DFFHQX1 \ram_reg[83][0]  (.Q(\ram[83][0] ), 
	.D(n1910), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][15]  (.Q(\ram[79][15] ), 
	.D(n1861), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][14]  (.Q(\ram[79][14] ), 
	.D(n1860), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][13]  (.Q(\ram[79][13] ), 
	.D(n1859), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][12]  (.Q(\ram[79][12] ), 
	.D(n1858), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][11]  (.Q(\ram[79][11] ), 
	.D(n1857), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][10]  (.Q(\ram[79][10] ), 
	.D(n1856), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][9]  (.Q(\ram[79][9] ), 
	.D(n1855), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][8]  (.Q(\ram[79][8] ), 
	.D(n1854), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][7]  (.Q(\ram[79][7] ), 
	.D(n1853), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][6]  (.Q(\ram[79][6] ), 
	.D(n1852), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][5]  (.Q(\ram[79][5] ), 
	.D(n1851), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][4]  (.Q(\ram[79][4] ), 
	.D(n1850), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][3]  (.Q(\ram[79][3] ), 
	.D(n1849), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][2]  (.Q(\ram[79][2] ), 
	.D(n1848), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][1]  (.Q(\ram[79][1] ), 
	.D(n1847), 
	.CK(clk));
   DFFHQX1 \ram_reg[79][0]  (.Q(\ram[79][0] ), 
	.D(n1846), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][15]  (.Q(\ram[75][15] ), 
	.D(n1797), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][14]  (.Q(\ram[75][14] ), 
	.D(n1796), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][13]  (.Q(\ram[75][13] ), 
	.D(n1795), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][12]  (.Q(\ram[75][12] ), 
	.D(n1794), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][11]  (.Q(\ram[75][11] ), 
	.D(n1793), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][10]  (.Q(\ram[75][10] ), 
	.D(n1792), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][9]  (.Q(\ram[75][9] ), 
	.D(n1791), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][8]  (.Q(\ram[75][8] ), 
	.D(n1790), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][7]  (.Q(\ram[75][7] ), 
	.D(n1789), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][6]  (.Q(\ram[75][6] ), 
	.D(n1788), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][5]  (.Q(\ram[75][5] ), 
	.D(n1787), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][4]  (.Q(\ram[75][4] ), 
	.D(n1786), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][3]  (.Q(\ram[75][3] ), 
	.D(n1785), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][2]  (.Q(\ram[75][2] ), 
	.D(n1784), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][1]  (.Q(\ram[75][1] ), 
	.D(n1783), 
	.CK(clk));
   DFFHQX1 \ram_reg[75][0]  (.Q(\ram[75][0] ), 
	.D(n1782), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][15]  (.Q(\ram[71][15] ), 
	.D(n1733), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][14]  (.Q(\ram[71][14] ), 
	.D(n1732), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][13]  (.Q(\ram[71][13] ), 
	.D(n1731), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][12]  (.Q(\ram[71][12] ), 
	.D(n1730), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][11]  (.Q(\ram[71][11] ), 
	.D(n1729), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][10]  (.Q(\ram[71][10] ), 
	.D(n1728), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][9]  (.Q(\ram[71][9] ), 
	.D(n1727), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][8]  (.Q(\ram[71][8] ), 
	.D(n1726), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][7]  (.Q(\ram[71][7] ), 
	.D(n1725), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][6]  (.Q(\ram[71][6] ), 
	.D(n1724), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][5]  (.Q(\ram[71][5] ), 
	.D(n1723), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][4]  (.Q(\ram[71][4] ), 
	.D(n1722), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][3]  (.Q(\ram[71][3] ), 
	.D(n1721), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][2]  (.Q(\ram[71][2] ), 
	.D(n1720), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][1]  (.Q(\ram[71][1] ), 
	.D(n1719), 
	.CK(clk));
   DFFHQX1 \ram_reg[71][0]  (.Q(\ram[71][0] ), 
	.D(n1718), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][15]  (.Q(\ram[67][15] ), 
	.D(n1669), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][14]  (.Q(\ram[67][14] ), 
	.D(n1668), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][13]  (.Q(\ram[67][13] ), 
	.D(n1667), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][12]  (.Q(\ram[67][12] ), 
	.D(n1666), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][11]  (.Q(\ram[67][11] ), 
	.D(n1665), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][10]  (.Q(\ram[67][10] ), 
	.D(n1664), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][9]  (.Q(\ram[67][9] ), 
	.D(n1663), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][8]  (.Q(\ram[67][8] ), 
	.D(n1662), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][7]  (.Q(\ram[67][7] ), 
	.D(n1661), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][6]  (.Q(\ram[67][6] ), 
	.D(n1660), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][5]  (.Q(\ram[67][5] ), 
	.D(n1659), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][4]  (.Q(\ram[67][4] ), 
	.D(n1658), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][3]  (.Q(\ram[67][3] ), 
	.D(n1657), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][2]  (.Q(\ram[67][2] ), 
	.D(n1656), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][1]  (.Q(\ram[67][1] ), 
	.D(n1655), 
	.CK(clk));
   DFFHQX1 \ram_reg[67][0]  (.Q(\ram[67][0] ), 
	.D(n1654), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][15]  (.Q(\ram[63][15] ), 
	.D(n1605), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][14]  (.Q(\ram[63][14] ), 
	.D(n1604), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][13]  (.Q(\ram[63][13] ), 
	.D(n1603), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][12]  (.Q(\ram[63][12] ), 
	.D(n1602), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][11]  (.Q(\ram[63][11] ), 
	.D(n1601), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][10]  (.Q(\ram[63][10] ), 
	.D(n1600), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][9]  (.Q(\ram[63][9] ), 
	.D(n1599), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][8]  (.Q(\ram[63][8] ), 
	.D(n1598), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][7]  (.Q(\ram[63][7] ), 
	.D(n1597), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][6]  (.Q(\ram[63][6] ), 
	.D(n1596), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][5]  (.Q(\ram[63][5] ), 
	.D(n1595), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][4]  (.Q(\ram[63][4] ), 
	.D(n1594), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][3]  (.Q(\ram[63][3] ), 
	.D(n1593), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][2]  (.Q(\ram[63][2] ), 
	.D(n1592), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][1]  (.Q(\ram[63][1] ), 
	.D(n1591), 
	.CK(clk));
   DFFHQX1 \ram_reg[63][0]  (.Q(\ram[63][0] ), 
	.D(n1590), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][15]  (.Q(\ram[59][15] ), 
	.D(n1541), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][14]  (.Q(\ram[59][14] ), 
	.D(n1540), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][13]  (.Q(\ram[59][13] ), 
	.D(n1539), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][12]  (.Q(\ram[59][12] ), 
	.D(n1538), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][11]  (.Q(\ram[59][11] ), 
	.D(n1537), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][10]  (.Q(\ram[59][10] ), 
	.D(n1536), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][9]  (.Q(\ram[59][9] ), 
	.D(n1535), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][8]  (.Q(\ram[59][8] ), 
	.D(n1534), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][7]  (.Q(\ram[59][7] ), 
	.D(n1533), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][6]  (.Q(\ram[59][6] ), 
	.D(n1532), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][5]  (.Q(\ram[59][5] ), 
	.D(n1531), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][4]  (.Q(\ram[59][4] ), 
	.D(n1530), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][3]  (.Q(\ram[59][3] ), 
	.D(n1529), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][2]  (.Q(\ram[59][2] ), 
	.D(n1528), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][1]  (.Q(\ram[59][1] ), 
	.D(n1527), 
	.CK(clk));
   DFFHQX1 \ram_reg[59][0]  (.Q(\ram[59][0] ), 
	.D(n1526), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][15]  (.Q(\ram[55][15] ), 
	.D(n1477), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][14]  (.Q(\ram[55][14] ), 
	.D(n1476), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][13]  (.Q(\ram[55][13] ), 
	.D(n1475), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][12]  (.Q(\ram[55][12] ), 
	.D(n1474), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][11]  (.Q(\ram[55][11] ), 
	.D(n1473), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][10]  (.Q(\ram[55][10] ), 
	.D(n1472), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][9]  (.Q(\ram[55][9] ), 
	.D(n1471), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][8]  (.Q(\ram[55][8] ), 
	.D(n1470), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][7]  (.Q(\ram[55][7] ), 
	.D(n1469), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][6]  (.Q(\ram[55][6] ), 
	.D(n1468), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][5]  (.Q(\ram[55][5] ), 
	.D(n1467), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][4]  (.Q(\ram[55][4] ), 
	.D(n1466), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][3]  (.Q(\ram[55][3] ), 
	.D(n1465), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][2]  (.Q(\ram[55][2] ), 
	.D(n1464), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][1]  (.Q(\ram[55][1] ), 
	.D(n1463), 
	.CK(clk));
   DFFHQX1 \ram_reg[55][0]  (.Q(\ram[55][0] ), 
	.D(n1462), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][15]  (.Q(\ram[51][15] ), 
	.D(n1413), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][14]  (.Q(\ram[51][14] ), 
	.D(n1412), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][13]  (.Q(\ram[51][13] ), 
	.D(n1411), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][12]  (.Q(\ram[51][12] ), 
	.D(n1410), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][11]  (.Q(\ram[51][11] ), 
	.D(n1409), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][10]  (.Q(\ram[51][10] ), 
	.D(n1408), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][9]  (.Q(\ram[51][9] ), 
	.D(n1407), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][8]  (.Q(\ram[51][8] ), 
	.D(n1406), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][7]  (.Q(\ram[51][7] ), 
	.D(n1405), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][6]  (.Q(\ram[51][6] ), 
	.D(n1404), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][5]  (.Q(\ram[51][5] ), 
	.D(n1403), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][4]  (.Q(\ram[51][4] ), 
	.D(n1402), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][3]  (.Q(\ram[51][3] ), 
	.D(n1401), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][2]  (.Q(\ram[51][2] ), 
	.D(n1400), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][1]  (.Q(\ram[51][1] ), 
	.D(n1399), 
	.CK(clk));
   DFFHQX1 \ram_reg[51][0]  (.Q(\ram[51][0] ), 
	.D(n1398), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][15]  (.Q(\ram[47][15] ), 
	.D(n1349), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][14]  (.Q(\ram[47][14] ), 
	.D(n1348), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][13]  (.Q(\ram[47][13] ), 
	.D(n1347), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][12]  (.Q(\ram[47][12] ), 
	.D(n1346), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][11]  (.Q(\ram[47][11] ), 
	.D(n1345), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][10]  (.Q(\ram[47][10] ), 
	.D(n1344), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][9]  (.Q(\ram[47][9] ), 
	.D(n1343), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][8]  (.Q(\ram[47][8] ), 
	.D(n1342), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][7]  (.Q(\ram[47][7] ), 
	.D(n1341), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][6]  (.Q(\ram[47][6] ), 
	.D(n1340), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][5]  (.Q(\ram[47][5] ), 
	.D(n1339), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][4]  (.Q(\ram[47][4] ), 
	.D(n1338), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][3]  (.Q(\ram[47][3] ), 
	.D(n1337), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][2]  (.Q(\ram[47][2] ), 
	.D(n1336), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][1]  (.Q(\ram[47][1] ), 
	.D(n1335), 
	.CK(clk));
   DFFHQX1 \ram_reg[47][0]  (.Q(\ram[47][0] ), 
	.D(n1334), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][15]  (.Q(\ram[43][15] ), 
	.D(n1285), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][14]  (.Q(\ram[43][14] ), 
	.D(n1284), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][13]  (.Q(\ram[43][13] ), 
	.D(n1283), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][12]  (.Q(\ram[43][12] ), 
	.D(n1282), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][11]  (.Q(\ram[43][11] ), 
	.D(n1281), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][10]  (.Q(\ram[43][10] ), 
	.D(n1280), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][9]  (.Q(\ram[43][9] ), 
	.D(n1279), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][8]  (.Q(\ram[43][8] ), 
	.D(n1278), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][7]  (.Q(\ram[43][7] ), 
	.D(n1277), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][6]  (.Q(\ram[43][6] ), 
	.D(n1276), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][5]  (.Q(\ram[43][5] ), 
	.D(n1275), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][4]  (.Q(\ram[43][4] ), 
	.D(n1274), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][3]  (.Q(\ram[43][3] ), 
	.D(n1273), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][2]  (.Q(\ram[43][2] ), 
	.D(n1272), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][1]  (.Q(\ram[43][1] ), 
	.D(n1271), 
	.CK(clk));
   DFFHQX1 \ram_reg[43][0]  (.Q(\ram[43][0] ), 
	.D(n1270), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][15]  (.Q(\ram[39][15] ), 
	.D(n1221), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][14]  (.Q(\ram[39][14] ), 
	.D(n1220), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][13]  (.Q(\ram[39][13] ), 
	.D(n1219), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][12]  (.Q(\ram[39][12] ), 
	.D(n1218), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][11]  (.Q(\ram[39][11] ), 
	.D(n1217), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][10]  (.Q(\ram[39][10] ), 
	.D(n1216), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][9]  (.Q(\ram[39][9] ), 
	.D(n1215), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][8]  (.Q(\ram[39][8] ), 
	.D(n1214), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][7]  (.Q(\ram[39][7] ), 
	.D(n1213), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][6]  (.Q(\ram[39][6] ), 
	.D(n1212), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][5]  (.Q(\ram[39][5] ), 
	.D(n1211), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][4]  (.Q(\ram[39][4] ), 
	.D(n1210), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][3]  (.Q(\ram[39][3] ), 
	.D(n1209), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][2]  (.Q(\ram[39][2] ), 
	.D(n1208), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][1]  (.Q(\ram[39][1] ), 
	.D(n1207), 
	.CK(clk));
   DFFHQX1 \ram_reg[39][0]  (.Q(\ram[39][0] ), 
	.D(n1206), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][15]  (.Q(\ram[35][15] ), 
	.D(n1157), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][14]  (.Q(\ram[35][14] ), 
	.D(n1156), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][13]  (.Q(\ram[35][13] ), 
	.D(n1155), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][12]  (.Q(\ram[35][12] ), 
	.D(n1154), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][11]  (.Q(\ram[35][11] ), 
	.D(n1153), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][10]  (.Q(\ram[35][10] ), 
	.D(n1152), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][9]  (.Q(\ram[35][9] ), 
	.D(n1151), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][8]  (.Q(\ram[35][8] ), 
	.D(n1150), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][7]  (.Q(\ram[35][7] ), 
	.D(n1149), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][6]  (.Q(\ram[35][6] ), 
	.D(n1148), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][5]  (.Q(\ram[35][5] ), 
	.D(n1147), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][4]  (.Q(\ram[35][4] ), 
	.D(n1146), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][3]  (.Q(\ram[35][3] ), 
	.D(n1145), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][2]  (.Q(\ram[35][2] ), 
	.D(n1144), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][1]  (.Q(\ram[35][1] ), 
	.D(n1143), 
	.CK(clk));
   DFFHQX1 \ram_reg[35][0]  (.Q(\ram[35][0] ), 
	.D(n1142), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][15]  (.Q(\ram[31][15] ), 
	.D(n1093), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][14]  (.Q(\ram[31][14] ), 
	.D(n1092), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][13]  (.Q(\ram[31][13] ), 
	.D(n1091), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][12]  (.Q(\ram[31][12] ), 
	.D(n1090), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][11]  (.Q(\ram[31][11] ), 
	.D(n1089), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][10]  (.Q(\ram[31][10] ), 
	.D(n1088), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][9]  (.Q(\ram[31][9] ), 
	.D(n1087), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][8]  (.Q(\ram[31][8] ), 
	.D(n1086), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][7]  (.Q(\ram[31][7] ), 
	.D(n1085), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][6]  (.Q(\ram[31][6] ), 
	.D(n1084), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][5]  (.Q(\ram[31][5] ), 
	.D(n1083), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][4]  (.Q(\ram[31][4] ), 
	.D(n1082), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][3]  (.Q(\ram[31][3] ), 
	.D(n1081), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][2]  (.Q(\ram[31][2] ), 
	.D(n1080), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][1]  (.Q(\ram[31][1] ), 
	.D(n1079), 
	.CK(clk));
   DFFHQX1 \ram_reg[31][0]  (.Q(\ram[31][0] ), 
	.D(n1078), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][15]  (.Q(\ram[27][15] ), 
	.D(n1029), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][14]  (.Q(\ram[27][14] ), 
	.D(n1028), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][13]  (.Q(\ram[27][13] ), 
	.D(n1027), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][12]  (.Q(\ram[27][12] ), 
	.D(n1026), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][11]  (.Q(\ram[27][11] ), 
	.D(n1025), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][10]  (.Q(\ram[27][10] ), 
	.D(n1024), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][9]  (.Q(\ram[27][9] ), 
	.D(n1023), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][8]  (.Q(\ram[27][8] ), 
	.D(n1022), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][7]  (.Q(\ram[27][7] ), 
	.D(n1021), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][6]  (.Q(\ram[27][6] ), 
	.D(n1020), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][5]  (.Q(\ram[27][5] ), 
	.D(n1019), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][4]  (.Q(\ram[27][4] ), 
	.D(n1018), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][3]  (.Q(\ram[27][3] ), 
	.D(n1017), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][2]  (.Q(\ram[27][2] ), 
	.D(n1016), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][1]  (.Q(\ram[27][1] ), 
	.D(n1015), 
	.CK(clk));
   DFFHQX1 \ram_reg[27][0]  (.Q(\ram[27][0] ), 
	.D(n1014), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][15]  (.Q(\ram[23][15] ), 
	.D(n965), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][14]  (.Q(\ram[23][14] ), 
	.D(n964), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][13]  (.Q(\ram[23][13] ), 
	.D(n963), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][12]  (.Q(\ram[23][12] ), 
	.D(n962), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][11]  (.Q(\ram[23][11] ), 
	.D(n961), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][10]  (.Q(\ram[23][10] ), 
	.D(n960), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][9]  (.Q(\ram[23][9] ), 
	.D(n959), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][8]  (.Q(\ram[23][8] ), 
	.D(n958), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][7]  (.Q(\ram[23][7] ), 
	.D(n957), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][6]  (.Q(\ram[23][6] ), 
	.D(n956), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][5]  (.Q(\ram[23][5] ), 
	.D(n955), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][4]  (.Q(\ram[23][4] ), 
	.D(n954), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][3]  (.Q(\ram[23][3] ), 
	.D(n953), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][2]  (.Q(\ram[23][2] ), 
	.D(n952), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][1]  (.Q(\ram[23][1] ), 
	.D(n951), 
	.CK(clk));
   DFFHQX1 \ram_reg[23][0]  (.Q(\ram[23][0] ), 
	.D(n950), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][15]  (.Q(\ram[19][15] ), 
	.D(n901), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][14]  (.Q(\ram[19][14] ), 
	.D(n900), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][13]  (.Q(\ram[19][13] ), 
	.D(n899), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][12]  (.Q(\ram[19][12] ), 
	.D(n898), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][11]  (.Q(\ram[19][11] ), 
	.D(n897), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][10]  (.Q(\ram[19][10] ), 
	.D(n896), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][9]  (.Q(\ram[19][9] ), 
	.D(n895), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][8]  (.Q(\ram[19][8] ), 
	.D(n894), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][7]  (.Q(\ram[19][7] ), 
	.D(n893), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][6]  (.Q(\ram[19][6] ), 
	.D(n892), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][5]  (.Q(\ram[19][5] ), 
	.D(n891), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][4]  (.Q(\ram[19][4] ), 
	.D(n890), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][3]  (.Q(\ram[19][3] ), 
	.D(n889), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][2]  (.Q(\ram[19][2] ), 
	.D(n888), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][1]  (.Q(\ram[19][1] ), 
	.D(n887), 
	.CK(clk));
   DFFHQX1 \ram_reg[19][0]  (.Q(\ram[19][0] ), 
	.D(n886), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][15]  (.Q(\ram[15][15] ), 
	.D(n837), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][14]  (.Q(\ram[15][14] ), 
	.D(n836), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][13]  (.Q(\ram[15][13] ), 
	.D(n835), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][12]  (.Q(\ram[15][12] ), 
	.D(n834), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][11]  (.Q(\ram[15][11] ), 
	.D(n833), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][10]  (.Q(\ram[15][10] ), 
	.D(n832), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][9]  (.Q(\ram[15][9] ), 
	.D(n831), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][8]  (.Q(\ram[15][8] ), 
	.D(n830), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][7]  (.Q(\ram[15][7] ), 
	.D(n829), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][6]  (.Q(\ram[15][6] ), 
	.D(n828), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][5]  (.Q(\ram[15][5] ), 
	.D(n827), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][4]  (.Q(\ram[15][4] ), 
	.D(n826), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][3]  (.Q(\ram[15][3] ), 
	.D(n825), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][2]  (.Q(\ram[15][2] ), 
	.D(n824), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][1]  (.Q(\ram[15][1] ), 
	.D(n823), 
	.CK(clk));
   DFFHQX1 \ram_reg[15][0]  (.Q(\ram[15][0] ), 
	.D(n822), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][15]  (.Q(\ram[11][15] ), 
	.D(n773), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][14]  (.Q(\ram[11][14] ), 
	.D(n772), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][13]  (.Q(\ram[11][13] ), 
	.D(n771), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][12]  (.Q(\ram[11][12] ), 
	.D(n770), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][11]  (.Q(\ram[11][11] ), 
	.D(n769), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][10]  (.Q(\ram[11][10] ), 
	.D(n768), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][9]  (.Q(\ram[11][9] ), 
	.D(n767), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][8]  (.Q(\ram[11][8] ), 
	.D(n766), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][7]  (.Q(\ram[11][7] ), 
	.D(n765), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][6]  (.Q(\ram[11][6] ), 
	.D(n764), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][5]  (.Q(\ram[11][5] ), 
	.D(n763), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][4]  (.Q(\ram[11][4] ), 
	.D(n762), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][3]  (.Q(\ram[11][3] ), 
	.D(n761), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][2]  (.Q(\ram[11][2] ), 
	.D(n760), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][1]  (.Q(\ram[11][1] ), 
	.D(n759), 
	.CK(clk));
   DFFHQX1 \ram_reg[11][0]  (.Q(\ram[11][0] ), 
	.D(n758), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][15]  (.Q(\ram[7][15] ), 
	.D(n709), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][14]  (.Q(\ram[7][14] ), 
	.D(n708), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][13]  (.Q(\ram[7][13] ), 
	.D(n707), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][12]  (.Q(\ram[7][12] ), 
	.D(n706), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][11]  (.Q(\ram[7][11] ), 
	.D(n705), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][10]  (.Q(\ram[7][10] ), 
	.D(n704), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][9]  (.Q(\ram[7][9] ), 
	.D(n703), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][8]  (.Q(\ram[7][8] ), 
	.D(n702), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][7]  (.Q(\ram[7][7] ), 
	.D(n701), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][6]  (.Q(\ram[7][6] ), 
	.D(n700), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][5]  (.Q(\ram[7][5] ), 
	.D(n699), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][4]  (.Q(\ram[7][4] ), 
	.D(n698), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][3]  (.Q(\ram[7][3] ), 
	.D(n697), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][2]  (.Q(\ram[7][2] ), 
	.D(n696), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][1]  (.Q(\ram[7][1] ), 
	.D(n695), 
	.CK(clk));
   DFFHQX1 \ram_reg[7][0]  (.Q(\ram[7][0] ), 
	.D(n694), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][15]  (.Q(\ram[3][15] ), 
	.D(n645), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][14]  (.Q(\ram[3][14] ), 
	.D(n644), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][13]  (.Q(\ram[3][13] ), 
	.D(n643), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][12]  (.Q(\ram[3][12] ), 
	.D(n642), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][11]  (.Q(\ram[3][11] ), 
	.D(n641), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][10]  (.Q(\ram[3][10] ), 
	.D(n640), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][9]  (.Q(\ram[3][9] ), 
	.D(n639), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][8]  (.Q(\ram[3][8] ), 
	.D(n638), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][7]  (.Q(\ram[3][7] ), 
	.D(n637), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][6]  (.Q(\ram[3][6] ), 
	.D(n636), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][5]  (.Q(\ram[3][5] ), 
	.D(n635), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][4]  (.Q(\ram[3][4] ), 
	.D(n634), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][3]  (.Q(\ram[3][3] ), 
	.D(n633), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][2]  (.Q(\ram[3][2] ), 
	.D(n632), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][1]  (.Q(\ram[3][1] ), 
	.D(n631), 
	.CK(clk));
   DFFHQX1 \ram_reg[3][0]  (.Q(\ram[3][0] ), 
	.D(n630), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][15]  (.Q(\ram[252][15] ), 
	.D(n4629), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][14]  (.Q(\ram[252][14] ), 
	.D(n4628), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][13]  (.Q(\ram[252][13] ), 
	.D(n4627), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][12]  (.Q(\ram[252][12] ), 
	.D(n4626), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][11]  (.Q(\ram[252][11] ), 
	.D(n4625), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][10]  (.Q(\ram[252][10] ), 
	.D(n4624), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][9]  (.Q(\ram[252][9] ), 
	.D(n4623), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][8]  (.Q(\ram[252][8] ), 
	.D(n4622), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][7]  (.Q(\ram[252][7] ), 
	.D(n4621), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][6]  (.Q(\ram[252][6] ), 
	.D(n4620), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][5]  (.Q(\ram[252][5] ), 
	.D(n4619), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][4]  (.Q(\ram[252][4] ), 
	.D(n4618), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][3]  (.Q(\ram[252][3] ), 
	.D(n4617), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][2]  (.Q(\ram[252][2] ), 
	.D(n4616), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][1]  (.Q(\ram[252][1] ), 
	.D(n4615), 
	.CK(clk));
   DFFHQX1 \ram_reg[252][0]  (.Q(\ram[252][0] ), 
	.D(n4614), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][15]  (.Q(\ram[248][15] ), 
	.D(n4565), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][14]  (.Q(\ram[248][14] ), 
	.D(n4564), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][13]  (.Q(\ram[248][13] ), 
	.D(n4563), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][12]  (.Q(\ram[248][12] ), 
	.D(n4562), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][11]  (.Q(\ram[248][11] ), 
	.D(n4561), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][10]  (.Q(\ram[248][10] ), 
	.D(n4560), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][9]  (.Q(\ram[248][9] ), 
	.D(n4559), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][8]  (.Q(\ram[248][8] ), 
	.D(n4558), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][7]  (.Q(\ram[248][7] ), 
	.D(n4557), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][6]  (.Q(\ram[248][6] ), 
	.D(n4556), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][5]  (.Q(\ram[248][5] ), 
	.D(n4555), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][4]  (.Q(\ram[248][4] ), 
	.D(n4554), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][3]  (.Q(\ram[248][3] ), 
	.D(n4553), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][2]  (.Q(\ram[248][2] ), 
	.D(n4552), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][1]  (.Q(\ram[248][1] ), 
	.D(n4551), 
	.CK(clk));
   DFFHQX1 \ram_reg[248][0]  (.Q(\ram[248][0] ), 
	.D(n4550), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][15]  (.Q(\ram[244][15] ), 
	.D(n4501), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][14]  (.Q(\ram[244][14] ), 
	.D(n4500), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][13]  (.Q(\ram[244][13] ), 
	.D(n4499), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][12]  (.Q(\ram[244][12] ), 
	.D(n4498), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][11]  (.Q(\ram[244][11] ), 
	.D(n4497), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][10]  (.Q(\ram[244][10] ), 
	.D(n4496), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][9]  (.Q(\ram[244][9] ), 
	.D(n4495), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][8]  (.Q(\ram[244][8] ), 
	.D(n4494), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][7]  (.Q(\ram[244][7] ), 
	.D(n4493), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][6]  (.Q(\ram[244][6] ), 
	.D(n4492), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][5]  (.Q(\ram[244][5] ), 
	.D(n4491), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][4]  (.Q(\ram[244][4] ), 
	.D(n4490), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][3]  (.Q(\ram[244][3] ), 
	.D(n4489), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][2]  (.Q(\ram[244][2] ), 
	.D(n4488), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][1]  (.Q(\ram[244][1] ), 
	.D(n4487), 
	.CK(clk));
   DFFHQX1 \ram_reg[244][0]  (.Q(\ram[244][0] ), 
	.D(n4486), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][15]  (.Q(\ram[240][15] ), 
	.D(n4437), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][14]  (.Q(\ram[240][14] ), 
	.D(n4436), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][13]  (.Q(\ram[240][13] ), 
	.D(n4435), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][12]  (.Q(\ram[240][12] ), 
	.D(n4434), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][11]  (.Q(\ram[240][11] ), 
	.D(n4433), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][10]  (.Q(\ram[240][10] ), 
	.D(n4432), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][9]  (.Q(\ram[240][9] ), 
	.D(n4431), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][8]  (.Q(\ram[240][8] ), 
	.D(n4430), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][7]  (.Q(\ram[240][7] ), 
	.D(n4429), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][6]  (.Q(\ram[240][6] ), 
	.D(n4428), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][5]  (.Q(\ram[240][5] ), 
	.D(n4427), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][4]  (.Q(\ram[240][4] ), 
	.D(n4426), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][3]  (.Q(\ram[240][3] ), 
	.D(n4425), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][2]  (.Q(\ram[240][2] ), 
	.D(n4424), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][1]  (.Q(\ram[240][1] ), 
	.D(n4423), 
	.CK(clk));
   DFFHQX1 \ram_reg[240][0]  (.Q(\ram[240][0] ), 
	.D(n4422), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][15]  (.Q(\ram[236][15] ), 
	.D(n4373), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][14]  (.Q(\ram[236][14] ), 
	.D(n4372), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][13]  (.Q(\ram[236][13] ), 
	.D(n4371), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][12]  (.Q(\ram[236][12] ), 
	.D(n4370), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][11]  (.Q(\ram[236][11] ), 
	.D(n4369), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][10]  (.Q(\ram[236][10] ), 
	.D(n4368), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][9]  (.Q(\ram[236][9] ), 
	.D(n4367), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][8]  (.Q(\ram[236][8] ), 
	.D(n4366), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][7]  (.Q(\ram[236][7] ), 
	.D(n4365), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][6]  (.Q(\ram[236][6] ), 
	.D(n4364), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][5]  (.Q(\ram[236][5] ), 
	.D(n4363), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][4]  (.Q(\ram[236][4] ), 
	.D(n4362), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][3]  (.Q(\ram[236][3] ), 
	.D(n4361), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][2]  (.Q(\ram[236][2] ), 
	.D(n4360), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][1]  (.Q(\ram[236][1] ), 
	.D(n4359), 
	.CK(clk));
   DFFHQX1 \ram_reg[236][0]  (.Q(\ram[236][0] ), 
	.D(n4358), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][15]  (.Q(\ram[232][15] ), 
	.D(n4309), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][14]  (.Q(\ram[232][14] ), 
	.D(n4308), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][13]  (.Q(\ram[232][13] ), 
	.D(n4307), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][12]  (.Q(\ram[232][12] ), 
	.D(n4306), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][11]  (.Q(\ram[232][11] ), 
	.D(n4305), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][10]  (.Q(\ram[232][10] ), 
	.D(n4304), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][9]  (.Q(\ram[232][9] ), 
	.D(n4303), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][8]  (.Q(\ram[232][8] ), 
	.D(n4302), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][7]  (.Q(\ram[232][7] ), 
	.D(n4301), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][6]  (.Q(\ram[232][6] ), 
	.D(n4300), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][5]  (.Q(\ram[232][5] ), 
	.D(n4299), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][4]  (.Q(\ram[232][4] ), 
	.D(n4298), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][3]  (.Q(\ram[232][3] ), 
	.D(n4297), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][2]  (.Q(\ram[232][2] ), 
	.D(n4296), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][1]  (.Q(\ram[232][1] ), 
	.D(n4295), 
	.CK(clk));
   DFFHQX1 \ram_reg[232][0]  (.Q(\ram[232][0] ), 
	.D(n4294), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][15]  (.Q(\ram[228][15] ), 
	.D(n4245), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][14]  (.Q(\ram[228][14] ), 
	.D(n4244), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][13]  (.Q(\ram[228][13] ), 
	.D(n4243), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][12]  (.Q(\ram[228][12] ), 
	.D(n4242), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][11]  (.Q(\ram[228][11] ), 
	.D(n4241), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][10]  (.Q(\ram[228][10] ), 
	.D(n4240), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][9]  (.Q(\ram[228][9] ), 
	.D(n4239), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][8]  (.Q(\ram[228][8] ), 
	.D(n4238), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][7]  (.Q(\ram[228][7] ), 
	.D(n4237), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][6]  (.Q(\ram[228][6] ), 
	.D(n4236), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][5]  (.Q(\ram[228][5] ), 
	.D(n4235), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][4]  (.Q(\ram[228][4] ), 
	.D(n4234), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][3]  (.Q(\ram[228][3] ), 
	.D(n4233), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][2]  (.Q(\ram[228][2] ), 
	.D(n4232), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][1]  (.Q(\ram[228][1] ), 
	.D(n4231), 
	.CK(clk));
   DFFHQX1 \ram_reg[228][0]  (.Q(\ram[228][0] ), 
	.D(n4230), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][15]  (.Q(\ram[224][15] ), 
	.D(n4181), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][14]  (.Q(\ram[224][14] ), 
	.D(n4180), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][13]  (.Q(\ram[224][13] ), 
	.D(n4179), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][12]  (.Q(\ram[224][12] ), 
	.D(n4178), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][11]  (.Q(\ram[224][11] ), 
	.D(n4177), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][10]  (.Q(\ram[224][10] ), 
	.D(n4176), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][9]  (.Q(\ram[224][9] ), 
	.D(n4175), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][8]  (.Q(\ram[224][8] ), 
	.D(n4174), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][7]  (.Q(\ram[224][7] ), 
	.D(n4173), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][6]  (.Q(\ram[224][6] ), 
	.D(n4172), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][5]  (.Q(\ram[224][5] ), 
	.D(n4171), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][4]  (.Q(\ram[224][4] ), 
	.D(n4170), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][3]  (.Q(\ram[224][3] ), 
	.D(n4169), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][2]  (.Q(\ram[224][2] ), 
	.D(n4168), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][1]  (.Q(\ram[224][1] ), 
	.D(n4167), 
	.CK(clk));
   DFFHQX1 \ram_reg[224][0]  (.Q(\ram[224][0] ), 
	.D(n4166), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][15]  (.Q(\ram[220][15] ), 
	.D(n4117), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][14]  (.Q(\ram[220][14] ), 
	.D(n4116), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][13]  (.Q(\ram[220][13] ), 
	.D(n4115), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][12]  (.Q(\ram[220][12] ), 
	.D(n4114), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][11]  (.Q(\ram[220][11] ), 
	.D(n4113), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][10]  (.Q(\ram[220][10] ), 
	.D(n4112), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][9]  (.Q(\ram[220][9] ), 
	.D(n4111), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][8]  (.Q(\ram[220][8] ), 
	.D(n4110), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][7]  (.Q(\ram[220][7] ), 
	.D(n4109), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][6]  (.Q(\ram[220][6] ), 
	.D(n4108), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][5]  (.Q(\ram[220][5] ), 
	.D(n4107), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][4]  (.Q(\ram[220][4] ), 
	.D(n4106), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][3]  (.Q(\ram[220][3] ), 
	.D(n4105), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][2]  (.Q(\ram[220][2] ), 
	.D(n4104), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][1]  (.Q(\ram[220][1] ), 
	.D(n4103), 
	.CK(clk));
   DFFHQX1 \ram_reg[220][0]  (.Q(\ram[220][0] ), 
	.D(n4102), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][15]  (.Q(\ram[216][15] ), 
	.D(n4053), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][14]  (.Q(\ram[216][14] ), 
	.D(n4052), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][13]  (.Q(\ram[216][13] ), 
	.D(n4051), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][12]  (.Q(\ram[216][12] ), 
	.D(n4050), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][11]  (.Q(\ram[216][11] ), 
	.D(n4049), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][10]  (.Q(\ram[216][10] ), 
	.D(n4048), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][9]  (.Q(\ram[216][9] ), 
	.D(n4047), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][8]  (.Q(\ram[216][8] ), 
	.D(n4046), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][7]  (.Q(\ram[216][7] ), 
	.D(n4045), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][6]  (.Q(\ram[216][6] ), 
	.D(n4044), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][5]  (.Q(\ram[216][5] ), 
	.D(n4043), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][4]  (.Q(\ram[216][4] ), 
	.D(n4042), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][3]  (.Q(\ram[216][3] ), 
	.D(n4041), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][2]  (.Q(\ram[216][2] ), 
	.D(n4040), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][1]  (.Q(\ram[216][1] ), 
	.D(n4039), 
	.CK(clk));
   DFFHQX1 \ram_reg[216][0]  (.Q(\ram[216][0] ), 
	.D(n4038), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][15]  (.Q(\ram[212][15] ), 
	.D(n3989), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][14]  (.Q(\ram[212][14] ), 
	.D(n3988), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][13]  (.Q(\ram[212][13] ), 
	.D(n3987), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][12]  (.Q(\ram[212][12] ), 
	.D(n3986), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][11]  (.Q(\ram[212][11] ), 
	.D(n3985), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][10]  (.Q(\ram[212][10] ), 
	.D(n3984), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][9]  (.Q(\ram[212][9] ), 
	.D(n3983), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][8]  (.Q(\ram[212][8] ), 
	.D(n3982), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][7]  (.Q(\ram[212][7] ), 
	.D(n3981), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][6]  (.Q(\ram[212][6] ), 
	.D(n3980), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][5]  (.Q(\ram[212][5] ), 
	.D(n3979), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][4]  (.Q(\ram[212][4] ), 
	.D(n3978), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][3]  (.Q(\ram[212][3] ), 
	.D(n3977), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][2]  (.Q(\ram[212][2] ), 
	.D(n3976), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][1]  (.Q(\ram[212][1] ), 
	.D(n3975), 
	.CK(clk));
   DFFHQX1 \ram_reg[212][0]  (.Q(\ram[212][0] ), 
	.D(n3974), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][15]  (.Q(\ram[208][15] ), 
	.D(n3925), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][14]  (.Q(\ram[208][14] ), 
	.D(n3924), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][13]  (.Q(\ram[208][13] ), 
	.D(n3923), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][12]  (.Q(\ram[208][12] ), 
	.D(n3922), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][11]  (.Q(\ram[208][11] ), 
	.D(n3921), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][10]  (.Q(\ram[208][10] ), 
	.D(n3920), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][9]  (.Q(\ram[208][9] ), 
	.D(n3919), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][8]  (.Q(\ram[208][8] ), 
	.D(n3918), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][7]  (.Q(\ram[208][7] ), 
	.D(n3917), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][6]  (.Q(\ram[208][6] ), 
	.D(n3916), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][5]  (.Q(\ram[208][5] ), 
	.D(n3915), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][4]  (.Q(\ram[208][4] ), 
	.D(n3914), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][3]  (.Q(\ram[208][3] ), 
	.D(n3913), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][2]  (.Q(\ram[208][2] ), 
	.D(n3912), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][1]  (.Q(\ram[208][1] ), 
	.D(n3911), 
	.CK(clk));
   DFFHQX1 \ram_reg[208][0]  (.Q(\ram[208][0] ), 
	.D(n3910), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][15]  (.Q(\ram[204][15] ), 
	.D(n3861), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][14]  (.Q(\ram[204][14] ), 
	.D(n3860), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][13]  (.Q(\ram[204][13] ), 
	.D(n3859), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][12]  (.Q(\ram[204][12] ), 
	.D(n3858), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][11]  (.Q(\ram[204][11] ), 
	.D(n3857), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][10]  (.Q(\ram[204][10] ), 
	.D(n3856), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][9]  (.Q(\ram[204][9] ), 
	.D(n3855), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][8]  (.Q(\ram[204][8] ), 
	.D(n3854), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][7]  (.Q(\ram[204][7] ), 
	.D(n3853), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][6]  (.Q(\ram[204][6] ), 
	.D(n3852), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][5]  (.Q(\ram[204][5] ), 
	.D(n3851), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][4]  (.Q(\ram[204][4] ), 
	.D(n3850), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][3]  (.Q(\ram[204][3] ), 
	.D(n3849), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][2]  (.Q(\ram[204][2] ), 
	.D(n3848), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][1]  (.Q(\ram[204][1] ), 
	.D(n3847), 
	.CK(clk));
   DFFHQX1 \ram_reg[204][0]  (.Q(\ram[204][0] ), 
	.D(n3846), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][15]  (.Q(\ram[200][15] ), 
	.D(n3797), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][14]  (.Q(\ram[200][14] ), 
	.D(n3796), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][13]  (.Q(\ram[200][13] ), 
	.D(n3795), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][12]  (.Q(\ram[200][12] ), 
	.D(n3794), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][11]  (.Q(\ram[200][11] ), 
	.D(n3793), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][10]  (.Q(\ram[200][10] ), 
	.D(n3792), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][9]  (.Q(\ram[200][9] ), 
	.D(n3791), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][8]  (.Q(\ram[200][8] ), 
	.D(n3790), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][7]  (.Q(\ram[200][7] ), 
	.D(n3789), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][6]  (.Q(\ram[200][6] ), 
	.D(n3788), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][5]  (.Q(\ram[200][5] ), 
	.D(n3787), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][4]  (.Q(\ram[200][4] ), 
	.D(n3786), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][3]  (.Q(\ram[200][3] ), 
	.D(n3785), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][2]  (.Q(\ram[200][2] ), 
	.D(n3784), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][1]  (.Q(\ram[200][1] ), 
	.D(n3783), 
	.CK(clk));
   DFFHQX1 \ram_reg[200][0]  (.Q(\ram[200][0] ), 
	.D(n3782), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][15]  (.Q(\ram[196][15] ), 
	.D(n3733), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][14]  (.Q(\ram[196][14] ), 
	.D(n3732), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][13]  (.Q(\ram[196][13] ), 
	.D(n3731), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][12]  (.Q(\ram[196][12] ), 
	.D(n3730), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][11]  (.Q(\ram[196][11] ), 
	.D(n3729), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][10]  (.Q(\ram[196][10] ), 
	.D(n3728), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][9]  (.Q(\ram[196][9] ), 
	.D(n3727), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][8]  (.Q(\ram[196][8] ), 
	.D(n3726), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][7]  (.Q(\ram[196][7] ), 
	.D(n3725), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][6]  (.Q(\ram[196][6] ), 
	.D(n3724), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][5]  (.Q(\ram[196][5] ), 
	.D(n3723), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][4]  (.Q(\ram[196][4] ), 
	.D(n3722), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][3]  (.Q(\ram[196][3] ), 
	.D(n3721), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][2]  (.Q(\ram[196][2] ), 
	.D(n3720), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][1]  (.Q(\ram[196][1] ), 
	.D(n3719), 
	.CK(clk));
   DFFHQX1 \ram_reg[196][0]  (.Q(\ram[196][0] ), 
	.D(n3718), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][15]  (.Q(\ram[192][15] ), 
	.D(n3669), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][14]  (.Q(\ram[192][14] ), 
	.D(n3668), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][13]  (.Q(\ram[192][13] ), 
	.D(n3667), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][12]  (.Q(\ram[192][12] ), 
	.D(n3666), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][11]  (.Q(\ram[192][11] ), 
	.D(n3665), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][10]  (.Q(\ram[192][10] ), 
	.D(n3664), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][9]  (.Q(\ram[192][9] ), 
	.D(n3663), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][8]  (.Q(\ram[192][8] ), 
	.D(n3662), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][7]  (.Q(\ram[192][7] ), 
	.D(n3661), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][6]  (.Q(\ram[192][6] ), 
	.D(n3660), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][5]  (.Q(\ram[192][5] ), 
	.D(n3659), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][4]  (.Q(\ram[192][4] ), 
	.D(n3658), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][3]  (.Q(\ram[192][3] ), 
	.D(n3657), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][2]  (.Q(\ram[192][2] ), 
	.D(n3656), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][1]  (.Q(\ram[192][1] ), 
	.D(n3655), 
	.CK(clk));
   DFFHQX1 \ram_reg[192][0]  (.Q(\ram[192][0] ), 
	.D(n3654), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][15]  (.Q(\ram[188][15] ), 
	.D(n3605), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][14]  (.Q(\ram[188][14] ), 
	.D(n3604), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][13]  (.Q(\ram[188][13] ), 
	.D(n3603), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][12]  (.Q(\ram[188][12] ), 
	.D(n3602), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][11]  (.Q(\ram[188][11] ), 
	.D(n3601), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][10]  (.Q(\ram[188][10] ), 
	.D(n3600), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][9]  (.Q(\ram[188][9] ), 
	.D(n3599), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][8]  (.Q(\ram[188][8] ), 
	.D(n3598), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][7]  (.Q(\ram[188][7] ), 
	.D(n3597), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][6]  (.Q(\ram[188][6] ), 
	.D(n3596), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][5]  (.Q(\ram[188][5] ), 
	.D(n3595), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][4]  (.Q(\ram[188][4] ), 
	.D(n3594), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][3]  (.Q(\ram[188][3] ), 
	.D(n3593), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][2]  (.Q(\ram[188][2] ), 
	.D(n3592), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][1]  (.Q(\ram[188][1] ), 
	.D(n3591), 
	.CK(clk));
   DFFHQX1 \ram_reg[188][0]  (.Q(\ram[188][0] ), 
	.D(n3590), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][15]  (.Q(\ram[184][15] ), 
	.D(n3541), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][14]  (.Q(\ram[184][14] ), 
	.D(n3540), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][13]  (.Q(\ram[184][13] ), 
	.D(n3539), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][12]  (.Q(\ram[184][12] ), 
	.D(n3538), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][11]  (.Q(\ram[184][11] ), 
	.D(n3537), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][10]  (.Q(\ram[184][10] ), 
	.D(n3536), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][9]  (.Q(\ram[184][9] ), 
	.D(n3535), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][8]  (.Q(\ram[184][8] ), 
	.D(n3534), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][7]  (.Q(\ram[184][7] ), 
	.D(n3533), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][6]  (.Q(\ram[184][6] ), 
	.D(n3532), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][5]  (.Q(\ram[184][5] ), 
	.D(n3531), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][4]  (.Q(\ram[184][4] ), 
	.D(n3530), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][3]  (.Q(\ram[184][3] ), 
	.D(n3529), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][2]  (.Q(\ram[184][2] ), 
	.D(n3528), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][1]  (.Q(\ram[184][1] ), 
	.D(n3527), 
	.CK(clk));
   DFFHQX1 \ram_reg[184][0]  (.Q(\ram[184][0] ), 
	.D(n3526), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][15]  (.Q(\ram[180][15] ), 
	.D(n3477), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][14]  (.Q(\ram[180][14] ), 
	.D(n3476), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][13]  (.Q(\ram[180][13] ), 
	.D(n3475), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][12]  (.Q(\ram[180][12] ), 
	.D(n3474), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][11]  (.Q(\ram[180][11] ), 
	.D(n3473), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][10]  (.Q(\ram[180][10] ), 
	.D(n3472), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][9]  (.Q(\ram[180][9] ), 
	.D(n3471), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][8]  (.Q(\ram[180][8] ), 
	.D(n3470), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][7]  (.Q(\ram[180][7] ), 
	.D(n3469), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][6]  (.Q(\ram[180][6] ), 
	.D(n3468), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][5]  (.Q(\ram[180][5] ), 
	.D(n3467), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][4]  (.Q(\ram[180][4] ), 
	.D(n3466), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][3]  (.Q(\ram[180][3] ), 
	.D(n3465), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][2]  (.Q(\ram[180][2] ), 
	.D(n3464), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][1]  (.Q(\ram[180][1] ), 
	.D(n3463), 
	.CK(clk));
   DFFHQX1 \ram_reg[180][0]  (.Q(\ram[180][0] ), 
	.D(n3462), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][15]  (.Q(\ram[176][15] ), 
	.D(n3413), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][14]  (.Q(\ram[176][14] ), 
	.D(n3412), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][13]  (.Q(\ram[176][13] ), 
	.D(n3411), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][12]  (.Q(\ram[176][12] ), 
	.D(n3410), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][11]  (.Q(\ram[176][11] ), 
	.D(n3409), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][10]  (.Q(\ram[176][10] ), 
	.D(n3408), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][9]  (.Q(\ram[176][9] ), 
	.D(n3407), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][8]  (.Q(\ram[176][8] ), 
	.D(n3406), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][7]  (.Q(\ram[176][7] ), 
	.D(n3405), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][6]  (.Q(\ram[176][6] ), 
	.D(n3404), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][5]  (.Q(\ram[176][5] ), 
	.D(n3403), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][4]  (.Q(\ram[176][4] ), 
	.D(n3402), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][3]  (.Q(\ram[176][3] ), 
	.D(n3401), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][2]  (.Q(\ram[176][2] ), 
	.D(n3400), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][1]  (.Q(\ram[176][1] ), 
	.D(n3399), 
	.CK(clk));
   DFFHQX1 \ram_reg[176][0]  (.Q(\ram[176][0] ), 
	.D(n3398), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][15]  (.Q(\ram[172][15] ), 
	.D(n3349), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][14]  (.Q(\ram[172][14] ), 
	.D(n3348), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][13]  (.Q(\ram[172][13] ), 
	.D(n3347), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][12]  (.Q(\ram[172][12] ), 
	.D(n3346), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][11]  (.Q(\ram[172][11] ), 
	.D(n3345), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][10]  (.Q(\ram[172][10] ), 
	.D(n3344), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][9]  (.Q(\ram[172][9] ), 
	.D(n3343), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][8]  (.Q(\ram[172][8] ), 
	.D(n3342), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][7]  (.Q(\ram[172][7] ), 
	.D(n3341), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][6]  (.Q(\ram[172][6] ), 
	.D(n3340), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][5]  (.Q(\ram[172][5] ), 
	.D(n3339), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][4]  (.Q(\ram[172][4] ), 
	.D(n3338), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][3]  (.Q(\ram[172][3] ), 
	.D(n3337), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][2]  (.Q(\ram[172][2] ), 
	.D(n3336), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][1]  (.Q(\ram[172][1] ), 
	.D(n3335), 
	.CK(clk));
   DFFHQX1 \ram_reg[172][0]  (.Q(\ram[172][0] ), 
	.D(n3334), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][15]  (.Q(\ram[168][15] ), 
	.D(n3285), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][14]  (.Q(\ram[168][14] ), 
	.D(n3284), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][13]  (.Q(\ram[168][13] ), 
	.D(n3283), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][12]  (.Q(\ram[168][12] ), 
	.D(n3282), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][11]  (.Q(\ram[168][11] ), 
	.D(n3281), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][10]  (.Q(\ram[168][10] ), 
	.D(n3280), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][9]  (.Q(\ram[168][9] ), 
	.D(n3279), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][8]  (.Q(\ram[168][8] ), 
	.D(n3278), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][7]  (.Q(\ram[168][7] ), 
	.D(n3277), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][6]  (.Q(\ram[168][6] ), 
	.D(n3276), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][5]  (.Q(\ram[168][5] ), 
	.D(n3275), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][4]  (.Q(\ram[168][4] ), 
	.D(n3274), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][3]  (.Q(\ram[168][3] ), 
	.D(n3273), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][2]  (.Q(\ram[168][2] ), 
	.D(n3272), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][1]  (.Q(\ram[168][1] ), 
	.D(n3271), 
	.CK(clk));
   DFFHQX1 \ram_reg[168][0]  (.Q(\ram[168][0] ), 
	.D(n3270), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][15]  (.Q(\ram[164][15] ), 
	.D(n3221), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][14]  (.Q(\ram[164][14] ), 
	.D(n3220), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][13]  (.Q(\ram[164][13] ), 
	.D(n3219), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][12]  (.Q(\ram[164][12] ), 
	.D(n3218), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][11]  (.Q(\ram[164][11] ), 
	.D(n3217), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][10]  (.Q(\ram[164][10] ), 
	.D(n3216), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][9]  (.Q(\ram[164][9] ), 
	.D(n3215), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][8]  (.Q(\ram[164][8] ), 
	.D(n3214), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][7]  (.Q(\ram[164][7] ), 
	.D(n3213), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][6]  (.Q(\ram[164][6] ), 
	.D(n3212), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][5]  (.Q(\ram[164][5] ), 
	.D(n3211), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][4]  (.Q(\ram[164][4] ), 
	.D(n3210), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][3]  (.Q(\ram[164][3] ), 
	.D(n3209), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][2]  (.Q(\ram[164][2] ), 
	.D(n3208), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][1]  (.Q(\ram[164][1] ), 
	.D(n3207), 
	.CK(clk));
   DFFHQX1 \ram_reg[164][0]  (.Q(\ram[164][0] ), 
	.D(n3206), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][15]  (.Q(\ram[160][15] ), 
	.D(n3157), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][14]  (.Q(\ram[160][14] ), 
	.D(n3156), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][13]  (.Q(\ram[160][13] ), 
	.D(n3155), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][12]  (.Q(\ram[160][12] ), 
	.D(n3154), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][11]  (.Q(\ram[160][11] ), 
	.D(n3153), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][10]  (.Q(\ram[160][10] ), 
	.D(n3152), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][9]  (.Q(\ram[160][9] ), 
	.D(n3151), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][8]  (.Q(\ram[160][8] ), 
	.D(n3150), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][7]  (.Q(\ram[160][7] ), 
	.D(n3149), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][6]  (.Q(\ram[160][6] ), 
	.D(n3148), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][5]  (.Q(\ram[160][5] ), 
	.D(n3147), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][4]  (.Q(\ram[160][4] ), 
	.D(n3146), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][3]  (.Q(\ram[160][3] ), 
	.D(n3145), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][2]  (.Q(\ram[160][2] ), 
	.D(n3144), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][1]  (.Q(\ram[160][1] ), 
	.D(n3143), 
	.CK(clk));
   DFFHQX1 \ram_reg[160][0]  (.Q(\ram[160][0] ), 
	.D(n3142), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][15]  (.Q(\ram[156][15] ), 
	.D(n3093), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][14]  (.Q(\ram[156][14] ), 
	.D(n3092), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][13]  (.Q(\ram[156][13] ), 
	.D(n3091), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][12]  (.Q(\ram[156][12] ), 
	.D(n3090), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][11]  (.Q(\ram[156][11] ), 
	.D(n3089), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][10]  (.Q(\ram[156][10] ), 
	.D(n3088), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][9]  (.Q(\ram[156][9] ), 
	.D(n3087), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][8]  (.Q(\ram[156][8] ), 
	.D(n3086), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][7]  (.Q(\ram[156][7] ), 
	.D(n3085), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][6]  (.Q(\ram[156][6] ), 
	.D(n3084), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][5]  (.Q(\ram[156][5] ), 
	.D(n3083), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][4]  (.Q(\ram[156][4] ), 
	.D(n3082), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][3]  (.Q(\ram[156][3] ), 
	.D(n3081), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][2]  (.Q(\ram[156][2] ), 
	.D(n3080), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][1]  (.Q(\ram[156][1] ), 
	.D(n3079), 
	.CK(clk));
   DFFHQX1 \ram_reg[156][0]  (.Q(\ram[156][0] ), 
	.D(n3078), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][15]  (.Q(\ram[152][15] ), 
	.D(n3029), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][14]  (.Q(\ram[152][14] ), 
	.D(n3028), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][13]  (.Q(\ram[152][13] ), 
	.D(n3027), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][12]  (.Q(\ram[152][12] ), 
	.D(n3026), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][11]  (.Q(\ram[152][11] ), 
	.D(n3025), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][10]  (.Q(\ram[152][10] ), 
	.D(n3024), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][9]  (.Q(\ram[152][9] ), 
	.D(n3023), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][8]  (.Q(\ram[152][8] ), 
	.D(n3022), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][7]  (.Q(\ram[152][7] ), 
	.D(n3021), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][6]  (.Q(\ram[152][6] ), 
	.D(n3020), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][5]  (.Q(\ram[152][5] ), 
	.D(n3019), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][4]  (.Q(\ram[152][4] ), 
	.D(n3018), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][3]  (.Q(\ram[152][3] ), 
	.D(n3017), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][2]  (.Q(\ram[152][2] ), 
	.D(n3016), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][1]  (.Q(\ram[152][1] ), 
	.D(n3015), 
	.CK(clk));
   DFFHQX1 \ram_reg[152][0]  (.Q(\ram[152][0] ), 
	.D(n3014), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][15]  (.Q(\ram[148][15] ), 
	.D(n2965), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][14]  (.Q(\ram[148][14] ), 
	.D(n2964), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][13]  (.Q(\ram[148][13] ), 
	.D(n2963), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][12]  (.Q(\ram[148][12] ), 
	.D(n2962), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][11]  (.Q(\ram[148][11] ), 
	.D(n2961), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][10]  (.Q(\ram[148][10] ), 
	.D(n2960), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][9]  (.Q(\ram[148][9] ), 
	.D(n2959), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][8]  (.Q(\ram[148][8] ), 
	.D(n2958), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][7]  (.Q(\ram[148][7] ), 
	.D(n2957), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][6]  (.Q(\ram[148][6] ), 
	.D(n2956), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][5]  (.Q(\ram[148][5] ), 
	.D(n2955), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][4]  (.Q(\ram[148][4] ), 
	.D(n2954), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][3]  (.Q(\ram[148][3] ), 
	.D(n2953), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][2]  (.Q(\ram[148][2] ), 
	.D(n2952), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][1]  (.Q(\ram[148][1] ), 
	.D(n2951), 
	.CK(clk));
   DFFHQX1 \ram_reg[148][0]  (.Q(\ram[148][0] ), 
	.D(n2950), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][15]  (.Q(\ram[144][15] ), 
	.D(n2901), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][14]  (.Q(\ram[144][14] ), 
	.D(n2900), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][13]  (.Q(\ram[144][13] ), 
	.D(n2899), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][12]  (.Q(\ram[144][12] ), 
	.D(n2898), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][11]  (.Q(\ram[144][11] ), 
	.D(n2897), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][10]  (.Q(\ram[144][10] ), 
	.D(n2896), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][9]  (.Q(\ram[144][9] ), 
	.D(n2895), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][8]  (.Q(\ram[144][8] ), 
	.D(n2894), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][7]  (.Q(\ram[144][7] ), 
	.D(n2893), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][6]  (.Q(\ram[144][6] ), 
	.D(n2892), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][5]  (.Q(\ram[144][5] ), 
	.D(n2891), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][4]  (.Q(\ram[144][4] ), 
	.D(n2890), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][3]  (.Q(\ram[144][3] ), 
	.D(n2889), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][2]  (.Q(\ram[144][2] ), 
	.D(n2888), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][1]  (.Q(\ram[144][1] ), 
	.D(n2887), 
	.CK(clk));
   DFFHQX1 \ram_reg[144][0]  (.Q(\ram[144][0] ), 
	.D(n2886), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][15]  (.Q(\ram[140][15] ), 
	.D(n2837), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][14]  (.Q(\ram[140][14] ), 
	.D(n2836), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][13]  (.Q(\ram[140][13] ), 
	.D(n2835), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][12]  (.Q(\ram[140][12] ), 
	.D(n2834), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][11]  (.Q(\ram[140][11] ), 
	.D(n2833), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][10]  (.Q(\ram[140][10] ), 
	.D(n2832), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][9]  (.Q(\ram[140][9] ), 
	.D(n2831), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][8]  (.Q(\ram[140][8] ), 
	.D(n2830), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][7]  (.Q(\ram[140][7] ), 
	.D(n2829), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][6]  (.Q(\ram[140][6] ), 
	.D(n2828), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][5]  (.Q(\ram[140][5] ), 
	.D(n2827), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][4]  (.Q(\ram[140][4] ), 
	.D(n2826), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][3]  (.Q(\ram[140][3] ), 
	.D(n2825), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][2]  (.Q(\ram[140][2] ), 
	.D(n2824), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][1]  (.Q(\ram[140][1] ), 
	.D(n2823), 
	.CK(clk));
   DFFHQX1 \ram_reg[140][0]  (.Q(\ram[140][0] ), 
	.D(n2822), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][15]  (.Q(\ram[136][15] ), 
	.D(n2773), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][14]  (.Q(\ram[136][14] ), 
	.D(n2772), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][13]  (.Q(\ram[136][13] ), 
	.D(n2771), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][12]  (.Q(\ram[136][12] ), 
	.D(n2770), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][11]  (.Q(\ram[136][11] ), 
	.D(n2769), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][10]  (.Q(\ram[136][10] ), 
	.D(n2768), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][9]  (.Q(\ram[136][9] ), 
	.D(n2767), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][8]  (.Q(\ram[136][8] ), 
	.D(n2766), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][7]  (.Q(\ram[136][7] ), 
	.D(n2765), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][6]  (.Q(\ram[136][6] ), 
	.D(n2764), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][5]  (.Q(\ram[136][5] ), 
	.D(n2763), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][4]  (.Q(\ram[136][4] ), 
	.D(n2762), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][3]  (.Q(\ram[136][3] ), 
	.D(n2761), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][2]  (.Q(\ram[136][2] ), 
	.D(n2760), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][1]  (.Q(\ram[136][1] ), 
	.D(n2759), 
	.CK(clk));
   DFFHQX1 \ram_reg[136][0]  (.Q(\ram[136][0] ), 
	.D(n2758), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][15]  (.Q(\ram[132][15] ), 
	.D(n2709), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][14]  (.Q(\ram[132][14] ), 
	.D(n2708), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][13]  (.Q(\ram[132][13] ), 
	.D(n2707), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][12]  (.Q(\ram[132][12] ), 
	.D(n2706), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][11]  (.Q(\ram[132][11] ), 
	.D(n2705), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][10]  (.Q(\ram[132][10] ), 
	.D(n2704), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][9]  (.Q(\ram[132][9] ), 
	.D(n2703), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][8]  (.Q(\ram[132][8] ), 
	.D(n2702), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][7]  (.Q(\ram[132][7] ), 
	.D(n2701), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][6]  (.Q(\ram[132][6] ), 
	.D(n2700), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][5]  (.Q(\ram[132][5] ), 
	.D(n2699), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][4]  (.Q(\ram[132][4] ), 
	.D(n2698), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][3]  (.Q(\ram[132][3] ), 
	.D(n2697), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][2]  (.Q(\ram[132][2] ), 
	.D(n2696), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][1]  (.Q(\ram[132][1] ), 
	.D(n2695), 
	.CK(clk));
   DFFHQX1 \ram_reg[132][0]  (.Q(\ram[132][0] ), 
	.D(n2694), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][15]  (.Q(\ram[128][15] ), 
	.D(n2645), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][14]  (.Q(\ram[128][14] ), 
	.D(n2644), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][13]  (.Q(\ram[128][13] ), 
	.D(n2643), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][12]  (.Q(\ram[128][12] ), 
	.D(n2642), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][11]  (.Q(\ram[128][11] ), 
	.D(n2641), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][10]  (.Q(\ram[128][10] ), 
	.D(n2640), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][9]  (.Q(\ram[128][9] ), 
	.D(n2639), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][8]  (.Q(\ram[128][8] ), 
	.D(n2638), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][7]  (.Q(\ram[128][7] ), 
	.D(n2637), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][6]  (.Q(\ram[128][6] ), 
	.D(n2636), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][5]  (.Q(\ram[128][5] ), 
	.D(n2635), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][4]  (.Q(\ram[128][4] ), 
	.D(n2634), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][3]  (.Q(\ram[128][3] ), 
	.D(n2633), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][2]  (.Q(\ram[128][2] ), 
	.D(n2632), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][1]  (.Q(\ram[128][1] ), 
	.D(n2631), 
	.CK(clk));
   DFFHQX1 \ram_reg[128][0]  (.Q(\ram[128][0] ), 
	.D(n2630), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][15]  (.Q(\ram[124][15] ), 
	.D(n2581), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][14]  (.Q(\ram[124][14] ), 
	.D(n2580), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][13]  (.Q(\ram[124][13] ), 
	.D(n2579), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][12]  (.Q(\ram[124][12] ), 
	.D(n2578), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][11]  (.Q(\ram[124][11] ), 
	.D(n2577), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][10]  (.Q(\ram[124][10] ), 
	.D(n2576), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][9]  (.Q(\ram[124][9] ), 
	.D(n2575), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][8]  (.Q(\ram[124][8] ), 
	.D(n2574), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][7]  (.Q(\ram[124][7] ), 
	.D(n2573), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][6]  (.Q(\ram[124][6] ), 
	.D(n2572), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][5]  (.Q(\ram[124][5] ), 
	.D(n2571), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][4]  (.Q(\ram[124][4] ), 
	.D(n2570), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][3]  (.Q(\ram[124][3] ), 
	.D(n2569), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][2]  (.Q(\ram[124][2] ), 
	.D(n2568), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][1]  (.Q(\ram[124][1] ), 
	.D(n2567), 
	.CK(clk));
   DFFHQX1 \ram_reg[124][0]  (.Q(\ram[124][0] ), 
	.D(n2566), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][15]  (.Q(\ram[120][15] ), 
	.D(n2517), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][14]  (.Q(\ram[120][14] ), 
	.D(n2516), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][13]  (.Q(\ram[120][13] ), 
	.D(n2515), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][12]  (.Q(\ram[120][12] ), 
	.D(n2514), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][11]  (.Q(\ram[120][11] ), 
	.D(n2513), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][10]  (.Q(\ram[120][10] ), 
	.D(n2512), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][9]  (.Q(\ram[120][9] ), 
	.D(n2511), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][8]  (.Q(\ram[120][8] ), 
	.D(n2510), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][7]  (.Q(\ram[120][7] ), 
	.D(n2509), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][6]  (.Q(\ram[120][6] ), 
	.D(n2508), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][5]  (.Q(\ram[120][5] ), 
	.D(n2507), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][4]  (.Q(\ram[120][4] ), 
	.D(n2506), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][3]  (.Q(\ram[120][3] ), 
	.D(n2505), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][2]  (.Q(\ram[120][2] ), 
	.D(n2504), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][1]  (.Q(\ram[120][1] ), 
	.D(n2503), 
	.CK(clk));
   DFFHQX1 \ram_reg[120][0]  (.Q(\ram[120][0] ), 
	.D(n2502), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][15]  (.Q(\ram[116][15] ), 
	.D(n2453), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][14]  (.Q(\ram[116][14] ), 
	.D(n2452), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][13]  (.Q(\ram[116][13] ), 
	.D(n2451), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][12]  (.Q(\ram[116][12] ), 
	.D(n2450), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][11]  (.Q(\ram[116][11] ), 
	.D(n2449), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][10]  (.Q(\ram[116][10] ), 
	.D(n2448), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][9]  (.Q(\ram[116][9] ), 
	.D(n2447), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][8]  (.Q(\ram[116][8] ), 
	.D(n2446), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][7]  (.Q(\ram[116][7] ), 
	.D(n2445), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][6]  (.Q(\ram[116][6] ), 
	.D(n2444), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][5]  (.Q(\ram[116][5] ), 
	.D(n2443), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][4]  (.Q(\ram[116][4] ), 
	.D(n2442), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][3]  (.Q(\ram[116][3] ), 
	.D(n2441), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][2]  (.Q(\ram[116][2] ), 
	.D(n2440), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][1]  (.Q(\ram[116][1] ), 
	.D(n2439), 
	.CK(clk));
   DFFHQX1 \ram_reg[116][0]  (.Q(\ram[116][0] ), 
	.D(n2438), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][15]  (.Q(\ram[112][15] ), 
	.D(n2389), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][14]  (.Q(\ram[112][14] ), 
	.D(n2388), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][13]  (.Q(\ram[112][13] ), 
	.D(n2387), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][12]  (.Q(\ram[112][12] ), 
	.D(n2386), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][11]  (.Q(\ram[112][11] ), 
	.D(n2385), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][10]  (.Q(\ram[112][10] ), 
	.D(n2384), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][9]  (.Q(\ram[112][9] ), 
	.D(n2383), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][8]  (.Q(\ram[112][8] ), 
	.D(n2382), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][7]  (.Q(\ram[112][7] ), 
	.D(n2381), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][6]  (.Q(\ram[112][6] ), 
	.D(n2380), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][5]  (.Q(\ram[112][5] ), 
	.D(n2379), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][4]  (.Q(\ram[112][4] ), 
	.D(n2378), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][3]  (.Q(\ram[112][3] ), 
	.D(n2377), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][2]  (.Q(\ram[112][2] ), 
	.D(n2376), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][1]  (.Q(\ram[112][1] ), 
	.D(n2375), 
	.CK(clk));
   DFFHQX1 \ram_reg[112][0]  (.Q(\ram[112][0] ), 
	.D(n2374), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][15]  (.Q(\ram[108][15] ), 
	.D(n2325), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][14]  (.Q(\ram[108][14] ), 
	.D(n2324), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][13]  (.Q(\ram[108][13] ), 
	.D(n2323), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][12]  (.Q(\ram[108][12] ), 
	.D(n2322), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][11]  (.Q(\ram[108][11] ), 
	.D(n2321), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][10]  (.Q(\ram[108][10] ), 
	.D(n2320), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][9]  (.Q(\ram[108][9] ), 
	.D(n2319), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][8]  (.Q(\ram[108][8] ), 
	.D(n2318), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][7]  (.Q(\ram[108][7] ), 
	.D(n2317), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][6]  (.Q(\ram[108][6] ), 
	.D(n2316), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][5]  (.Q(\ram[108][5] ), 
	.D(n2315), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][4]  (.Q(\ram[108][4] ), 
	.D(n2314), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][3]  (.Q(\ram[108][3] ), 
	.D(n2313), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][2]  (.Q(\ram[108][2] ), 
	.D(n2312), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][1]  (.Q(\ram[108][1] ), 
	.D(n2311), 
	.CK(clk));
   DFFHQX1 \ram_reg[108][0]  (.Q(\ram[108][0] ), 
	.D(n2310), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][15]  (.Q(\ram[104][15] ), 
	.D(n2261), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][14]  (.Q(\ram[104][14] ), 
	.D(n2260), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][13]  (.Q(\ram[104][13] ), 
	.D(n2259), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][12]  (.Q(\ram[104][12] ), 
	.D(n2258), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][11]  (.Q(\ram[104][11] ), 
	.D(n2257), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][10]  (.Q(\ram[104][10] ), 
	.D(n2256), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][9]  (.Q(\ram[104][9] ), 
	.D(n2255), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][8]  (.Q(\ram[104][8] ), 
	.D(n2254), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][7]  (.Q(\ram[104][7] ), 
	.D(n2253), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][6]  (.Q(\ram[104][6] ), 
	.D(n2252), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][5]  (.Q(\ram[104][5] ), 
	.D(n2251), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][4]  (.Q(\ram[104][4] ), 
	.D(n2250), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][3]  (.Q(\ram[104][3] ), 
	.D(n2249), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][2]  (.Q(\ram[104][2] ), 
	.D(n2248), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][1]  (.Q(\ram[104][1] ), 
	.D(n2247), 
	.CK(clk));
   DFFHQX1 \ram_reg[104][0]  (.Q(\ram[104][0] ), 
	.D(n2246), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][15]  (.Q(\ram[100][15] ), 
	.D(n2197), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][14]  (.Q(\ram[100][14] ), 
	.D(n2196), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][13]  (.Q(\ram[100][13] ), 
	.D(n2195), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][12]  (.Q(\ram[100][12] ), 
	.D(n2194), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][11]  (.Q(\ram[100][11] ), 
	.D(n2193), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][10]  (.Q(\ram[100][10] ), 
	.D(n2192), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][9]  (.Q(\ram[100][9] ), 
	.D(n2191), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][8]  (.Q(\ram[100][8] ), 
	.D(n2190), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][7]  (.Q(\ram[100][7] ), 
	.D(n2189), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][6]  (.Q(\ram[100][6] ), 
	.D(n2188), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][5]  (.Q(\ram[100][5] ), 
	.D(n2187), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][4]  (.Q(\ram[100][4] ), 
	.D(n2186), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][3]  (.Q(\ram[100][3] ), 
	.D(n2185), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][2]  (.Q(\ram[100][2] ), 
	.D(n2184), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][1]  (.Q(\ram[100][1] ), 
	.D(n2183), 
	.CK(clk));
   DFFHQX1 \ram_reg[100][0]  (.Q(\ram[100][0] ), 
	.D(n2182), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][15]  (.Q(\ram[96][15] ), 
	.D(n2133), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][14]  (.Q(\ram[96][14] ), 
	.D(n2132), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][13]  (.Q(\ram[96][13] ), 
	.D(n2131), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][12]  (.Q(\ram[96][12] ), 
	.D(n2130), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][11]  (.Q(\ram[96][11] ), 
	.D(n2129), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][10]  (.Q(\ram[96][10] ), 
	.D(n2128), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][9]  (.Q(\ram[96][9] ), 
	.D(n2127), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][8]  (.Q(\ram[96][8] ), 
	.D(n2126), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][7]  (.Q(\ram[96][7] ), 
	.D(n2125), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][6]  (.Q(\ram[96][6] ), 
	.D(n2124), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][5]  (.Q(\ram[96][5] ), 
	.D(n2123), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][4]  (.Q(\ram[96][4] ), 
	.D(n2122), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][3]  (.Q(\ram[96][3] ), 
	.D(n2121), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][2]  (.Q(\ram[96][2] ), 
	.D(n2120), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][1]  (.Q(\ram[96][1] ), 
	.D(n2119), 
	.CK(clk));
   DFFHQX1 \ram_reg[96][0]  (.Q(\ram[96][0] ), 
	.D(n2118), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][15]  (.Q(\ram[92][15] ), 
	.D(n2069), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][14]  (.Q(\ram[92][14] ), 
	.D(n2068), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][13]  (.Q(\ram[92][13] ), 
	.D(n2067), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][12]  (.Q(\ram[92][12] ), 
	.D(n2066), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][11]  (.Q(\ram[92][11] ), 
	.D(n2065), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][10]  (.Q(\ram[92][10] ), 
	.D(n2064), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][9]  (.Q(\ram[92][9] ), 
	.D(n2063), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][8]  (.Q(\ram[92][8] ), 
	.D(n2062), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][7]  (.Q(\ram[92][7] ), 
	.D(n2061), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][6]  (.Q(\ram[92][6] ), 
	.D(n2060), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][5]  (.Q(\ram[92][5] ), 
	.D(n2059), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][4]  (.Q(\ram[92][4] ), 
	.D(n2058), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][3]  (.Q(\ram[92][3] ), 
	.D(n2057), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][2]  (.Q(\ram[92][2] ), 
	.D(n2056), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][1]  (.Q(\ram[92][1] ), 
	.D(n2055), 
	.CK(clk));
   DFFHQX1 \ram_reg[92][0]  (.Q(\ram[92][0] ), 
	.D(n2054), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][15]  (.Q(\ram[88][15] ), 
	.D(n2005), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][14]  (.Q(\ram[88][14] ), 
	.D(n2004), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][13]  (.Q(\ram[88][13] ), 
	.D(n2003), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][12]  (.Q(\ram[88][12] ), 
	.D(n2002), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][11]  (.Q(\ram[88][11] ), 
	.D(n2001), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][10]  (.Q(\ram[88][10] ), 
	.D(n2000), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][9]  (.Q(\ram[88][9] ), 
	.D(n1999), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][8]  (.Q(\ram[88][8] ), 
	.D(n1998), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][7]  (.Q(\ram[88][7] ), 
	.D(n1997), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][6]  (.Q(\ram[88][6] ), 
	.D(n1996), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][5]  (.Q(\ram[88][5] ), 
	.D(n1995), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][4]  (.Q(\ram[88][4] ), 
	.D(n1994), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][3]  (.Q(\ram[88][3] ), 
	.D(n1993), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][2]  (.Q(\ram[88][2] ), 
	.D(n1992), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][1]  (.Q(\ram[88][1] ), 
	.D(n1991), 
	.CK(clk));
   DFFHQX1 \ram_reg[88][0]  (.Q(\ram[88][0] ), 
	.D(n1990), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][15]  (.Q(\ram[84][15] ), 
	.D(n1941), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][14]  (.Q(\ram[84][14] ), 
	.D(n1940), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][13]  (.Q(\ram[84][13] ), 
	.D(n1939), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][12]  (.Q(\ram[84][12] ), 
	.D(n1938), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][11]  (.Q(\ram[84][11] ), 
	.D(n1937), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][10]  (.Q(\ram[84][10] ), 
	.D(n1936), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][9]  (.Q(\ram[84][9] ), 
	.D(n1935), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][8]  (.Q(\ram[84][8] ), 
	.D(n1934), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][7]  (.Q(\ram[84][7] ), 
	.D(n1933), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][6]  (.Q(\ram[84][6] ), 
	.D(n1932), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][5]  (.Q(\ram[84][5] ), 
	.D(n1931), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][4]  (.Q(\ram[84][4] ), 
	.D(n1930), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][3]  (.Q(\ram[84][3] ), 
	.D(n1929), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][2]  (.Q(\ram[84][2] ), 
	.D(n1928), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][1]  (.Q(\ram[84][1] ), 
	.D(n1927), 
	.CK(clk));
   DFFHQX1 \ram_reg[84][0]  (.Q(\ram[84][0] ), 
	.D(n1926), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][15]  (.Q(\ram[80][15] ), 
	.D(n1877), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][14]  (.Q(\ram[80][14] ), 
	.D(n1876), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][13]  (.Q(\ram[80][13] ), 
	.D(n1875), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][12]  (.Q(\ram[80][12] ), 
	.D(n1874), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][11]  (.Q(\ram[80][11] ), 
	.D(n1873), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][10]  (.Q(\ram[80][10] ), 
	.D(n1872), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][9]  (.Q(\ram[80][9] ), 
	.D(n1871), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][8]  (.Q(\ram[80][8] ), 
	.D(n1870), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][7]  (.Q(\ram[80][7] ), 
	.D(n1869), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][6]  (.Q(\ram[80][6] ), 
	.D(n1868), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][5]  (.Q(\ram[80][5] ), 
	.D(n1867), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][4]  (.Q(\ram[80][4] ), 
	.D(n1866), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][3]  (.Q(\ram[80][3] ), 
	.D(n1865), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][2]  (.Q(\ram[80][2] ), 
	.D(n1864), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][1]  (.Q(\ram[80][1] ), 
	.D(n1863), 
	.CK(clk));
   DFFHQX1 \ram_reg[80][0]  (.Q(\ram[80][0] ), 
	.D(n1862), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][15]  (.Q(\ram[76][15] ), 
	.D(n1813), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][14]  (.Q(\ram[76][14] ), 
	.D(n1812), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][13]  (.Q(\ram[76][13] ), 
	.D(n1811), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][12]  (.Q(\ram[76][12] ), 
	.D(n1810), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][11]  (.Q(\ram[76][11] ), 
	.D(n1809), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][10]  (.Q(\ram[76][10] ), 
	.D(n1808), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][9]  (.Q(\ram[76][9] ), 
	.D(n1807), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][8]  (.Q(\ram[76][8] ), 
	.D(n1806), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][7]  (.Q(\ram[76][7] ), 
	.D(n1805), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][6]  (.Q(\ram[76][6] ), 
	.D(n1804), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][5]  (.Q(\ram[76][5] ), 
	.D(n1803), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][4]  (.Q(\ram[76][4] ), 
	.D(n1802), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][3]  (.Q(\ram[76][3] ), 
	.D(n1801), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][2]  (.Q(\ram[76][2] ), 
	.D(n1800), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][1]  (.Q(\ram[76][1] ), 
	.D(n1799), 
	.CK(clk));
   DFFHQX1 \ram_reg[76][0]  (.Q(\ram[76][0] ), 
	.D(n1798), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][15]  (.Q(\ram[72][15] ), 
	.D(n1749), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][14]  (.Q(\ram[72][14] ), 
	.D(n1748), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][13]  (.Q(\ram[72][13] ), 
	.D(n1747), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][12]  (.Q(\ram[72][12] ), 
	.D(n1746), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][11]  (.Q(\ram[72][11] ), 
	.D(n1745), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][10]  (.Q(\ram[72][10] ), 
	.D(n1744), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][9]  (.Q(\ram[72][9] ), 
	.D(n1743), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][8]  (.Q(\ram[72][8] ), 
	.D(n1742), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][7]  (.Q(\ram[72][7] ), 
	.D(n1741), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][6]  (.Q(\ram[72][6] ), 
	.D(n1740), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][5]  (.Q(\ram[72][5] ), 
	.D(n1739), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][4]  (.Q(\ram[72][4] ), 
	.D(n1738), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][3]  (.Q(\ram[72][3] ), 
	.D(n1737), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][2]  (.Q(\ram[72][2] ), 
	.D(n1736), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][1]  (.Q(\ram[72][1] ), 
	.D(n1735), 
	.CK(clk));
   DFFHQX1 \ram_reg[72][0]  (.Q(\ram[72][0] ), 
	.D(n1734), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][15]  (.Q(\ram[68][15] ), 
	.D(n1685), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][14]  (.Q(\ram[68][14] ), 
	.D(n1684), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][13]  (.Q(\ram[68][13] ), 
	.D(n1683), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][12]  (.Q(\ram[68][12] ), 
	.D(n1682), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][11]  (.Q(\ram[68][11] ), 
	.D(n1681), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][10]  (.Q(\ram[68][10] ), 
	.D(n1680), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][9]  (.Q(\ram[68][9] ), 
	.D(n1679), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][8]  (.Q(\ram[68][8] ), 
	.D(n1678), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][7]  (.Q(\ram[68][7] ), 
	.D(n1677), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][6]  (.Q(\ram[68][6] ), 
	.D(n1676), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][5]  (.Q(\ram[68][5] ), 
	.D(n1675), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][4]  (.Q(\ram[68][4] ), 
	.D(n1674), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][3]  (.Q(\ram[68][3] ), 
	.D(n1673), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][2]  (.Q(\ram[68][2] ), 
	.D(n1672), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][1]  (.Q(\ram[68][1] ), 
	.D(n1671), 
	.CK(clk));
   DFFHQX1 \ram_reg[68][0]  (.Q(\ram[68][0] ), 
	.D(n1670), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][15]  (.Q(\ram[64][15] ), 
	.D(n1621), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][14]  (.Q(\ram[64][14] ), 
	.D(n1620), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][13]  (.Q(\ram[64][13] ), 
	.D(n1619), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][12]  (.Q(\ram[64][12] ), 
	.D(n1618), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][11]  (.Q(\ram[64][11] ), 
	.D(n1617), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][10]  (.Q(\ram[64][10] ), 
	.D(n1616), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][9]  (.Q(\ram[64][9] ), 
	.D(n1615), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][8]  (.Q(\ram[64][8] ), 
	.D(n1614), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][7]  (.Q(\ram[64][7] ), 
	.D(n1613), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][6]  (.Q(\ram[64][6] ), 
	.D(n1612), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][5]  (.Q(\ram[64][5] ), 
	.D(n1611), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][4]  (.Q(\ram[64][4] ), 
	.D(n1610), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][3]  (.Q(\ram[64][3] ), 
	.D(n1609), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][2]  (.Q(\ram[64][2] ), 
	.D(n1608), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][1]  (.Q(\ram[64][1] ), 
	.D(n1607), 
	.CK(clk));
   DFFHQX1 \ram_reg[64][0]  (.Q(\ram[64][0] ), 
	.D(n1606), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][15]  (.Q(\ram[60][15] ), 
	.D(n1557), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][14]  (.Q(\ram[60][14] ), 
	.D(n1556), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][13]  (.Q(\ram[60][13] ), 
	.D(n1555), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][12]  (.Q(\ram[60][12] ), 
	.D(n1554), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][11]  (.Q(\ram[60][11] ), 
	.D(n1553), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][10]  (.Q(\ram[60][10] ), 
	.D(n1552), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][9]  (.Q(\ram[60][9] ), 
	.D(n1551), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][8]  (.Q(\ram[60][8] ), 
	.D(n1550), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][7]  (.Q(\ram[60][7] ), 
	.D(n1549), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][6]  (.Q(\ram[60][6] ), 
	.D(n1548), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][5]  (.Q(\ram[60][5] ), 
	.D(n1547), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][4]  (.Q(\ram[60][4] ), 
	.D(n1546), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][3]  (.Q(\ram[60][3] ), 
	.D(n1545), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][2]  (.Q(\ram[60][2] ), 
	.D(n1544), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][1]  (.Q(\ram[60][1] ), 
	.D(n1543), 
	.CK(clk));
   DFFHQX1 \ram_reg[60][0]  (.Q(\ram[60][0] ), 
	.D(n1542), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][15]  (.Q(\ram[56][15] ), 
	.D(n1493), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][14]  (.Q(\ram[56][14] ), 
	.D(n1492), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][13]  (.Q(\ram[56][13] ), 
	.D(n1491), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][12]  (.Q(\ram[56][12] ), 
	.D(n1490), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][11]  (.Q(\ram[56][11] ), 
	.D(n1489), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][10]  (.Q(\ram[56][10] ), 
	.D(n1488), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][9]  (.Q(\ram[56][9] ), 
	.D(n1487), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][8]  (.Q(\ram[56][8] ), 
	.D(n1486), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][7]  (.Q(\ram[56][7] ), 
	.D(n1485), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][6]  (.Q(\ram[56][6] ), 
	.D(n1484), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][5]  (.Q(\ram[56][5] ), 
	.D(n1483), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][4]  (.Q(\ram[56][4] ), 
	.D(n1482), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][3]  (.Q(\ram[56][3] ), 
	.D(n1481), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][2]  (.Q(\ram[56][2] ), 
	.D(n1480), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][1]  (.Q(\ram[56][1] ), 
	.D(n1479), 
	.CK(clk));
   DFFHQX1 \ram_reg[56][0]  (.Q(\ram[56][0] ), 
	.D(n1478), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][15]  (.Q(\ram[52][15] ), 
	.D(n1429), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][14]  (.Q(\ram[52][14] ), 
	.D(n1428), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][13]  (.Q(\ram[52][13] ), 
	.D(n1427), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][12]  (.Q(\ram[52][12] ), 
	.D(n1426), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][11]  (.Q(\ram[52][11] ), 
	.D(n1425), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][10]  (.Q(\ram[52][10] ), 
	.D(n1424), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][9]  (.Q(\ram[52][9] ), 
	.D(n1423), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][8]  (.Q(\ram[52][8] ), 
	.D(n1422), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][7]  (.Q(\ram[52][7] ), 
	.D(n1421), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][6]  (.Q(\ram[52][6] ), 
	.D(n1420), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][5]  (.Q(\ram[52][5] ), 
	.D(n1419), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][4]  (.Q(\ram[52][4] ), 
	.D(n1418), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][3]  (.Q(\ram[52][3] ), 
	.D(n1417), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][2]  (.Q(\ram[52][2] ), 
	.D(n1416), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][1]  (.Q(\ram[52][1] ), 
	.D(n1415), 
	.CK(clk));
   DFFHQX1 \ram_reg[52][0]  (.Q(\ram[52][0] ), 
	.D(n1414), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][15]  (.Q(\ram[48][15] ), 
	.D(n1365), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][14]  (.Q(\ram[48][14] ), 
	.D(n1364), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][13]  (.Q(\ram[48][13] ), 
	.D(n1363), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][12]  (.Q(\ram[48][12] ), 
	.D(n1362), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][11]  (.Q(\ram[48][11] ), 
	.D(n1361), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][10]  (.Q(\ram[48][10] ), 
	.D(n1360), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][9]  (.Q(\ram[48][9] ), 
	.D(n1359), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][8]  (.Q(\ram[48][8] ), 
	.D(n1358), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][7]  (.Q(\ram[48][7] ), 
	.D(n1357), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][6]  (.Q(\ram[48][6] ), 
	.D(n1356), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][5]  (.Q(\ram[48][5] ), 
	.D(n1355), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][4]  (.Q(\ram[48][4] ), 
	.D(n1354), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][3]  (.Q(\ram[48][3] ), 
	.D(n1353), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][2]  (.Q(\ram[48][2] ), 
	.D(n1352), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][1]  (.Q(\ram[48][1] ), 
	.D(n1351), 
	.CK(clk));
   DFFHQX1 \ram_reg[48][0]  (.Q(\ram[48][0] ), 
	.D(n1350), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][15]  (.Q(\ram[44][15] ), 
	.D(n1301), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][14]  (.Q(\ram[44][14] ), 
	.D(n1300), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][13]  (.Q(\ram[44][13] ), 
	.D(n1299), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][12]  (.Q(\ram[44][12] ), 
	.D(n1298), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][11]  (.Q(\ram[44][11] ), 
	.D(n1297), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][10]  (.Q(\ram[44][10] ), 
	.D(n1296), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][9]  (.Q(\ram[44][9] ), 
	.D(n1295), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][8]  (.Q(\ram[44][8] ), 
	.D(n1294), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][7]  (.Q(\ram[44][7] ), 
	.D(n1293), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][6]  (.Q(\ram[44][6] ), 
	.D(n1292), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][5]  (.Q(\ram[44][5] ), 
	.D(n1291), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][4]  (.Q(\ram[44][4] ), 
	.D(n1290), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][3]  (.Q(\ram[44][3] ), 
	.D(n1289), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][2]  (.Q(\ram[44][2] ), 
	.D(n1288), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][1]  (.Q(\ram[44][1] ), 
	.D(n1287), 
	.CK(clk));
   DFFHQX1 \ram_reg[44][0]  (.Q(\ram[44][0] ), 
	.D(n1286), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][15]  (.Q(\ram[40][15] ), 
	.D(n1237), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][14]  (.Q(\ram[40][14] ), 
	.D(n1236), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][13]  (.Q(\ram[40][13] ), 
	.D(n1235), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][12]  (.Q(\ram[40][12] ), 
	.D(n1234), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][11]  (.Q(\ram[40][11] ), 
	.D(n1233), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][10]  (.Q(\ram[40][10] ), 
	.D(n1232), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][9]  (.Q(\ram[40][9] ), 
	.D(n1231), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][8]  (.Q(\ram[40][8] ), 
	.D(n1230), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][7]  (.Q(\ram[40][7] ), 
	.D(n1229), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][6]  (.Q(\ram[40][6] ), 
	.D(n1228), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][5]  (.Q(\ram[40][5] ), 
	.D(n1227), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][4]  (.Q(\ram[40][4] ), 
	.D(n1226), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][3]  (.Q(\ram[40][3] ), 
	.D(n1225), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][2]  (.Q(\ram[40][2] ), 
	.D(n1224), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][1]  (.Q(\ram[40][1] ), 
	.D(n1223), 
	.CK(clk));
   DFFHQX1 \ram_reg[40][0]  (.Q(\ram[40][0] ), 
	.D(n1222), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][15]  (.Q(\ram[36][15] ), 
	.D(n1173), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][14]  (.Q(\ram[36][14] ), 
	.D(n1172), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][13]  (.Q(\ram[36][13] ), 
	.D(n1171), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][12]  (.Q(\ram[36][12] ), 
	.D(n1170), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][11]  (.Q(\ram[36][11] ), 
	.D(n1169), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][10]  (.Q(\ram[36][10] ), 
	.D(n1168), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][9]  (.Q(\ram[36][9] ), 
	.D(n1167), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][8]  (.Q(\ram[36][8] ), 
	.D(n1166), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][7]  (.Q(\ram[36][7] ), 
	.D(n1165), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][6]  (.Q(\ram[36][6] ), 
	.D(n1164), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][5]  (.Q(\ram[36][5] ), 
	.D(n1163), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][4]  (.Q(\ram[36][4] ), 
	.D(n1162), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][3]  (.Q(\ram[36][3] ), 
	.D(n1161), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][2]  (.Q(\ram[36][2] ), 
	.D(n1160), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][1]  (.Q(\ram[36][1] ), 
	.D(n1159), 
	.CK(clk));
   DFFHQX1 \ram_reg[36][0]  (.Q(\ram[36][0] ), 
	.D(n1158), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][15]  (.Q(\ram[32][15] ), 
	.D(n1109), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][14]  (.Q(\ram[32][14] ), 
	.D(n1108), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][13]  (.Q(\ram[32][13] ), 
	.D(n1107), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][12]  (.Q(\ram[32][12] ), 
	.D(n1106), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][11]  (.Q(\ram[32][11] ), 
	.D(n1105), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][10]  (.Q(\ram[32][10] ), 
	.D(n1104), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][9]  (.Q(\ram[32][9] ), 
	.D(n1103), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][8]  (.Q(\ram[32][8] ), 
	.D(n1102), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][7]  (.Q(\ram[32][7] ), 
	.D(n1101), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][6]  (.Q(\ram[32][6] ), 
	.D(n1100), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][5]  (.Q(\ram[32][5] ), 
	.D(n1099), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][4]  (.Q(\ram[32][4] ), 
	.D(n1098), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][3]  (.Q(\ram[32][3] ), 
	.D(n1097), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][2]  (.Q(\ram[32][2] ), 
	.D(n1096), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][1]  (.Q(\ram[32][1] ), 
	.D(n1095), 
	.CK(clk));
   DFFHQX1 \ram_reg[32][0]  (.Q(\ram[32][0] ), 
	.D(n1094), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][15]  (.Q(\ram[28][15] ), 
	.D(n1045), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][14]  (.Q(\ram[28][14] ), 
	.D(n1044), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][13]  (.Q(\ram[28][13] ), 
	.D(n1043), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][12]  (.Q(\ram[28][12] ), 
	.D(n1042), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][11]  (.Q(\ram[28][11] ), 
	.D(n1041), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][10]  (.Q(\ram[28][10] ), 
	.D(n1040), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][9]  (.Q(\ram[28][9] ), 
	.D(n1039), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][8]  (.Q(\ram[28][8] ), 
	.D(n1038), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][7]  (.Q(\ram[28][7] ), 
	.D(n1037), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][6]  (.Q(\ram[28][6] ), 
	.D(n1036), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][5]  (.Q(\ram[28][5] ), 
	.D(n1035), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][4]  (.Q(\ram[28][4] ), 
	.D(n1034), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][3]  (.Q(\ram[28][3] ), 
	.D(n1033), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][2]  (.Q(\ram[28][2] ), 
	.D(n1032), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][1]  (.Q(\ram[28][1] ), 
	.D(n1031), 
	.CK(clk));
   DFFHQX1 \ram_reg[28][0]  (.Q(\ram[28][0] ), 
	.D(n1030), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][15]  (.Q(\ram[24][15] ), 
	.D(n981), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][14]  (.Q(\ram[24][14] ), 
	.D(n980), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][13]  (.Q(\ram[24][13] ), 
	.D(n979), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][12]  (.Q(\ram[24][12] ), 
	.D(n978), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][11]  (.Q(\ram[24][11] ), 
	.D(n977), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][10]  (.Q(\ram[24][10] ), 
	.D(n976), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][9]  (.Q(\ram[24][9] ), 
	.D(n975), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][8]  (.Q(\ram[24][8] ), 
	.D(n974), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][7]  (.Q(\ram[24][7] ), 
	.D(n973), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][6]  (.Q(\ram[24][6] ), 
	.D(n972), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][5]  (.Q(\ram[24][5] ), 
	.D(n971), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][4]  (.Q(\ram[24][4] ), 
	.D(n970), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][3]  (.Q(\ram[24][3] ), 
	.D(n969), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][2]  (.Q(\ram[24][2] ), 
	.D(n968), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][1]  (.Q(\ram[24][1] ), 
	.D(n967), 
	.CK(clk));
   DFFHQX1 \ram_reg[24][0]  (.Q(\ram[24][0] ), 
	.D(n966), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][15]  (.Q(\ram[20][15] ), 
	.D(n917), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][14]  (.Q(\ram[20][14] ), 
	.D(n916), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][13]  (.Q(\ram[20][13] ), 
	.D(n915), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][12]  (.Q(\ram[20][12] ), 
	.D(n914), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][11]  (.Q(\ram[20][11] ), 
	.D(n913), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][10]  (.Q(\ram[20][10] ), 
	.D(n912), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][9]  (.Q(\ram[20][9] ), 
	.D(n911), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][8]  (.Q(\ram[20][8] ), 
	.D(n910), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][7]  (.Q(\ram[20][7] ), 
	.D(n909), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][6]  (.Q(\ram[20][6] ), 
	.D(n908), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][5]  (.Q(\ram[20][5] ), 
	.D(n907), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][4]  (.Q(\ram[20][4] ), 
	.D(n906), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][3]  (.Q(\ram[20][3] ), 
	.D(n905), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][2]  (.Q(\ram[20][2] ), 
	.D(n904), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][1]  (.Q(\ram[20][1] ), 
	.D(n903), 
	.CK(clk));
   DFFHQX1 \ram_reg[20][0]  (.Q(\ram[20][0] ), 
	.D(n902), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][15]  (.Q(\ram[16][15] ), 
	.D(n853), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][14]  (.Q(\ram[16][14] ), 
	.D(n852), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][13]  (.Q(\ram[16][13] ), 
	.D(n851), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][12]  (.Q(\ram[16][12] ), 
	.D(n850), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][11]  (.Q(\ram[16][11] ), 
	.D(n849), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][10]  (.Q(\ram[16][10] ), 
	.D(n848), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][9]  (.Q(\ram[16][9] ), 
	.D(n847), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][8]  (.Q(\ram[16][8] ), 
	.D(n846), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][7]  (.Q(\ram[16][7] ), 
	.D(n845), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][6]  (.Q(\ram[16][6] ), 
	.D(n844), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][5]  (.Q(\ram[16][5] ), 
	.D(n843), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][4]  (.Q(\ram[16][4] ), 
	.D(n842), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][3]  (.Q(\ram[16][3] ), 
	.D(n841), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][2]  (.Q(\ram[16][2] ), 
	.D(n840), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][1]  (.Q(\ram[16][1] ), 
	.D(n839), 
	.CK(clk));
   DFFHQX1 \ram_reg[16][0]  (.Q(\ram[16][0] ), 
	.D(n838), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][15]  (.Q(\ram[12][15] ), 
	.D(n789), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][14]  (.Q(\ram[12][14] ), 
	.D(n788), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][13]  (.Q(\ram[12][13] ), 
	.D(n787), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][12]  (.Q(\ram[12][12] ), 
	.D(n786), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][11]  (.Q(\ram[12][11] ), 
	.D(n785), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][10]  (.Q(\ram[12][10] ), 
	.D(n784), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][9]  (.Q(\ram[12][9] ), 
	.D(n783), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][8]  (.Q(\ram[12][8] ), 
	.D(n782), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][7]  (.Q(\ram[12][7] ), 
	.D(n781), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][6]  (.Q(\ram[12][6] ), 
	.D(n780), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][5]  (.Q(\ram[12][5] ), 
	.D(n779), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][4]  (.Q(\ram[12][4] ), 
	.D(n778), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][3]  (.Q(\ram[12][3] ), 
	.D(n777), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][2]  (.Q(\ram[12][2] ), 
	.D(n776), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][1]  (.Q(\ram[12][1] ), 
	.D(n775), 
	.CK(clk));
   DFFHQX1 \ram_reg[12][0]  (.Q(\ram[12][0] ), 
	.D(n774), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][15]  (.Q(\ram[8][15] ), 
	.D(n725), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][14]  (.Q(\ram[8][14] ), 
	.D(n724), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][13]  (.Q(\ram[8][13] ), 
	.D(n723), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][12]  (.Q(\ram[8][12] ), 
	.D(n722), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][11]  (.Q(\ram[8][11] ), 
	.D(n721), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][10]  (.Q(\ram[8][10] ), 
	.D(n720), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][9]  (.Q(\ram[8][9] ), 
	.D(n719), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][8]  (.Q(\ram[8][8] ), 
	.D(n718), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][7]  (.Q(\ram[8][7] ), 
	.D(n717), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][6]  (.Q(\ram[8][6] ), 
	.D(n716), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][5]  (.Q(\ram[8][5] ), 
	.D(n715), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][4]  (.Q(\ram[8][4] ), 
	.D(n714), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][3]  (.Q(\ram[8][3] ), 
	.D(n713), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][2]  (.Q(\ram[8][2] ), 
	.D(n712), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][1]  (.Q(\ram[8][1] ), 
	.D(n711), 
	.CK(clk));
   DFFHQX1 \ram_reg[8][0]  (.Q(\ram[8][0] ), 
	.D(n710), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][15]  (.Q(\ram[4][15] ), 
	.D(n661), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][14]  (.Q(\ram[4][14] ), 
	.D(n660), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][13]  (.Q(\ram[4][13] ), 
	.D(n659), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][12]  (.Q(\ram[4][12] ), 
	.D(n658), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][11]  (.Q(\ram[4][11] ), 
	.D(n657), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][10]  (.Q(\ram[4][10] ), 
	.D(n656), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][9]  (.Q(\ram[4][9] ), 
	.D(n655), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][8]  (.Q(\ram[4][8] ), 
	.D(n654), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][7]  (.Q(\ram[4][7] ), 
	.D(n653), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][6]  (.Q(\ram[4][6] ), 
	.D(n652), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][5]  (.Q(\ram[4][5] ), 
	.D(n651), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][4]  (.Q(\ram[4][4] ), 
	.D(n650), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][3]  (.Q(\ram[4][3] ), 
	.D(n649), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][2]  (.Q(\ram[4][2] ), 
	.D(n648), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][1]  (.Q(\ram[4][1] ), 
	.D(n647), 
	.CK(clk));
   DFFHQX1 \ram_reg[4][0]  (.Q(\ram[4][0] ), 
	.D(n646), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][15]  (.Q(\ram[0][15] ), 
	.D(n597), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][14]  (.Q(\ram[0][14] ), 
	.D(n596), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][13]  (.Q(\ram[0][13] ), 
	.D(n595), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][12]  (.Q(\ram[0][12] ), 
	.D(n594), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][11]  (.Q(\ram[0][11] ), 
	.D(n593), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][10]  (.Q(\ram[0][10] ), 
	.D(n592), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][9]  (.Q(\ram[0][9] ), 
	.D(n591), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][8]  (.Q(\ram[0][8] ), 
	.D(n590), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][7]  (.Q(\ram[0][7] ), 
	.D(n589), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][6]  (.Q(\ram[0][6] ), 
	.D(n588), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][5]  (.Q(\ram[0][5] ), 
	.D(n587), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][4]  (.Q(\ram[0][4] ), 
	.D(n586), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][3]  (.Q(\ram[0][3] ), 
	.D(n585), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][2]  (.Q(\ram[0][2] ), 
	.D(n584), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][1]  (.Q(\ram[0][1] ), 
	.D(n583), 
	.CK(clk));
   DFFHQX1 \ram_reg[0][0]  (.Q(\ram[0][0] ), 
	.D(n582), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][15]  (.Q(\ram[254][15] ), 
	.D(n4661), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][14]  (.Q(\ram[254][14] ), 
	.D(n4660), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][13]  (.Q(\ram[254][13] ), 
	.D(n4659), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][12]  (.Q(\ram[254][12] ), 
	.D(n4658), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][11]  (.Q(\ram[254][11] ), 
	.D(n4657), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][10]  (.Q(\ram[254][10] ), 
	.D(n4656), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][9]  (.Q(\ram[254][9] ), 
	.D(n4655), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][8]  (.Q(\ram[254][8] ), 
	.D(n4654), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][7]  (.Q(\ram[254][7] ), 
	.D(n4653), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][6]  (.Q(\ram[254][6] ), 
	.D(n4652), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][5]  (.Q(\ram[254][5] ), 
	.D(n4651), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][4]  (.Q(\ram[254][4] ), 
	.D(n4650), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][3]  (.Q(\ram[254][3] ), 
	.D(n4649), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][2]  (.Q(\ram[254][2] ), 
	.D(n4648), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][1]  (.Q(\ram[254][1] ), 
	.D(n4647), 
	.CK(clk));
   DFFHQX1 \ram_reg[254][0]  (.Q(\ram[254][0] ), 
	.D(n4646), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][15]  (.Q(\ram[250][15] ), 
	.D(n4597), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][14]  (.Q(\ram[250][14] ), 
	.D(n4596), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][13]  (.Q(\ram[250][13] ), 
	.D(n4595), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][12]  (.Q(\ram[250][12] ), 
	.D(n4594), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][11]  (.Q(\ram[250][11] ), 
	.D(n4593), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][10]  (.Q(\ram[250][10] ), 
	.D(n4592), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][9]  (.Q(\ram[250][9] ), 
	.D(n4591), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][8]  (.Q(\ram[250][8] ), 
	.D(n4590), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][7]  (.Q(\ram[250][7] ), 
	.D(n4589), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][6]  (.Q(\ram[250][6] ), 
	.D(n4588), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][5]  (.Q(\ram[250][5] ), 
	.D(n4587), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][4]  (.Q(\ram[250][4] ), 
	.D(n4586), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][3]  (.Q(\ram[250][3] ), 
	.D(n4585), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][2]  (.Q(\ram[250][2] ), 
	.D(n4584), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][1]  (.Q(\ram[250][1] ), 
	.D(n4583), 
	.CK(clk));
   DFFHQX1 \ram_reg[250][0]  (.Q(\ram[250][0] ), 
	.D(n4582), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][15]  (.Q(\ram[246][15] ), 
	.D(n4533), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][14]  (.Q(\ram[246][14] ), 
	.D(n4532), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][13]  (.Q(\ram[246][13] ), 
	.D(n4531), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][12]  (.Q(\ram[246][12] ), 
	.D(n4530), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][11]  (.Q(\ram[246][11] ), 
	.D(n4529), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][10]  (.Q(\ram[246][10] ), 
	.D(n4528), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][9]  (.Q(\ram[246][9] ), 
	.D(n4527), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][8]  (.Q(\ram[246][8] ), 
	.D(n4526), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][7]  (.Q(\ram[246][7] ), 
	.D(n4525), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][6]  (.Q(\ram[246][6] ), 
	.D(n4524), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][5]  (.Q(\ram[246][5] ), 
	.D(n4523), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][4]  (.Q(\ram[246][4] ), 
	.D(n4522), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][3]  (.Q(\ram[246][3] ), 
	.D(n4521), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][2]  (.Q(\ram[246][2] ), 
	.D(n4520), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][1]  (.Q(\ram[246][1] ), 
	.D(n4519), 
	.CK(clk));
   DFFHQX1 \ram_reg[246][0]  (.Q(\ram[246][0] ), 
	.D(n4518), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][15]  (.Q(\ram[242][15] ), 
	.D(n4469), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][14]  (.Q(\ram[242][14] ), 
	.D(n4468), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][13]  (.Q(\ram[242][13] ), 
	.D(n4467), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][12]  (.Q(\ram[242][12] ), 
	.D(n4466), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][11]  (.Q(\ram[242][11] ), 
	.D(n4465), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][10]  (.Q(\ram[242][10] ), 
	.D(n4464), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][9]  (.Q(\ram[242][9] ), 
	.D(n4463), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][8]  (.Q(\ram[242][8] ), 
	.D(n4462), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][7]  (.Q(\ram[242][7] ), 
	.D(n4461), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][6]  (.Q(\ram[242][6] ), 
	.D(n4460), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][5]  (.Q(\ram[242][5] ), 
	.D(n4459), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][4]  (.Q(\ram[242][4] ), 
	.D(n4458), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][3]  (.Q(\ram[242][3] ), 
	.D(n4457), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][2]  (.Q(\ram[242][2] ), 
	.D(n4456), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][1]  (.Q(\ram[242][1] ), 
	.D(n4455), 
	.CK(clk));
   DFFHQX1 \ram_reg[242][0]  (.Q(\ram[242][0] ), 
	.D(n4454), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][15]  (.Q(\ram[238][15] ), 
	.D(n4405), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][14]  (.Q(\ram[238][14] ), 
	.D(n4404), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][13]  (.Q(\ram[238][13] ), 
	.D(n4403), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][12]  (.Q(\ram[238][12] ), 
	.D(n4402), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][11]  (.Q(\ram[238][11] ), 
	.D(n4401), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][10]  (.Q(\ram[238][10] ), 
	.D(n4400), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][9]  (.Q(\ram[238][9] ), 
	.D(n4399), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][8]  (.Q(\ram[238][8] ), 
	.D(n4398), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][7]  (.Q(\ram[238][7] ), 
	.D(n4397), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][6]  (.Q(\ram[238][6] ), 
	.D(n4396), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][5]  (.Q(\ram[238][5] ), 
	.D(n4395), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][4]  (.Q(\ram[238][4] ), 
	.D(n4394), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][3]  (.Q(\ram[238][3] ), 
	.D(n4393), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][2]  (.Q(\ram[238][2] ), 
	.D(n4392), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][1]  (.Q(\ram[238][1] ), 
	.D(n4391), 
	.CK(clk));
   DFFHQX1 \ram_reg[238][0]  (.Q(\ram[238][0] ), 
	.D(n4390), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][15]  (.Q(\ram[234][15] ), 
	.D(n4341), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][14]  (.Q(\ram[234][14] ), 
	.D(n4340), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][13]  (.Q(\ram[234][13] ), 
	.D(n4339), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][12]  (.Q(\ram[234][12] ), 
	.D(n4338), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][11]  (.Q(\ram[234][11] ), 
	.D(n4337), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][10]  (.Q(\ram[234][10] ), 
	.D(n4336), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][9]  (.Q(\ram[234][9] ), 
	.D(n4335), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][8]  (.Q(\ram[234][8] ), 
	.D(n4334), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][7]  (.Q(\ram[234][7] ), 
	.D(n4333), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][6]  (.Q(\ram[234][6] ), 
	.D(n4332), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][5]  (.Q(\ram[234][5] ), 
	.D(n4331), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][4]  (.Q(\ram[234][4] ), 
	.D(n4330), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][3]  (.Q(\ram[234][3] ), 
	.D(n4329), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][2]  (.Q(\ram[234][2] ), 
	.D(n4328), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][1]  (.Q(\ram[234][1] ), 
	.D(n4327), 
	.CK(clk));
   DFFHQX1 \ram_reg[234][0]  (.Q(\ram[234][0] ), 
	.D(n4326), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][15]  (.Q(\ram[230][15] ), 
	.D(n4277), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][14]  (.Q(\ram[230][14] ), 
	.D(n4276), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][13]  (.Q(\ram[230][13] ), 
	.D(n4275), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][12]  (.Q(\ram[230][12] ), 
	.D(n4274), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][11]  (.Q(\ram[230][11] ), 
	.D(n4273), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][10]  (.Q(\ram[230][10] ), 
	.D(n4272), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][9]  (.Q(\ram[230][9] ), 
	.D(n4271), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][8]  (.Q(\ram[230][8] ), 
	.D(n4270), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][7]  (.Q(\ram[230][7] ), 
	.D(n4269), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][6]  (.Q(\ram[230][6] ), 
	.D(n4268), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][5]  (.Q(\ram[230][5] ), 
	.D(n4267), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][4]  (.Q(\ram[230][4] ), 
	.D(n4266), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][3]  (.Q(\ram[230][3] ), 
	.D(n4265), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][2]  (.Q(\ram[230][2] ), 
	.D(n4264), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][1]  (.Q(\ram[230][1] ), 
	.D(n4263), 
	.CK(clk));
   DFFHQX1 \ram_reg[230][0]  (.Q(\ram[230][0] ), 
	.D(n4262), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][15]  (.Q(\ram[226][15] ), 
	.D(n4213), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][14]  (.Q(\ram[226][14] ), 
	.D(n4212), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][13]  (.Q(\ram[226][13] ), 
	.D(n4211), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][12]  (.Q(\ram[226][12] ), 
	.D(n4210), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][11]  (.Q(\ram[226][11] ), 
	.D(n4209), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][10]  (.Q(\ram[226][10] ), 
	.D(n4208), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][9]  (.Q(\ram[226][9] ), 
	.D(n4207), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][8]  (.Q(\ram[226][8] ), 
	.D(n4206), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][7]  (.Q(\ram[226][7] ), 
	.D(n4205), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][6]  (.Q(\ram[226][6] ), 
	.D(n4204), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][5]  (.Q(\ram[226][5] ), 
	.D(n4203), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][4]  (.Q(\ram[226][4] ), 
	.D(n4202), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][3]  (.Q(\ram[226][3] ), 
	.D(n4201), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][2]  (.Q(\ram[226][2] ), 
	.D(n4200), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][1]  (.Q(\ram[226][1] ), 
	.D(n4199), 
	.CK(clk));
   DFFHQX1 \ram_reg[226][0]  (.Q(\ram[226][0] ), 
	.D(n4198), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][15]  (.Q(\ram[222][15] ), 
	.D(n4149), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][14]  (.Q(\ram[222][14] ), 
	.D(n4148), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][13]  (.Q(\ram[222][13] ), 
	.D(n4147), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][12]  (.Q(\ram[222][12] ), 
	.D(n4146), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][11]  (.Q(\ram[222][11] ), 
	.D(n4145), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][10]  (.Q(\ram[222][10] ), 
	.D(n4144), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][9]  (.Q(\ram[222][9] ), 
	.D(n4143), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][8]  (.Q(\ram[222][8] ), 
	.D(n4142), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][7]  (.Q(\ram[222][7] ), 
	.D(n4141), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][6]  (.Q(\ram[222][6] ), 
	.D(n4140), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][5]  (.Q(\ram[222][5] ), 
	.D(n4139), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][4]  (.Q(\ram[222][4] ), 
	.D(n4138), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][3]  (.Q(\ram[222][3] ), 
	.D(n4137), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][2]  (.Q(\ram[222][2] ), 
	.D(n4136), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][1]  (.Q(\ram[222][1] ), 
	.D(n4135), 
	.CK(clk));
   DFFHQX1 \ram_reg[222][0]  (.Q(\ram[222][0] ), 
	.D(n4134), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][15]  (.Q(\ram[218][15] ), 
	.D(n4085), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][14]  (.Q(\ram[218][14] ), 
	.D(n4084), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][13]  (.Q(\ram[218][13] ), 
	.D(n4083), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][12]  (.Q(\ram[218][12] ), 
	.D(n4082), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][11]  (.Q(\ram[218][11] ), 
	.D(n4081), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][10]  (.Q(\ram[218][10] ), 
	.D(n4080), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][9]  (.Q(\ram[218][9] ), 
	.D(n4079), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][8]  (.Q(\ram[218][8] ), 
	.D(n4078), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][7]  (.Q(\ram[218][7] ), 
	.D(n4077), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][6]  (.Q(\ram[218][6] ), 
	.D(n4076), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][5]  (.Q(\ram[218][5] ), 
	.D(n4075), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][4]  (.Q(\ram[218][4] ), 
	.D(n4074), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][3]  (.Q(\ram[218][3] ), 
	.D(n4073), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][2]  (.Q(\ram[218][2] ), 
	.D(n4072), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][1]  (.Q(\ram[218][1] ), 
	.D(n4071), 
	.CK(clk));
   DFFHQX1 \ram_reg[218][0]  (.Q(\ram[218][0] ), 
	.D(n4070), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][15]  (.Q(\ram[214][15] ), 
	.D(n4021), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][14]  (.Q(\ram[214][14] ), 
	.D(n4020), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][13]  (.Q(\ram[214][13] ), 
	.D(n4019), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][12]  (.Q(\ram[214][12] ), 
	.D(n4018), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][11]  (.Q(\ram[214][11] ), 
	.D(n4017), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][10]  (.Q(\ram[214][10] ), 
	.D(n4016), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][9]  (.Q(\ram[214][9] ), 
	.D(n4015), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][8]  (.Q(\ram[214][8] ), 
	.D(n4014), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][7]  (.Q(\ram[214][7] ), 
	.D(n4013), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][6]  (.Q(\ram[214][6] ), 
	.D(n4012), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][5]  (.Q(\ram[214][5] ), 
	.D(n4011), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][4]  (.Q(\ram[214][4] ), 
	.D(n4010), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][3]  (.Q(\ram[214][3] ), 
	.D(n4009), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][2]  (.Q(\ram[214][2] ), 
	.D(n4008), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][1]  (.Q(\ram[214][1] ), 
	.D(n4007), 
	.CK(clk));
   DFFHQX1 \ram_reg[214][0]  (.Q(\ram[214][0] ), 
	.D(n4006), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][15]  (.Q(\ram[210][15] ), 
	.D(n3957), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][14]  (.Q(\ram[210][14] ), 
	.D(n3956), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][13]  (.Q(\ram[210][13] ), 
	.D(n3955), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][12]  (.Q(\ram[210][12] ), 
	.D(n3954), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][11]  (.Q(\ram[210][11] ), 
	.D(n3953), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][10]  (.Q(\ram[210][10] ), 
	.D(n3952), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][9]  (.Q(\ram[210][9] ), 
	.D(n3951), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][8]  (.Q(\ram[210][8] ), 
	.D(n3950), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][7]  (.Q(\ram[210][7] ), 
	.D(n3949), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][6]  (.Q(\ram[210][6] ), 
	.D(n3948), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][5]  (.Q(\ram[210][5] ), 
	.D(n3947), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][4]  (.Q(\ram[210][4] ), 
	.D(n3946), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][3]  (.Q(\ram[210][3] ), 
	.D(n3945), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][2]  (.Q(\ram[210][2] ), 
	.D(n3944), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][1]  (.Q(\ram[210][1] ), 
	.D(n3943), 
	.CK(clk));
   DFFHQX1 \ram_reg[210][0]  (.Q(\ram[210][0] ), 
	.D(n3942), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][15]  (.Q(\ram[206][15] ), 
	.D(n3893), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][14]  (.Q(\ram[206][14] ), 
	.D(n3892), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][13]  (.Q(\ram[206][13] ), 
	.D(n3891), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][12]  (.Q(\ram[206][12] ), 
	.D(n3890), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][11]  (.Q(\ram[206][11] ), 
	.D(n3889), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][10]  (.Q(\ram[206][10] ), 
	.D(n3888), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][9]  (.Q(\ram[206][9] ), 
	.D(n3887), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][8]  (.Q(\ram[206][8] ), 
	.D(n3886), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][7]  (.Q(\ram[206][7] ), 
	.D(n3885), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][6]  (.Q(\ram[206][6] ), 
	.D(n3884), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][5]  (.Q(\ram[206][5] ), 
	.D(n3883), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][4]  (.Q(\ram[206][4] ), 
	.D(n3882), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][3]  (.Q(\ram[206][3] ), 
	.D(n3881), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][2]  (.Q(\ram[206][2] ), 
	.D(n3880), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][1]  (.Q(\ram[206][1] ), 
	.D(n3879), 
	.CK(clk));
   DFFHQX1 \ram_reg[206][0]  (.Q(\ram[206][0] ), 
	.D(n3878), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][15]  (.Q(\ram[202][15] ), 
	.D(n3829), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][14]  (.Q(\ram[202][14] ), 
	.D(n3828), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][13]  (.Q(\ram[202][13] ), 
	.D(n3827), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][12]  (.Q(\ram[202][12] ), 
	.D(n3826), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][11]  (.Q(\ram[202][11] ), 
	.D(n3825), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][10]  (.Q(\ram[202][10] ), 
	.D(n3824), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][9]  (.Q(\ram[202][9] ), 
	.D(n3823), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][8]  (.Q(\ram[202][8] ), 
	.D(n3822), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][7]  (.Q(\ram[202][7] ), 
	.D(n3821), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][6]  (.Q(\ram[202][6] ), 
	.D(n3820), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][5]  (.Q(\ram[202][5] ), 
	.D(n3819), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][4]  (.Q(\ram[202][4] ), 
	.D(n3818), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][3]  (.Q(\ram[202][3] ), 
	.D(n3817), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][2]  (.Q(\ram[202][2] ), 
	.D(n3816), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][1]  (.Q(\ram[202][1] ), 
	.D(n3815), 
	.CK(clk));
   DFFHQX1 \ram_reg[202][0]  (.Q(\ram[202][0] ), 
	.D(n3814), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][15]  (.Q(\ram[198][15] ), 
	.D(n3765), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][14]  (.Q(\ram[198][14] ), 
	.D(n3764), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][13]  (.Q(\ram[198][13] ), 
	.D(n3763), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][12]  (.Q(\ram[198][12] ), 
	.D(n3762), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][11]  (.Q(\ram[198][11] ), 
	.D(n3761), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][10]  (.Q(\ram[198][10] ), 
	.D(n3760), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][9]  (.Q(\ram[198][9] ), 
	.D(n3759), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][8]  (.Q(\ram[198][8] ), 
	.D(n3758), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][7]  (.Q(\ram[198][7] ), 
	.D(n3757), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][6]  (.Q(\ram[198][6] ), 
	.D(n3756), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][5]  (.Q(\ram[198][5] ), 
	.D(n3755), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][4]  (.Q(\ram[198][4] ), 
	.D(n3754), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][3]  (.Q(\ram[198][3] ), 
	.D(n3753), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][2]  (.Q(\ram[198][2] ), 
	.D(n3752), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][1]  (.Q(\ram[198][1] ), 
	.D(n3751), 
	.CK(clk));
   DFFHQX1 \ram_reg[198][0]  (.Q(\ram[198][0] ), 
	.D(n3750), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][15]  (.Q(\ram[194][15] ), 
	.D(n3701), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][14]  (.Q(\ram[194][14] ), 
	.D(n3700), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][13]  (.Q(\ram[194][13] ), 
	.D(n3699), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][12]  (.Q(\ram[194][12] ), 
	.D(n3698), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][11]  (.Q(\ram[194][11] ), 
	.D(n3697), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][10]  (.Q(\ram[194][10] ), 
	.D(n3696), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][9]  (.Q(\ram[194][9] ), 
	.D(n3695), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][8]  (.Q(\ram[194][8] ), 
	.D(n3694), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][7]  (.Q(\ram[194][7] ), 
	.D(n3693), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][6]  (.Q(\ram[194][6] ), 
	.D(n3692), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][5]  (.Q(\ram[194][5] ), 
	.D(n3691), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][4]  (.Q(\ram[194][4] ), 
	.D(n3690), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][3]  (.Q(\ram[194][3] ), 
	.D(n3689), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][2]  (.Q(\ram[194][2] ), 
	.D(n3688), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][1]  (.Q(\ram[194][1] ), 
	.D(n3687), 
	.CK(clk));
   DFFHQX1 \ram_reg[194][0]  (.Q(\ram[194][0] ), 
	.D(n3686), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][15]  (.Q(\ram[190][15] ), 
	.D(n3637), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][14]  (.Q(\ram[190][14] ), 
	.D(n3636), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][13]  (.Q(\ram[190][13] ), 
	.D(n3635), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][12]  (.Q(\ram[190][12] ), 
	.D(n3634), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][11]  (.Q(\ram[190][11] ), 
	.D(n3633), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][10]  (.Q(\ram[190][10] ), 
	.D(n3632), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][9]  (.Q(\ram[190][9] ), 
	.D(n3631), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][8]  (.Q(\ram[190][8] ), 
	.D(n3630), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][7]  (.Q(\ram[190][7] ), 
	.D(n3629), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][6]  (.Q(\ram[190][6] ), 
	.D(n3628), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][5]  (.Q(\ram[190][5] ), 
	.D(n3627), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][4]  (.Q(\ram[190][4] ), 
	.D(n3626), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][3]  (.Q(\ram[190][3] ), 
	.D(n3625), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][2]  (.Q(\ram[190][2] ), 
	.D(n3624), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][1]  (.Q(\ram[190][1] ), 
	.D(n3623), 
	.CK(clk));
   DFFHQX1 \ram_reg[190][0]  (.Q(\ram[190][0] ), 
	.D(n3622), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][15]  (.Q(\ram[186][15] ), 
	.D(n3573), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][14]  (.Q(\ram[186][14] ), 
	.D(n3572), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][13]  (.Q(\ram[186][13] ), 
	.D(n3571), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][12]  (.Q(\ram[186][12] ), 
	.D(n3570), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][11]  (.Q(\ram[186][11] ), 
	.D(n3569), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][10]  (.Q(\ram[186][10] ), 
	.D(n3568), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][9]  (.Q(\ram[186][9] ), 
	.D(n3567), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][8]  (.Q(\ram[186][8] ), 
	.D(n3566), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][7]  (.Q(\ram[186][7] ), 
	.D(n3565), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][6]  (.Q(\ram[186][6] ), 
	.D(n3564), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][5]  (.Q(\ram[186][5] ), 
	.D(n3563), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][4]  (.Q(\ram[186][4] ), 
	.D(n3562), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][3]  (.Q(\ram[186][3] ), 
	.D(n3561), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][2]  (.Q(\ram[186][2] ), 
	.D(n3560), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][1]  (.Q(\ram[186][1] ), 
	.D(n3559), 
	.CK(clk));
   DFFHQX1 \ram_reg[186][0]  (.Q(\ram[186][0] ), 
	.D(n3558), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][15]  (.Q(\ram[182][15] ), 
	.D(n3509), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][14]  (.Q(\ram[182][14] ), 
	.D(n3508), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][13]  (.Q(\ram[182][13] ), 
	.D(n3507), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][12]  (.Q(\ram[182][12] ), 
	.D(n3506), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][11]  (.Q(\ram[182][11] ), 
	.D(n3505), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][10]  (.Q(\ram[182][10] ), 
	.D(n3504), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][9]  (.Q(\ram[182][9] ), 
	.D(n3503), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][8]  (.Q(\ram[182][8] ), 
	.D(n3502), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][7]  (.Q(\ram[182][7] ), 
	.D(n3501), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][6]  (.Q(\ram[182][6] ), 
	.D(n3500), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][5]  (.Q(\ram[182][5] ), 
	.D(n3499), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][4]  (.Q(\ram[182][4] ), 
	.D(n3498), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][3]  (.Q(\ram[182][3] ), 
	.D(n3497), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][2]  (.Q(\ram[182][2] ), 
	.D(n3496), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][1]  (.Q(\ram[182][1] ), 
	.D(n3495), 
	.CK(clk));
   DFFHQX1 \ram_reg[182][0]  (.Q(\ram[182][0] ), 
	.D(n3494), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][15]  (.Q(\ram[178][15] ), 
	.D(n3445), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][14]  (.Q(\ram[178][14] ), 
	.D(n3444), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][13]  (.Q(\ram[178][13] ), 
	.D(n3443), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][12]  (.Q(\ram[178][12] ), 
	.D(n3442), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][11]  (.Q(\ram[178][11] ), 
	.D(n3441), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][10]  (.Q(\ram[178][10] ), 
	.D(n3440), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][9]  (.Q(\ram[178][9] ), 
	.D(n3439), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][8]  (.Q(\ram[178][8] ), 
	.D(n3438), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][7]  (.Q(\ram[178][7] ), 
	.D(n3437), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][6]  (.Q(\ram[178][6] ), 
	.D(n3436), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][5]  (.Q(\ram[178][5] ), 
	.D(n3435), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][4]  (.Q(\ram[178][4] ), 
	.D(n3434), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][3]  (.Q(\ram[178][3] ), 
	.D(n3433), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][2]  (.Q(\ram[178][2] ), 
	.D(n3432), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][1]  (.Q(\ram[178][1] ), 
	.D(n3431), 
	.CK(clk));
   DFFHQX1 \ram_reg[178][0]  (.Q(\ram[178][0] ), 
	.D(n3430), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][15]  (.Q(\ram[174][15] ), 
	.D(n3381), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][14]  (.Q(\ram[174][14] ), 
	.D(n3380), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][13]  (.Q(\ram[174][13] ), 
	.D(n3379), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][12]  (.Q(\ram[174][12] ), 
	.D(n3378), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][11]  (.Q(\ram[174][11] ), 
	.D(n3377), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][10]  (.Q(\ram[174][10] ), 
	.D(n3376), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][9]  (.Q(\ram[174][9] ), 
	.D(n3375), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][8]  (.Q(\ram[174][8] ), 
	.D(n3374), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][7]  (.Q(\ram[174][7] ), 
	.D(n3373), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][6]  (.Q(\ram[174][6] ), 
	.D(n3372), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][5]  (.Q(\ram[174][5] ), 
	.D(n3371), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][4]  (.Q(\ram[174][4] ), 
	.D(n3370), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][3]  (.Q(\ram[174][3] ), 
	.D(n3369), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][2]  (.Q(\ram[174][2] ), 
	.D(n3368), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][1]  (.Q(\ram[174][1] ), 
	.D(n3367), 
	.CK(clk));
   DFFHQX1 \ram_reg[174][0]  (.Q(\ram[174][0] ), 
	.D(n3366), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][15]  (.Q(\ram[170][15] ), 
	.D(n3317), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][14]  (.Q(\ram[170][14] ), 
	.D(n3316), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][13]  (.Q(\ram[170][13] ), 
	.D(n3315), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][12]  (.Q(\ram[170][12] ), 
	.D(n3314), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][11]  (.Q(\ram[170][11] ), 
	.D(n3313), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][10]  (.Q(\ram[170][10] ), 
	.D(n3312), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][9]  (.Q(\ram[170][9] ), 
	.D(n3311), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][8]  (.Q(\ram[170][8] ), 
	.D(n3310), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][7]  (.Q(\ram[170][7] ), 
	.D(n3309), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][6]  (.Q(\ram[170][6] ), 
	.D(n3308), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][5]  (.Q(\ram[170][5] ), 
	.D(n3307), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][4]  (.Q(\ram[170][4] ), 
	.D(n3306), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][3]  (.Q(\ram[170][3] ), 
	.D(n3305), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][2]  (.Q(\ram[170][2] ), 
	.D(n3304), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][1]  (.Q(\ram[170][1] ), 
	.D(n3303), 
	.CK(clk));
   DFFHQX1 \ram_reg[170][0]  (.Q(\ram[170][0] ), 
	.D(n3302), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][15]  (.Q(\ram[166][15] ), 
	.D(n3253), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][14]  (.Q(\ram[166][14] ), 
	.D(n3252), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][13]  (.Q(\ram[166][13] ), 
	.D(n3251), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][12]  (.Q(\ram[166][12] ), 
	.D(n3250), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][11]  (.Q(\ram[166][11] ), 
	.D(n3249), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][10]  (.Q(\ram[166][10] ), 
	.D(n3248), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][9]  (.Q(\ram[166][9] ), 
	.D(n3247), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][8]  (.Q(\ram[166][8] ), 
	.D(n3246), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][7]  (.Q(\ram[166][7] ), 
	.D(n3245), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][6]  (.Q(\ram[166][6] ), 
	.D(n3244), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][5]  (.Q(\ram[166][5] ), 
	.D(n3243), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][4]  (.Q(\ram[166][4] ), 
	.D(n3242), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][3]  (.Q(\ram[166][3] ), 
	.D(n3241), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][2]  (.Q(\ram[166][2] ), 
	.D(n3240), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][1]  (.Q(\ram[166][1] ), 
	.D(n3239), 
	.CK(clk));
   DFFHQX1 \ram_reg[166][0]  (.Q(\ram[166][0] ), 
	.D(n3238), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][15]  (.Q(\ram[162][15] ), 
	.D(n3189), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][14]  (.Q(\ram[162][14] ), 
	.D(n3188), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][13]  (.Q(\ram[162][13] ), 
	.D(n3187), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][12]  (.Q(\ram[162][12] ), 
	.D(n3186), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][11]  (.Q(\ram[162][11] ), 
	.D(n3185), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][10]  (.Q(\ram[162][10] ), 
	.D(n3184), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][9]  (.Q(\ram[162][9] ), 
	.D(n3183), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][8]  (.Q(\ram[162][8] ), 
	.D(n3182), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][7]  (.Q(\ram[162][7] ), 
	.D(n3181), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][6]  (.Q(\ram[162][6] ), 
	.D(n3180), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][5]  (.Q(\ram[162][5] ), 
	.D(n3179), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][4]  (.Q(\ram[162][4] ), 
	.D(n3178), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][3]  (.Q(\ram[162][3] ), 
	.D(n3177), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][2]  (.Q(\ram[162][2] ), 
	.D(n3176), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][1]  (.Q(\ram[162][1] ), 
	.D(n3175), 
	.CK(clk));
   DFFHQX1 \ram_reg[162][0]  (.Q(\ram[162][0] ), 
	.D(n3174), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][15]  (.Q(\ram[158][15] ), 
	.D(n3125), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][14]  (.Q(\ram[158][14] ), 
	.D(n3124), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][13]  (.Q(\ram[158][13] ), 
	.D(n3123), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][12]  (.Q(\ram[158][12] ), 
	.D(n3122), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][11]  (.Q(\ram[158][11] ), 
	.D(n3121), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][10]  (.Q(\ram[158][10] ), 
	.D(n3120), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][9]  (.Q(\ram[158][9] ), 
	.D(n3119), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][8]  (.Q(\ram[158][8] ), 
	.D(n3118), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][7]  (.Q(\ram[158][7] ), 
	.D(n3117), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][6]  (.Q(\ram[158][6] ), 
	.D(n3116), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][5]  (.Q(\ram[158][5] ), 
	.D(n3115), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][4]  (.Q(\ram[158][4] ), 
	.D(n3114), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][3]  (.Q(\ram[158][3] ), 
	.D(n3113), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][2]  (.Q(\ram[158][2] ), 
	.D(n3112), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][1]  (.Q(\ram[158][1] ), 
	.D(n3111), 
	.CK(clk));
   DFFHQX1 \ram_reg[158][0]  (.Q(\ram[158][0] ), 
	.D(n3110), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][15]  (.Q(\ram[154][15] ), 
	.D(n3061), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][14]  (.Q(\ram[154][14] ), 
	.D(n3060), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][13]  (.Q(\ram[154][13] ), 
	.D(n3059), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][12]  (.Q(\ram[154][12] ), 
	.D(n3058), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][11]  (.Q(\ram[154][11] ), 
	.D(n3057), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][10]  (.Q(\ram[154][10] ), 
	.D(n3056), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][9]  (.Q(\ram[154][9] ), 
	.D(n3055), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][8]  (.Q(\ram[154][8] ), 
	.D(n3054), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][7]  (.Q(\ram[154][7] ), 
	.D(n3053), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][6]  (.Q(\ram[154][6] ), 
	.D(n3052), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][5]  (.Q(\ram[154][5] ), 
	.D(n3051), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][4]  (.Q(\ram[154][4] ), 
	.D(n3050), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][3]  (.Q(\ram[154][3] ), 
	.D(n3049), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][2]  (.Q(\ram[154][2] ), 
	.D(n3048), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][1]  (.Q(\ram[154][1] ), 
	.D(n3047), 
	.CK(clk));
   DFFHQX1 \ram_reg[154][0]  (.Q(\ram[154][0] ), 
	.D(n3046), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][15]  (.Q(\ram[150][15] ), 
	.D(n2997), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][14]  (.Q(\ram[150][14] ), 
	.D(n2996), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][13]  (.Q(\ram[150][13] ), 
	.D(n2995), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][12]  (.Q(\ram[150][12] ), 
	.D(n2994), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][11]  (.Q(\ram[150][11] ), 
	.D(n2993), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][10]  (.Q(\ram[150][10] ), 
	.D(n2992), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][9]  (.Q(\ram[150][9] ), 
	.D(n2991), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][8]  (.Q(\ram[150][8] ), 
	.D(n2990), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][7]  (.Q(\ram[150][7] ), 
	.D(n2989), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][6]  (.Q(\ram[150][6] ), 
	.D(n2988), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][5]  (.Q(\ram[150][5] ), 
	.D(n2987), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][4]  (.Q(\ram[150][4] ), 
	.D(n2986), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][3]  (.Q(\ram[150][3] ), 
	.D(n2985), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][2]  (.Q(\ram[150][2] ), 
	.D(n2984), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][1]  (.Q(\ram[150][1] ), 
	.D(n2983), 
	.CK(clk));
   DFFHQX1 \ram_reg[150][0]  (.Q(\ram[150][0] ), 
	.D(n2982), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][15]  (.Q(\ram[146][15] ), 
	.D(n2933), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][14]  (.Q(\ram[146][14] ), 
	.D(n2932), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][13]  (.Q(\ram[146][13] ), 
	.D(n2931), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][12]  (.Q(\ram[146][12] ), 
	.D(n2930), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][11]  (.Q(\ram[146][11] ), 
	.D(n2929), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][10]  (.Q(\ram[146][10] ), 
	.D(n2928), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][9]  (.Q(\ram[146][9] ), 
	.D(n2927), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][8]  (.Q(\ram[146][8] ), 
	.D(n2926), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][7]  (.Q(\ram[146][7] ), 
	.D(n2925), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][6]  (.Q(\ram[146][6] ), 
	.D(n2924), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][5]  (.Q(\ram[146][5] ), 
	.D(n2923), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][4]  (.Q(\ram[146][4] ), 
	.D(n2922), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][3]  (.Q(\ram[146][3] ), 
	.D(n2921), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][2]  (.Q(\ram[146][2] ), 
	.D(n2920), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][1]  (.Q(\ram[146][1] ), 
	.D(n2919), 
	.CK(clk));
   DFFHQX1 \ram_reg[146][0]  (.Q(\ram[146][0] ), 
	.D(n2918), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][15]  (.Q(\ram[142][15] ), 
	.D(n2869), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][14]  (.Q(\ram[142][14] ), 
	.D(n2868), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][13]  (.Q(\ram[142][13] ), 
	.D(n2867), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][12]  (.Q(\ram[142][12] ), 
	.D(n2866), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][11]  (.Q(\ram[142][11] ), 
	.D(n2865), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][10]  (.Q(\ram[142][10] ), 
	.D(n2864), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][9]  (.Q(\ram[142][9] ), 
	.D(n2863), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][8]  (.Q(\ram[142][8] ), 
	.D(n2862), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][7]  (.Q(\ram[142][7] ), 
	.D(n2861), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][6]  (.Q(\ram[142][6] ), 
	.D(n2860), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][5]  (.Q(\ram[142][5] ), 
	.D(n2859), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][4]  (.Q(\ram[142][4] ), 
	.D(n2858), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][3]  (.Q(\ram[142][3] ), 
	.D(n2857), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][2]  (.Q(\ram[142][2] ), 
	.D(n2856), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][1]  (.Q(\ram[142][1] ), 
	.D(n2855), 
	.CK(clk));
   DFFHQX1 \ram_reg[142][0]  (.Q(\ram[142][0] ), 
	.D(n2854), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][15]  (.Q(\ram[138][15] ), 
	.D(n2805), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][14]  (.Q(\ram[138][14] ), 
	.D(n2804), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][13]  (.Q(\ram[138][13] ), 
	.D(n2803), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][12]  (.Q(\ram[138][12] ), 
	.D(n2802), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][11]  (.Q(\ram[138][11] ), 
	.D(n2801), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][10]  (.Q(\ram[138][10] ), 
	.D(n2800), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][9]  (.Q(\ram[138][9] ), 
	.D(n2799), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][8]  (.Q(\ram[138][8] ), 
	.D(n2798), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][7]  (.Q(\ram[138][7] ), 
	.D(n2797), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][6]  (.Q(\ram[138][6] ), 
	.D(n2796), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][5]  (.Q(\ram[138][5] ), 
	.D(n2795), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][4]  (.Q(\ram[138][4] ), 
	.D(n2794), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][3]  (.Q(\ram[138][3] ), 
	.D(n2793), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][2]  (.Q(\ram[138][2] ), 
	.D(n2792), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][1]  (.Q(\ram[138][1] ), 
	.D(n2791), 
	.CK(clk));
   DFFHQX1 \ram_reg[138][0]  (.Q(\ram[138][0] ), 
	.D(n2790), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][15]  (.Q(\ram[134][15] ), 
	.D(n2741), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][14]  (.Q(\ram[134][14] ), 
	.D(n2740), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][13]  (.Q(\ram[134][13] ), 
	.D(n2739), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][12]  (.Q(\ram[134][12] ), 
	.D(n2738), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][11]  (.Q(\ram[134][11] ), 
	.D(n2737), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][10]  (.Q(\ram[134][10] ), 
	.D(n2736), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][9]  (.Q(\ram[134][9] ), 
	.D(n2735), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][8]  (.Q(\ram[134][8] ), 
	.D(n2734), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][7]  (.Q(\ram[134][7] ), 
	.D(n2733), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][6]  (.Q(\ram[134][6] ), 
	.D(n2732), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][5]  (.Q(\ram[134][5] ), 
	.D(n2731), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][4]  (.Q(\ram[134][4] ), 
	.D(n2730), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][3]  (.Q(\ram[134][3] ), 
	.D(n2729), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][2]  (.Q(\ram[134][2] ), 
	.D(n2728), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][1]  (.Q(\ram[134][1] ), 
	.D(n2727), 
	.CK(clk));
   DFFHQX1 \ram_reg[134][0]  (.Q(\ram[134][0] ), 
	.D(n2726), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][15]  (.Q(\ram[130][15] ), 
	.D(n2677), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][14]  (.Q(\ram[130][14] ), 
	.D(n2676), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][13]  (.Q(\ram[130][13] ), 
	.D(n2675), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][12]  (.Q(\ram[130][12] ), 
	.D(n2674), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][11]  (.Q(\ram[130][11] ), 
	.D(n2673), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][10]  (.Q(\ram[130][10] ), 
	.D(n2672), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][9]  (.Q(\ram[130][9] ), 
	.D(n2671), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][8]  (.Q(\ram[130][8] ), 
	.D(n2670), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][7]  (.Q(\ram[130][7] ), 
	.D(n2669), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][6]  (.Q(\ram[130][6] ), 
	.D(n2668), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][5]  (.Q(\ram[130][5] ), 
	.D(n2667), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][4]  (.Q(\ram[130][4] ), 
	.D(n2666), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][3]  (.Q(\ram[130][3] ), 
	.D(n2665), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][2]  (.Q(\ram[130][2] ), 
	.D(n2664), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][1]  (.Q(\ram[130][1] ), 
	.D(n2663), 
	.CK(clk));
   DFFHQX1 \ram_reg[130][0]  (.Q(\ram[130][0] ), 
	.D(n2662), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][15]  (.Q(\ram[126][15] ), 
	.D(n2613), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][14]  (.Q(\ram[126][14] ), 
	.D(n2612), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][13]  (.Q(\ram[126][13] ), 
	.D(n2611), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][12]  (.Q(\ram[126][12] ), 
	.D(n2610), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][11]  (.Q(\ram[126][11] ), 
	.D(n2609), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][10]  (.Q(\ram[126][10] ), 
	.D(n2608), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][9]  (.Q(\ram[126][9] ), 
	.D(n2607), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][8]  (.Q(\ram[126][8] ), 
	.D(n2606), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][7]  (.Q(\ram[126][7] ), 
	.D(n2605), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][6]  (.Q(\ram[126][6] ), 
	.D(n2604), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][5]  (.Q(\ram[126][5] ), 
	.D(n2603), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][4]  (.Q(\ram[126][4] ), 
	.D(n2602), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][3]  (.Q(\ram[126][3] ), 
	.D(n2601), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][2]  (.Q(\ram[126][2] ), 
	.D(n2600), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][1]  (.Q(\ram[126][1] ), 
	.D(n2599), 
	.CK(clk));
   DFFHQX1 \ram_reg[126][0]  (.Q(\ram[126][0] ), 
	.D(n2598), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][15]  (.Q(\ram[122][15] ), 
	.D(n2549), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][14]  (.Q(\ram[122][14] ), 
	.D(n2548), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][13]  (.Q(\ram[122][13] ), 
	.D(n2547), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][12]  (.Q(\ram[122][12] ), 
	.D(n2546), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][11]  (.Q(\ram[122][11] ), 
	.D(n2545), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][10]  (.Q(\ram[122][10] ), 
	.D(n2544), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][9]  (.Q(\ram[122][9] ), 
	.D(n2543), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][8]  (.Q(\ram[122][8] ), 
	.D(n2542), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][7]  (.Q(\ram[122][7] ), 
	.D(n2541), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][6]  (.Q(\ram[122][6] ), 
	.D(n2540), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][5]  (.Q(\ram[122][5] ), 
	.D(n2539), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][4]  (.Q(\ram[122][4] ), 
	.D(n2538), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][3]  (.Q(\ram[122][3] ), 
	.D(n2537), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][2]  (.Q(\ram[122][2] ), 
	.D(n2536), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][1]  (.Q(\ram[122][1] ), 
	.D(n2535), 
	.CK(clk));
   DFFHQX1 \ram_reg[122][0]  (.Q(\ram[122][0] ), 
	.D(n2534), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][15]  (.Q(\ram[118][15] ), 
	.D(n2485), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][14]  (.Q(\ram[118][14] ), 
	.D(n2484), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][13]  (.Q(\ram[118][13] ), 
	.D(n2483), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][12]  (.Q(\ram[118][12] ), 
	.D(n2482), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][11]  (.Q(\ram[118][11] ), 
	.D(n2481), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][10]  (.Q(\ram[118][10] ), 
	.D(n2480), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][9]  (.Q(\ram[118][9] ), 
	.D(n2479), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][8]  (.Q(\ram[118][8] ), 
	.D(n2478), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][7]  (.Q(\ram[118][7] ), 
	.D(n2477), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][6]  (.Q(\ram[118][6] ), 
	.D(n2476), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][5]  (.Q(\ram[118][5] ), 
	.D(n2475), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][4]  (.Q(\ram[118][4] ), 
	.D(n2474), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][3]  (.Q(\ram[118][3] ), 
	.D(n2473), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][2]  (.Q(\ram[118][2] ), 
	.D(n2472), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][1]  (.Q(\ram[118][1] ), 
	.D(n2471), 
	.CK(clk));
   DFFHQX1 \ram_reg[118][0]  (.Q(\ram[118][0] ), 
	.D(n2470), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][15]  (.Q(\ram[114][15] ), 
	.D(n2421), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][14]  (.Q(\ram[114][14] ), 
	.D(n2420), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][13]  (.Q(\ram[114][13] ), 
	.D(n2419), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][12]  (.Q(\ram[114][12] ), 
	.D(n2418), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][11]  (.Q(\ram[114][11] ), 
	.D(n2417), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][10]  (.Q(\ram[114][10] ), 
	.D(n2416), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][9]  (.Q(\ram[114][9] ), 
	.D(n2415), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][8]  (.Q(\ram[114][8] ), 
	.D(n2414), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][7]  (.Q(\ram[114][7] ), 
	.D(n2413), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][6]  (.Q(\ram[114][6] ), 
	.D(n2412), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][5]  (.Q(\ram[114][5] ), 
	.D(n2411), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][4]  (.Q(\ram[114][4] ), 
	.D(n2410), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][3]  (.Q(\ram[114][3] ), 
	.D(n2409), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][2]  (.Q(\ram[114][2] ), 
	.D(n2408), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][1]  (.Q(\ram[114][1] ), 
	.D(n2407), 
	.CK(clk));
   DFFHQX1 \ram_reg[114][0]  (.Q(\ram[114][0] ), 
	.D(n2406), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][15]  (.Q(\ram[110][15] ), 
	.D(n2357), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][14]  (.Q(\ram[110][14] ), 
	.D(n2356), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][13]  (.Q(\ram[110][13] ), 
	.D(n2355), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][12]  (.Q(\ram[110][12] ), 
	.D(n2354), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][11]  (.Q(\ram[110][11] ), 
	.D(n2353), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][10]  (.Q(\ram[110][10] ), 
	.D(n2352), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][9]  (.Q(\ram[110][9] ), 
	.D(n2351), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][8]  (.Q(\ram[110][8] ), 
	.D(n2350), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][7]  (.Q(\ram[110][7] ), 
	.D(n2349), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][6]  (.Q(\ram[110][6] ), 
	.D(n2348), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][5]  (.Q(\ram[110][5] ), 
	.D(n2347), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][4]  (.Q(\ram[110][4] ), 
	.D(n2346), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][3]  (.Q(\ram[110][3] ), 
	.D(n2345), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][2]  (.Q(\ram[110][2] ), 
	.D(n2344), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][1]  (.Q(\ram[110][1] ), 
	.D(n2343), 
	.CK(clk));
   DFFHQX1 \ram_reg[110][0]  (.Q(\ram[110][0] ), 
	.D(n2342), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][15]  (.Q(\ram[106][15] ), 
	.D(n2293), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][14]  (.Q(\ram[106][14] ), 
	.D(n2292), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][13]  (.Q(\ram[106][13] ), 
	.D(n2291), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][12]  (.Q(\ram[106][12] ), 
	.D(n2290), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][11]  (.Q(\ram[106][11] ), 
	.D(n2289), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][10]  (.Q(\ram[106][10] ), 
	.D(n2288), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][9]  (.Q(\ram[106][9] ), 
	.D(n2287), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][8]  (.Q(\ram[106][8] ), 
	.D(n2286), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][7]  (.Q(\ram[106][7] ), 
	.D(n2285), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][6]  (.Q(\ram[106][6] ), 
	.D(n2284), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][5]  (.Q(\ram[106][5] ), 
	.D(n2283), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][4]  (.Q(\ram[106][4] ), 
	.D(n2282), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][3]  (.Q(\ram[106][3] ), 
	.D(n2281), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][2]  (.Q(\ram[106][2] ), 
	.D(n2280), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][1]  (.Q(\ram[106][1] ), 
	.D(n2279), 
	.CK(clk));
   DFFHQX1 \ram_reg[106][0]  (.Q(\ram[106][0] ), 
	.D(n2278), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][15]  (.Q(\ram[102][15] ), 
	.D(n2229), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][14]  (.Q(\ram[102][14] ), 
	.D(n2228), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][13]  (.Q(\ram[102][13] ), 
	.D(n2227), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][12]  (.Q(\ram[102][12] ), 
	.D(n2226), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][11]  (.Q(\ram[102][11] ), 
	.D(n2225), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][10]  (.Q(\ram[102][10] ), 
	.D(n2224), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][9]  (.Q(\ram[102][9] ), 
	.D(n2223), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][8]  (.Q(\ram[102][8] ), 
	.D(n2222), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][7]  (.Q(\ram[102][7] ), 
	.D(n2221), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][6]  (.Q(\ram[102][6] ), 
	.D(n2220), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][5]  (.Q(\ram[102][5] ), 
	.D(n2219), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][4]  (.Q(\ram[102][4] ), 
	.D(n2218), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][3]  (.Q(\ram[102][3] ), 
	.D(n2217), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][2]  (.Q(\ram[102][2] ), 
	.D(n2216), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][1]  (.Q(\ram[102][1] ), 
	.D(n2215), 
	.CK(clk));
   DFFHQX1 \ram_reg[102][0]  (.Q(\ram[102][0] ), 
	.D(n2214), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][15]  (.Q(\ram[98][15] ), 
	.D(n2165), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][14]  (.Q(\ram[98][14] ), 
	.D(n2164), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][13]  (.Q(\ram[98][13] ), 
	.D(n2163), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][12]  (.Q(\ram[98][12] ), 
	.D(n2162), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][11]  (.Q(\ram[98][11] ), 
	.D(n2161), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][10]  (.Q(\ram[98][10] ), 
	.D(n2160), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][9]  (.Q(\ram[98][9] ), 
	.D(n2159), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][8]  (.Q(\ram[98][8] ), 
	.D(n2158), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][7]  (.Q(\ram[98][7] ), 
	.D(n2157), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][6]  (.Q(\ram[98][6] ), 
	.D(n2156), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][5]  (.Q(\ram[98][5] ), 
	.D(n2155), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][4]  (.Q(\ram[98][4] ), 
	.D(n2154), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][3]  (.Q(\ram[98][3] ), 
	.D(n2153), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][2]  (.Q(\ram[98][2] ), 
	.D(n2152), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][1]  (.Q(\ram[98][1] ), 
	.D(n2151), 
	.CK(clk));
   DFFHQX1 \ram_reg[98][0]  (.Q(\ram[98][0] ), 
	.D(n2150), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][15]  (.Q(\ram[94][15] ), 
	.D(n2101), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][14]  (.Q(\ram[94][14] ), 
	.D(n2100), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][13]  (.Q(\ram[94][13] ), 
	.D(n2099), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][12]  (.Q(\ram[94][12] ), 
	.D(n2098), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][11]  (.Q(\ram[94][11] ), 
	.D(n2097), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][10]  (.Q(\ram[94][10] ), 
	.D(n2096), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][9]  (.Q(\ram[94][9] ), 
	.D(n2095), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][8]  (.Q(\ram[94][8] ), 
	.D(n2094), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][7]  (.Q(\ram[94][7] ), 
	.D(n2093), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][6]  (.Q(\ram[94][6] ), 
	.D(n2092), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][5]  (.Q(\ram[94][5] ), 
	.D(n2091), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][4]  (.Q(\ram[94][4] ), 
	.D(n2090), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][3]  (.Q(\ram[94][3] ), 
	.D(n2089), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][2]  (.Q(\ram[94][2] ), 
	.D(n2088), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][1]  (.Q(\ram[94][1] ), 
	.D(n2087), 
	.CK(clk));
   DFFHQX1 \ram_reg[94][0]  (.Q(\ram[94][0] ), 
	.D(n2086), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][15]  (.Q(\ram[90][15] ), 
	.D(n2037), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][14]  (.Q(\ram[90][14] ), 
	.D(n2036), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][13]  (.Q(\ram[90][13] ), 
	.D(n2035), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][12]  (.Q(\ram[90][12] ), 
	.D(n2034), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][11]  (.Q(\ram[90][11] ), 
	.D(n2033), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][10]  (.Q(\ram[90][10] ), 
	.D(n2032), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][9]  (.Q(\ram[90][9] ), 
	.D(n2031), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][8]  (.Q(\ram[90][8] ), 
	.D(n2030), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][7]  (.Q(\ram[90][7] ), 
	.D(n2029), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][6]  (.Q(\ram[90][6] ), 
	.D(n2028), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][5]  (.Q(\ram[90][5] ), 
	.D(n2027), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][4]  (.Q(\ram[90][4] ), 
	.D(n2026), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][3]  (.Q(\ram[90][3] ), 
	.D(n2025), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][2]  (.Q(\ram[90][2] ), 
	.D(n2024), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][1]  (.Q(\ram[90][1] ), 
	.D(n2023), 
	.CK(clk));
   DFFHQX1 \ram_reg[90][0]  (.Q(\ram[90][0] ), 
	.D(n2022), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][15]  (.Q(\ram[86][15] ), 
	.D(n1973), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][14]  (.Q(\ram[86][14] ), 
	.D(n1972), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][13]  (.Q(\ram[86][13] ), 
	.D(n1971), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][12]  (.Q(\ram[86][12] ), 
	.D(n1970), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][11]  (.Q(\ram[86][11] ), 
	.D(n1969), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][10]  (.Q(\ram[86][10] ), 
	.D(n1968), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][9]  (.Q(\ram[86][9] ), 
	.D(n1967), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][8]  (.Q(\ram[86][8] ), 
	.D(n1966), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][7]  (.Q(\ram[86][7] ), 
	.D(n1965), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][6]  (.Q(\ram[86][6] ), 
	.D(n1964), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][5]  (.Q(\ram[86][5] ), 
	.D(n1963), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][4]  (.Q(\ram[86][4] ), 
	.D(n1962), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][3]  (.Q(\ram[86][3] ), 
	.D(n1961), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][2]  (.Q(\ram[86][2] ), 
	.D(n1960), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][1]  (.Q(\ram[86][1] ), 
	.D(n1959), 
	.CK(clk));
   DFFHQX1 \ram_reg[86][0]  (.Q(\ram[86][0] ), 
	.D(n1958), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][15]  (.Q(\ram[82][15] ), 
	.D(n1909), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][14]  (.Q(\ram[82][14] ), 
	.D(n1908), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][13]  (.Q(\ram[82][13] ), 
	.D(n1907), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][12]  (.Q(\ram[82][12] ), 
	.D(n1906), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][11]  (.Q(\ram[82][11] ), 
	.D(n1905), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][10]  (.Q(\ram[82][10] ), 
	.D(n1904), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][9]  (.Q(\ram[82][9] ), 
	.D(n1903), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][8]  (.Q(\ram[82][8] ), 
	.D(n1902), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][7]  (.Q(\ram[82][7] ), 
	.D(n1901), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][6]  (.Q(\ram[82][6] ), 
	.D(n1900), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][5]  (.Q(\ram[82][5] ), 
	.D(n1899), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][4]  (.Q(\ram[82][4] ), 
	.D(n1898), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][3]  (.Q(\ram[82][3] ), 
	.D(n1897), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][2]  (.Q(\ram[82][2] ), 
	.D(n1896), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][1]  (.Q(\ram[82][1] ), 
	.D(n1895), 
	.CK(clk));
   DFFHQX1 \ram_reg[82][0]  (.Q(\ram[82][0] ), 
	.D(n1894), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][15]  (.Q(\ram[78][15] ), 
	.D(n1845), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][14]  (.Q(\ram[78][14] ), 
	.D(n1844), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][13]  (.Q(\ram[78][13] ), 
	.D(n1843), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][12]  (.Q(\ram[78][12] ), 
	.D(n1842), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][11]  (.Q(\ram[78][11] ), 
	.D(n1841), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][10]  (.Q(\ram[78][10] ), 
	.D(n1840), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][9]  (.Q(\ram[78][9] ), 
	.D(n1839), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][8]  (.Q(\ram[78][8] ), 
	.D(n1838), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][7]  (.Q(\ram[78][7] ), 
	.D(n1837), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][6]  (.Q(\ram[78][6] ), 
	.D(n1836), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][5]  (.Q(\ram[78][5] ), 
	.D(n1835), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][4]  (.Q(\ram[78][4] ), 
	.D(n1834), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][3]  (.Q(\ram[78][3] ), 
	.D(n1833), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][2]  (.Q(\ram[78][2] ), 
	.D(n1832), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][1]  (.Q(\ram[78][1] ), 
	.D(n1831), 
	.CK(clk));
   DFFHQX1 \ram_reg[78][0]  (.Q(\ram[78][0] ), 
	.D(n1830), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][15]  (.Q(\ram[74][15] ), 
	.D(n1781), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][14]  (.Q(\ram[74][14] ), 
	.D(n1780), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][13]  (.Q(\ram[74][13] ), 
	.D(n1779), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][12]  (.Q(\ram[74][12] ), 
	.D(n1778), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][11]  (.Q(\ram[74][11] ), 
	.D(n1777), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][10]  (.Q(\ram[74][10] ), 
	.D(n1776), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][9]  (.Q(\ram[74][9] ), 
	.D(n1775), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][8]  (.Q(\ram[74][8] ), 
	.D(n1774), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][7]  (.Q(\ram[74][7] ), 
	.D(n1773), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][6]  (.Q(\ram[74][6] ), 
	.D(n1772), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][5]  (.Q(\ram[74][5] ), 
	.D(n1771), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][4]  (.Q(\ram[74][4] ), 
	.D(n1770), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][3]  (.Q(\ram[74][3] ), 
	.D(n1769), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][2]  (.Q(\ram[74][2] ), 
	.D(n1768), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][1]  (.Q(\ram[74][1] ), 
	.D(n1767), 
	.CK(clk));
   DFFHQX1 \ram_reg[74][0]  (.Q(\ram[74][0] ), 
	.D(n1766), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][15]  (.Q(\ram[70][15] ), 
	.D(n1717), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][14]  (.Q(\ram[70][14] ), 
	.D(n1716), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][13]  (.Q(\ram[70][13] ), 
	.D(n1715), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][12]  (.Q(\ram[70][12] ), 
	.D(n1714), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][11]  (.Q(\ram[70][11] ), 
	.D(n1713), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][10]  (.Q(\ram[70][10] ), 
	.D(n1712), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][9]  (.Q(\ram[70][9] ), 
	.D(n1711), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][8]  (.Q(\ram[70][8] ), 
	.D(n1710), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][7]  (.Q(\ram[70][7] ), 
	.D(n1709), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][6]  (.Q(\ram[70][6] ), 
	.D(n1708), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][5]  (.Q(\ram[70][5] ), 
	.D(n1707), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][4]  (.Q(\ram[70][4] ), 
	.D(n1706), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][3]  (.Q(\ram[70][3] ), 
	.D(n1705), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][2]  (.Q(\ram[70][2] ), 
	.D(n1704), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][1]  (.Q(\ram[70][1] ), 
	.D(n1703), 
	.CK(clk));
   DFFHQX1 \ram_reg[70][0]  (.Q(\ram[70][0] ), 
	.D(n1702), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][15]  (.Q(\ram[66][15] ), 
	.D(n1653), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][14]  (.Q(\ram[66][14] ), 
	.D(n1652), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][13]  (.Q(\ram[66][13] ), 
	.D(n1651), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][12]  (.Q(\ram[66][12] ), 
	.D(n1650), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][11]  (.Q(\ram[66][11] ), 
	.D(n1649), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][10]  (.Q(\ram[66][10] ), 
	.D(n1648), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][9]  (.Q(\ram[66][9] ), 
	.D(n1647), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][8]  (.Q(\ram[66][8] ), 
	.D(n1646), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][7]  (.Q(\ram[66][7] ), 
	.D(n1645), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][6]  (.Q(\ram[66][6] ), 
	.D(n1644), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][5]  (.Q(\ram[66][5] ), 
	.D(n1643), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][4]  (.Q(\ram[66][4] ), 
	.D(n1642), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][3]  (.Q(\ram[66][3] ), 
	.D(n1641), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][2]  (.Q(\ram[66][2] ), 
	.D(n1640), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][1]  (.Q(\ram[66][1] ), 
	.D(n1639), 
	.CK(clk));
   DFFHQX1 \ram_reg[66][0]  (.Q(\ram[66][0] ), 
	.D(n1638), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][15]  (.Q(\ram[62][15] ), 
	.D(n1589), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][14]  (.Q(\ram[62][14] ), 
	.D(n1588), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][13]  (.Q(\ram[62][13] ), 
	.D(n1587), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][12]  (.Q(\ram[62][12] ), 
	.D(n1586), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][11]  (.Q(\ram[62][11] ), 
	.D(n1585), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][10]  (.Q(\ram[62][10] ), 
	.D(n1584), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][9]  (.Q(\ram[62][9] ), 
	.D(n1583), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][8]  (.Q(\ram[62][8] ), 
	.D(n1582), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][7]  (.Q(\ram[62][7] ), 
	.D(n1581), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][6]  (.Q(\ram[62][6] ), 
	.D(n1580), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][5]  (.Q(\ram[62][5] ), 
	.D(n1579), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][4]  (.Q(\ram[62][4] ), 
	.D(n1578), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][3]  (.Q(\ram[62][3] ), 
	.D(n1577), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][2]  (.Q(\ram[62][2] ), 
	.D(n1576), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][1]  (.Q(\ram[62][1] ), 
	.D(n1575), 
	.CK(clk));
   DFFHQX1 \ram_reg[62][0]  (.Q(\ram[62][0] ), 
	.D(n1574), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][15]  (.Q(\ram[58][15] ), 
	.D(n1525), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][14]  (.Q(\ram[58][14] ), 
	.D(n1524), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][13]  (.Q(\ram[58][13] ), 
	.D(n1523), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][12]  (.Q(\ram[58][12] ), 
	.D(n1522), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][11]  (.Q(\ram[58][11] ), 
	.D(n1521), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][10]  (.Q(\ram[58][10] ), 
	.D(n1520), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][9]  (.Q(\ram[58][9] ), 
	.D(n1519), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][8]  (.Q(\ram[58][8] ), 
	.D(n1518), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][7]  (.Q(\ram[58][7] ), 
	.D(n1517), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][6]  (.Q(\ram[58][6] ), 
	.D(n1516), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][5]  (.Q(\ram[58][5] ), 
	.D(n1515), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][4]  (.Q(\ram[58][4] ), 
	.D(n1514), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][3]  (.Q(\ram[58][3] ), 
	.D(n1513), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][2]  (.Q(\ram[58][2] ), 
	.D(n1512), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][1]  (.Q(\ram[58][1] ), 
	.D(n1511), 
	.CK(clk));
   DFFHQX1 \ram_reg[58][0]  (.Q(\ram[58][0] ), 
	.D(n1510), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][15]  (.Q(\ram[54][15] ), 
	.D(n1461), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][14]  (.Q(\ram[54][14] ), 
	.D(n1460), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][13]  (.Q(\ram[54][13] ), 
	.D(n1459), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][12]  (.Q(\ram[54][12] ), 
	.D(n1458), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][11]  (.Q(\ram[54][11] ), 
	.D(n1457), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][10]  (.Q(\ram[54][10] ), 
	.D(n1456), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][9]  (.Q(\ram[54][9] ), 
	.D(n1455), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][8]  (.Q(\ram[54][8] ), 
	.D(n1454), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][7]  (.Q(\ram[54][7] ), 
	.D(n1453), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][6]  (.Q(\ram[54][6] ), 
	.D(n1452), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][5]  (.Q(\ram[54][5] ), 
	.D(n1451), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][4]  (.Q(\ram[54][4] ), 
	.D(n1450), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][3]  (.Q(\ram[54][3] ), 
	.D(n1449), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][2]  (.Q(\ram[54][2] ), 
	.D(n1448), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][1]  (.Q(\ram[54][1] ), 
	.D(n1447), 
	.CK(clk));
   DFFHQX1 \ram_reg[54][0]  (.Q(\ram[54][0] ), 
	.D(n1446), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][15]  (.Q(\ram[50][15] ), 
	.D(n1397), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][14]  (.Q(\ram[50][14] ), 
	.D(n1396), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][13]  (.Q(\ram[50][13] ), 
	.D(n1395), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][12]  (.Q(\ram[50][12] ), 
	.D(n1394), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][11]  (.Q(\ram[50][11] ), 
	.D(n1393), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][10]  (.Q(\ram[50][10] ), 
	.D(n1392), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][9]  (.Q(\ram[50][9] ), 
	.D(n1391), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][8]  (.Q(\ram[50][8] ), 
	.D(n1390), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][7]  (.Q(\ram[50][7] ), 
	.D(n1389), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][6]  (.Q(\ram[50][6] ), 
	.D(n1388), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][5]  (.Q(\ram[50][5] ), 
	.D(n1387), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][4]  (.Q(\ram[50][4] ), 
	.D(n1386), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][3]  (.Q(\ram[50][3] ), 
	.D(n1385), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][2]  (.Q(\ram[50][2] ), 
	.D(n1384), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][1]  (.Q(\ram[50][1] ), 
	.D(n1383), 
	.CK(clk));
   DFFHQX1 \ram_reg[50][0]  (.Q(\ram[50][0] ), 
	.D(n1382), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][15]  (.Q(\ram[46][15] ), 
	.D(n1333), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][14]  (.Q(\ram[46][14] ), 
	.D(n1332), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][13]  (.Q(\ram[46][13] ), 
	.D(n1331), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][12]  (.Q(\ram[46][12] ), 
	.D(n1330), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][11]  (.Q(\ram[46][11] ), 
	.D(n1329), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][10]  (.Q(\ram[46][10] ), 
	.D(n1328), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][9]  (.Q(\ram[46][9] ), 
	.D(n1327), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][8]  (.Q(\ram[46][8] ), 
	.D(n1326), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][7]  (.Q(\ram[46][7] ), 
	.D(n1325), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][6]  (.Q(\ram[46][6] ), 
	.D(n1324), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][5]  (.Q(\ram[46][5] ), 
	.D(n1323), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][4]  (.Q(\ram[46][4] ), 
	.D(n1322), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][3]  (.Q(\ram[46][3] ), 
	.D(n1321), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][2]  (.Q(\ram[46][2] ), 
	.D(n1320), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][1]  (.Q(\ram[46][1] ), 
	.D(n1319), 
	.CK(clk));
   DFFHQX1 \ram_reg[46][0]  (.Q(\ram[46][0] ), 
	.D(n1318), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][15]  (.Q(\ram[42][15] ), 
	.D(n1269), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][14]  (.Q(\ram[42][14] ), 
	.D(n1268), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][13]  (.Q(\ram[42][13] ), 
	.D(n1267), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][12]  (.Q(\ram[42][12] ), 
	.D(n1266), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][11]  (.Q(\ram[42][11] ), 
	.D(n1265), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][10]  (.Q(\ram[42][10] ), 
	.D(n1264), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][9]  (.Q(\ram[42][9] ), 
	.D(n1263), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][8]  (.Q(\ram[42][8] ), 
	.D(n1262), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][7]  (.Q(\ram[42][7] ), 
	.D(n1261), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][6]  (.Q(\ram[42][6] ), 
	.D(n1260), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][5]  (.Q(\ram[42][5] ), 
	.D(n1259), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][4]  (.Q(\ram[42][4] ), 
	.D(n1258), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][3]  (.Q(\ram[42][3] ), 
	.D(n1257), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][2]  (.Q(\ram[42][2] ), 
	.D(n1256), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][1]  (.Q(\ram[42][1] ), 
	.D(n1255), 
	.CK(clk));
   DFFHQX1 \ram_reg[42][0]  (.Q(\ram[42][0] ), 
	.D(n1254), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][15]  (.Q(\ram[38][15] ), 
	.D(n1205), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][14]  (.Q(\ram[38][14] ), 
	.D(n1204), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][13]  (.Q(\ram[38][13] ), 
	.D(n1203), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][12]  (.Q(\ram[38][12] ), 
	.D(n1202), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][11]  (.Q(\ram[38][11] ), 
	.D(n1201), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][10]  (.Q(\ram[38][10] ), 
	.D(n1200), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][9]  (.Q(\ram[38][9] ), 
	.D(n1199), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][8]  (.Q(\ram[38][8] ), 
	.D(n1198), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][7]  (.Q(\ram[38][7] ), 
	.D(n1197), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][6]  (.Q(\ram[38][6] ), 
	.D(n1196), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][5]  (.Q(\ram[38][5] ), 
	.D(n1195), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][4]  (.Q(\ram[38][4] ), 
	.D(n1194), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][3]  (.Q(\ram[38][3] ), 
	.D(n1193), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][2]  (.Q(\ram[38][2] ), 
	.D(n1192), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][1]  (.Q(\ram[38][1] ), 
	.D(n1191), 
	.CK(clk));
   DFFHQX1 \ram_reg[38][0]  (.Q(\ram[38][0] ), 
	.D(n1190), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][15]  (.Q(\ram[34][15] ), 
	.D(n1141), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][14]  (.Q(\ram[34][14] ), 
	.D(n1140), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][13]  (.Q(\ram[34][13] ), 
	.D(n1139), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][12]  (.Q(\ram[34][12] ), 
	.D(n1138), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][11]  (.Q(\ram[34][11] ), 
	.D(n1137), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][10]  (.Q(\ram[34][10] ), 
	.D(n1136), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][9]  (.Q(\ram[34][9] ), 
	.D(n1135), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][8]  (.Q(\ram[34][8] ), 
	.D(n1134), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][7]  (.Q(\ram[34][7] ), 
	.D(n1133), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][6]  (.Q(\ram[34][6] ), 
	.D(n1132), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][5]  (.Q(\ram[34][5] ), 
	.D(n1131), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][4]  (.Q(\ram[34][4] ), 
	.D(n1130), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][3]  (.Q(\ram[34][3] ), 
	.D(n1129), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][2]  (.Q(\ram[34][2] ), 
	.D(n1128), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][1]  (.Q(\ram[34][1] ), 
	.D(n1127), 
	.CK(clk));
   DFFHQX1 \ram_reg[34][0]  (.Q(\ram[34][0] ), 
	.D(n1126), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][15]  (.Q(\ram[30][15] ), 
	.D(n1077), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][14]  (.Q(\ram[30][14] ), 
	.D(n1076), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][13]  (.Q(\ram[30][13] ), 
	.D(n1075), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][12]  (.Q(\ram[30][12] ), 
	.D(n1074), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][11]  (.Q(\ram[30][11] ), 
	.D(n1073), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][10]  (.Q(\ram[30][10] ), 
	.D(n1072), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][9]  (.Q(\ram[30][9] ), 
	.D(n1071), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][8]  (.Q(\ram[30][8] ), 
	.D(n1070), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][7]  (.Q(\ram[30][7] ), 
	.D(n1069), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][6]  (.Q(\ram[30][6] ), 
	.D(n1068), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][5]  (.Q(\ram[30][5] ), 
	.D(n1067), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][4]  (.Q(\ram[30][4] ), 
	.D(n1066), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][3]  (.Q(\ram[30][3] ), 
	.D(n1065), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][2]  (.Q(\ram[30][2] ), 
	.D(n1064), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][1]  (.Q(\ram[30][1] ), 
	.D(n1063), 
	.CK(clk));
   DFFHQX1 \ram_reg[30][0]  (.Q(\ram[30][0] ), 
	.D(n1062), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][15]  (.Q(\ram[26][15] ), 
	.D(n1013), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][14]  (.Q(\ram[26][14] ), 
	.D(n1012), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][13]  (.Q(\ram[26][13] ), 
	.D(n1011), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][12]  (.Q(\ram[26][12] ), 
	.D(n1010), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][11]  (.Q(\ram[26][11] ), 
	.D(n1009), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][10]  (.Q(\ram[26][10] ), 
	.D(n1008), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][9]  (.Q(\ram[26][9] ), 
	.D(n1007), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][8]  (.Q(\ram[26][8] ), 
	.D(n1006), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][7]  (.Q(\ram[26][7] ), 
	.D(n1005), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][6]  (.Q(\ram[26][6] ), 
	.D(n1004), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][5]  (.Q(\ram[26][5] ), 
	.D(n1003), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][4]  (.Q(\ram[26][4] ), 
	.D(n1002), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][3]  (.Q(\ram[26][3] ), 
	.D(n1001), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][2]  (.Q(\ram[26][2] ), 
	.D(n1000), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][1]  (.Q(\ram[26][1] ), 
	.D(n999), 
	.CK(clk));
   DFFHQX1 \ram_reg[26][0]  (.Q(\ram[26][0] ), 
	.D(n998), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][15]  (.Q(\ram[22][15] ), 
	.D(n949), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][14]  (.Q(\ram[22][14] ), 
	.D(n948), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][13]  (.Q(\ram[22][13] ), 
	.D(n947), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][12]  (.Q(\ram[22][12] ), 
	.D(n946), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][11]  (.Q(\ram[22][11] ), 
	.D(n945), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][10]  (.Q(\ram[22][10] ), 
	.D(n944), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][9]  (.Q(\ram[22][9] ), 
	.D(n943), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][8]  (.Q(\ram[22][8] ), 
	.D(n942), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][7]  (.Q(\ram[22][7] ), 
	.D(n941), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][6]  (.Q(\ram[22][6] ), 
	.D(n940), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][5]  (.Q(\ram[22][5] ), 
	.D(n939), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][4]  (.Q(\ram[22][4] ), 
	.D(n938), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][3]  (.Q(\ram[22][3] ), 
	.D(n937), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][2]  (.Q(\ram[22][2] ), 
	.D(n936), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][1]  (.Q(\ram[22][1] ), 
	.D(n935), 
	.CK(clk));
   DFFHQX1 \ram_reg[22][0]  (.Q(\ram[22][0] ), 
	.D(n934), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][15]  (.Q(\ram[18][15] ), 
	.D(n885), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][14]  (.Q(\ram[18][14] ), 
	.D(n884), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][13]  (.Q(\ram[18][13] ), 
	.D(n883), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][12]  (.Q(\ram[18][12] ), 
	.D(n882), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][11]  (.Q(\ram[18][11] ), 
	.D(n881), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][10]  (.Q(\ram[18][10] ), 
	.D(n880), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][9]  (.Q(\ram[18][9] ), 
	.D(n879), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][8]  (.Q(\ram[18][8] ), 
	.D(n878), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][7]  (.Q(\ram[18][7] ), 
	.D(n877), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][6]  (.Q(\ram[18][6] ), 
	.D(n876), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][5]  (.Q(\ram[18][5] ), 
	.D(n875), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][4]  (.Q(\ram[18][4] ), 
	.D(n874), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][3]  (.Q(\ram[18][3] ), 
	.D(n873), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][2]  (.Q(\ram[18][2] ), 
	.D(n872), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][1]  (.Q(\ram[18][1] ), 
	.D(n871), 
	.CK(clk));
   DFFHQX1 \ram_reg[18][0]  (.Q(\ram[18][0] ), 
	.D(n870), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][15]  (.Q(\ram[14][15] ), 
	.D(n821), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][14]  (.Q(\ram[14][14] ), 
	.D(n820), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][13]  (.Q(\ram[14][13] ), 
	.D(n819), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][12]  (.Q(\ram[14][12] ), 
	.D(n818), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][11]  (.Q(\ram[14][11] ), 
	.D(n817), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][10]  (.Q(\ram[14][10] ), 
	.D(n816), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][9]  (.Q(\ram[14][9] ), 
	.D(n815), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][8]  (.Q(\ram[14][8] ), 
	.D(n814), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][7]  (.Q(\ram[14][7] ), 
	.D(n813), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][6]  (.Q(\ram[14][6] ), 
	.D(n812), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][5]  (.Q(\ram[14][5] ), 
	.D(n811), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][4]  (.Q(\ram[14][4] ), 
	.D(n810), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][3]  (.Q(\ram[14][3] ), 
	.D(n809), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][2]  (.Q(\ram[14][2] ), 
	.D(n808), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][1]  (.Q(\ram[14][1] ), 
	.D(n807), 
	.CK(clk));
   DFFHQX1 \ram_reg[14][0]  (.Q(\ram[14][0] ), 
	.D(n806), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][15]  (.Q(\ram[10][15] ), 
	.D(n757), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][14]  (.Q(\ram[10][14] ), 
	.D(n756), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][13]  (.Q(\ram[10][13] ), 
	.D(n755), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][12]  (.Q(\ram[10][12] ), 
	.D(n754), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][11]  (.Q(\ram[10][11] ), 
	.D(n753), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][10]  (.Q(\ram[10][10] ), 
	.D(n752), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][9]  (.Q(\ram[10][9] ), 
	.D(n751), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][8]  (.Q(\ram[10][8] ), 
	.D(n750), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][7]  (.Q(\ram[10][7] ), 
	.D(n749), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][6]  (.Q(\ram[10][6] ), 
	.D(n748), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][5]  (.Q(\ram[10][5] ), 
	.D(n747), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][4]  (.Q(\ram[10][4] ), 
	.D(n746), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][3]  (.Q(\ram[10][3] ), 
	.D(n745), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][2]  (.Q(\ram[10][2] ), 
	.D(n744), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][1]  (.Q(\ram[10][1] ), 
	.D(n743), 
	.CK(clk));
   DFFHQX1 \ram_reg[10][0]  (.Q(\ram[10][0] ), 
	.D(n742), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][15]  (.Q(\ram[6][15] ), 
	.D(n693), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][14]  (.Q(\ram[6][14] ), 
	.D(n692), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][13]  (.Q(\ram[6][13] ), 
	.D(n691), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][12]  (.Q(\ram[6][12] ), 
	.D(n690), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][11]  (.Q(\ram[6][11] ), 
	.D(n689), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][10]  (.Q(\ram[6][10] ), 
	.D(n688), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][9]  (.Q(\ram[6][9] ), 
	.D(n687), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][8]  (.Q(\ram[6][8] ), 
	.D(n686), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][7]  (.Q(\ram[6][7] ), 
	.D(n685), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][6]  (.Q(\ram[6][6] ), 
	.D(n684), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][5]  (.Q(\ram[6][5] ), 
	.D(n683), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][4]  (.Q(\ram[6][4] ), 
	.D(n682), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][3]  (.Q(\ram[6][3] ), 
	.D(n681), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][2]  (.Q(\ram[6][2] ), 
	.D(n680), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][1]  (.Q(\ram[6][1] ), 
	.D(n679), 
	.CK(clk));
   DFFHQX1 \ram_reg[6][0]  (.Q(\ram[6][0] ), 
	.D(n678), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][15]  (.Q(\ram[2][15] ), 
	.D(n629), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][14]  (.Q(\ram[2][14] ), 
	.D(n628), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][13]  (.Q(\ram[2][13] ), 
	.D(n627), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][12]  (.Q(\ram[2][12] ), 
	.D(n626), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][11]  (.Q(\ram[2][11] ), 
	.D(n625), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][10]  (.Q(\ram[2][10] ), 
	.D(n624), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][9]  (.Q(\ram[2][9] ), 
	.D(n623), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][8]  (.Q(\ram[2][8] ), 
	.D(n622), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][7]  (.Q(\ram[2][7] ), 
	.D(n621), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][6]  (.Q(\ram[2][6] ), 
	.D(n620), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][5]  (.Q(\ram[2][5] ), 
	.D(n619), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][4]  (.Q(\ram[2][4] ), 
	.D(n618), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][3]  (.Q(\ram[2][3] ), 
	.D(n617), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][2]  (.Q(\ram[2][2] ), 
	.D(n616), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][1]  (.Q(\ram[2][1] ), 
	.D(n615), 
	.CK(clk));
   DFFHQX1 \ram_reg[2][0]  (.Q(\ram[2][0] ), 
	.D(n614), 
	.CK(clk));
   OAI22X1 U138 (.Y(n999), 
	.B1(n6307), 
	.B0(n6306), 
	.A1(n6305), 
	.A0(n6304));
   INVX1 U139 (.Y(n6305), 
	.A(\ram[26][1] ));
   OAI22X1 U140 (.Y(n998), 
	.B1(n6309), 
	.B0(n6307), 
	.A1(n6308), 
	.A0(n6304));
   INVX1 U141 (.Y(n6308), 
	.A(\ram[26][0] ));
   OAI22X1 U142 (.Y(n997), 
	.B1(n6313), 
	.B0(n6312), 
	.A1(n6311), 
	.A0(n6310));
   INVX1 U143 (.Y(n6313), 
	.A(\ram[25][15] ));
   OAI22X1 U144 (.Y(n996), 
	.B1(n6315), 
	.B0(n6312), 
	.A1(n6314), 
	.A0(n6310));
   INVX1 U145 (.Y(n6315), 
	.A(\ram[25][14] ));
   OAI22X1 U146 (.Y(n995), 
	.B1(n6317), 
	.B0(n6312), 
	.A1(n6316), 
	.A0(n6310));
   INVX1 U147 (.Y(n6317), 
	.A(\ram[25][13] ));
   OAI22X1 U148 (.Y(n994), 
	.B1(n6319), 
	.B0(n6312), 
	.A1(n6318), 
	.A0(n6310));
   INVX1 U149 (.Y(n6319), 
	.A(\ram[25][12] ));
   OAI22X1 U150 (.Y(n993), 
	.B1(n6321), 
	.B0(n6312), 
	.A1(n6320), 
	.A0(n6310));
   INVX1 U151 (.Y(n6321), 
	.A(\ram[25][11] ));
   OAI22X1 U152 (.Y(n992), 
	.B1(n6323), 
	.B0(n6312), 
	.A1(n6322), 
	.A0(n6310));
   INVX1 U153 (.Y(n6323), 
	.A(\ram[25][10] ));
   OAI22X1 U154 (.Y(n991), 
	.B1(n6325), 
	.B0(n6312), 
	.A1(n6324), 
	.A0(n6310));
   INVX1 U155 (.Y(n6325), 
	.A(\ram[25][9] ));
   OAI22X1 U156 (.Y(n990), 
	.B1(n6327), 
	.B0(n6312), 
	.A1(n6326), 
	.A0(n6310));
   INVX1 U157 (.Y(n6327), 
	.A(\ram[25][8] ));
   OAI22X1 U158 (.Y(n989), 
	.B1(n6329), 
	.B0(n6312), 
	.A1(n6328), 
	.A0(n6310));
   INVX1 U159 (.Y(n6329), 
	.A(\ram[25][7] ));
   OAI22X1 U160 (.Y(n988), 
	.B1(n6331), 
	.B0(n6312), 
	.A1(n6330), 
	.A0(n6310));
   INVX1 U161 (.Y(n6331), 
	.A(\ram[25][6] ));
   OAI22X1 U162 (.Y(n987), 
	.B1(n6333), 
	.B0(n6312), 
	.A1(n6332), 
	.A0(n6310));
   INVX1 U163 (.Y(n6333), 
	.A(\ram[25][5] ));
   OAI22X1 U164 (.Y(n986), 
	.B1(n6335), 
	.B0(n6312), 
	.A1(n6334), 
	.A0(n6310));
   INVX1 U165 (.Y(n6335), 
	.A(\ram[25][4] ));
   OAI22X1 U166 (.Y(n985), 
	.B1(n6337), 
	.B0(n6312), 
	.A1(n6336), 
	.A0(n6310));
   INVX1 U167 (.Y(n6337), 
	.A(\ram[25][3] ));
   OAI22X1 U168 (.Y(n984), 
	.B1(n6339), 
	.B0(n6312), 
	.A1(n6338), 
	.A0(n6310));
   INVX1 U169 (.Y(n6339), 
	.A(\ram[25][2] ));
   OAI22X1 U170 (.Y(n983), 
	.B1(n6340), 
	.B0(n6312), 
	.A1(n6310), 
	.A0(n6306));
   INVX1 U171 (.Y(n6340), 
	.A(\ram[25][1] ));
   OAI22X1 U172 (.Y(n982), 
	.B1(n6341), 
	.B0(n6312), 
	.A1(n6310), 
	.A0(n6309));
   INVX1 U173 (.Y(n6341), 
	.A(\ram[25][0] ));
   NOR2BX1 U174 (.Y(n6312), 
	.B(n6310), 
	.AN(mem_write_en));
   NAND2X1 U175 (.Y(n6310), 
	.B(n6343), 
	.A(n6342));
   OAI22X1 U176 (.Y(n981), 
	.B1(n6346), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6311));
   INVX1 U177 (.Y(n6346), 
	.A(\ram[24][15] ));
   OAI22X1 U178 (.Y(n980), 
	.B1(n6347), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6314));
   INVX1 U179 (.Y(n6347), 
	.A(\ram[24][14] ));
   OAI22X1 U180 (.Y(n979), 
	.B1(n6348), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6316));
   INVX1 U181 (.Y(n6348), 
	.A(\ram[24][13] ));
   OAI22X1 U182 (.Y(n978), 
	.B1(n6349), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6318));
   INVX1 U183 (.Y(n6349), 
	.A(\ram[24][12] ));
   OAI22X1 U184 (.Y(n977), 
	.B1(n6350), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6320));
   INVX1 U185 (.Y(n6350), 
	.A(\ram[24][11] ));
   OAI22X1 U186 (.Y(n976), 
	.B1(n6351), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6322));
   INVX1 U187 (.Y(n6351), 
	.A(\ram[24][10] ));
   OAI22X1 U188 (.Y(n975), 
	.B1(n6352), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6324));
   INVX1 U189 (.Y(n6352), 
	.A(\ram[24][9] ));
   OAI22X1 U190 (.Y(n974), 
	.B1(n6353), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6326));
   INVX1 U191 (.Y(n6353), 
	.A(\ram[24][8] ));
   OAI22X1 U192 (.Y(n973), 
	.B1(n6354), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6328));
   INVX1 U193 (.Y(n6354), 
	.A(\ram[24][7] ));
   OAI22X1 U194 (.Y(n972), 
	.B1(n6355), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6330));
   INVX1 U195 (.Y(n6355), 
	.A(\ram[24][6] ));
   OAI22X1 U196 (.Y(n971), 
	.B1(n6356), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6332));
   INVX1 U197 (.Y(n6356), 
	.A(\ram[24][5] ));
   OAI22X1 U198 (.Y(n970), 
	.B1(n6357), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6334));
   INVX1 U199 (.Y(n6357), 
	.A(\ram[24][4] ));
   OAI22X1 U200 (.Y(n969), 
	.B1(n6358), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6336));
   INVX1 U201 (.Y(n6358), 
	.A(\ram[24][3] ));
   OAI22X1 U202 (.Y(n968), 
	.B1(n6359), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6338));
   INVX1 U203 (.Y(n6359), 
	.A(\ram[24][2] ));
   OAI22X1 U204 (.Y(n967), 
	.B1(n6360), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6306));
   INVX1 U205 (.Y(n6360), 
	.A(\ram[24][1] ));
   OAI22X1 U206 (.Y(n966), 
	.B1(n6361), 
	.B0(n6345), 
	.A1(n6344), 
	.A0(n6309));
   INVX1 U207 (.Y(n6361), 
	.A(\ram[24][0] ));
   NOR2BX1 U208 (.Y(n6345), 
	.B(n6344), 
	.AN(mem_write_en));
   NAND2X1 U209 (.Y(n6344), 
	.B(n6343), 
	.A(n6362));
   OAI22X1 U210 (.Y(n965), 
	.B1(n6365), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6311));
   INVX1 U211 (.Y(n6365), 
	.A(\ram[23][15] ));
   OAI22X1 U212 (.Y(n964), 
	.B1(n6366), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6314));
   INVX1 U213 (.Y(n6366), 
	.A(\ram[23][14] ));
   OAI22X1 U214 (.Y(n963), 
	.B1(n6367), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6316));
   INVX1 U215 (.Y(n6367), 
	.A(\ram[23][13] ));
   OAI22X1 U216 (.Y(n962), 
	.B1(n6368), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6318));
   INVX1 U217 (.Y(n6368), 
	.A(\ram[23][12] ));
   OAI22X1 U218 (.Y(n961), 
	.B1(n6369), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6320));
   INVX1 U219 (.Y(n6369), 
	.A(\ram[23][11] ));
   OAI22X1 U220 (.Y(n960), 
	.B1(n6370), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6322));
   INVX1 U221 (.Y(n6370), 
	.A(\ram[23][10] ));
   OAI22X1 U222 (.Y(n959), 
	.B1(n6371), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6324));
   INVX1 U223 (.Y(n6371), 
	.A(\ram[23][9] ));
   OAI22X1 U224 (.Y(n958), 
	.B1(n6372), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6326));
   INVX1 U225 (.Y(n6372), 
	.A(\ram[23][8] ));
   OAI22X1 U226 (.Y(n957), 
	.B1(n6373), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6328));
   INVX1 U227 (.Y(n6373), 
	.A(\ram[23][7] ));
   OAI22X1 U228 (.Y(n956), 
	.B1(n6374), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6330));
   INVX1 U229 (.Y(n6374), 
	.A(\ram[23][6] ));
   OAI22X1 U230 (.Y(n955), 
	.B1(n6375), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6332));
   INVX1 U231 (.Y(n6375), 
	.A(\ram[23][5] ));
   OAI22X1 U232 (.Y(n954), 
	.B1(n6376), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6334));
   INVX1 U233 (.Y(n6376), 
	.A(\ram[23][4] ));
   OAI22X1 U234 (.Y(n953), 
	.B1(n6377), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6336));
   INVX1 U235 (.Y(n6377), 
	.A(\ram[23][3] ));
   OAI22X1 U236 (.Y(n952), 
	.B1(n6378), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6338));
   INVX1 U237 (.Y(n6378), 
	.A(\ram[23][2] ));
   OAI22X1 U238 (.Y(n951), 
	.B1(n6379), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6306));
   INVX1 U239 (.Y(n6379), 
	.A(\ram[23][1] ));
   OAI22X1 U240 (.Y(n950), 
	.B1(n6380), 
	.B0(n6364), 
	.A1(n6363), 
	.A0(n6309));
   INVX1 U241 (.Y(n6380), 
	.A(\ram[23][0] ));
   NOR2BX1 U242 (.Y(n6364), 
	.B(n6363), 
	.AN(mem_write_en));
   NAND2X1 U243 (.Y(n6363), 
	.B(n6343), 
	.A(n6381));
   OAI22X1 U244 (.Y(n949), 
	.B1(n6384), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6311));
   INVX1 U245 (.Y(n6384), 
	.A(\ram[22][15] ));
   OAI22X1 U246 (.Y(n948), 
	.B1(n6385), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6314));
   INVX1 U247 (.Y(n6385), 
	.A(\ram[22][14] ));
   OAI22X1 U248 (.Y(n947), 
	.B1(n6386), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6316));
   INVX1 U249 (.Y(n6386), 
	.A(\ram[22][13] ));
   OAI22X1 U250 (.Y(n946), 
	.B1(n6387), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6318));
   INVX1 U251 (.Y(n6387), 
	.A(\ram[22][12] ));
   OAI22X1 U252 (.Y(n945), 
	.B1(n6388), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6320));
   INVX1 U253 (.Y(n6388), 
	.A(\ram[22][11] ));
   OAI22X1 U254 (.Y(n944), 
	.B1(n6389), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6322));
   INVX1 U255 (.Y(n6389), 
	.A(\ram[22][10] ));
   OAI22X1 U256 (.Y(n943), 
	.B1(n6390), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6324));
   INVX1 U257 (.Y(n6390), 
	.A(\ram[22][9] ));
   OAI22X1 U258 (.Y(n942), 
	.B1(n6391), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6326));
   INVX1 U259 (.Y(n6391), 
	.A(\ram[22][8] ));
   OAI22X1 U260 (.Y(n941), 
	.B1(n6392), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6328));
   INVX1 U261 (.Y(n6392), 
	.A(\ram[22][7] ));
   OAI22X1 U262 (.Y(n940), 
	.B1(n6393), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6330));
   INVX1 U263 (.Y(n6393), 
	.A(\ram[22][6] ));
   OAI22X1 U264 (.Y(n939), 
	.B1(n6394), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6332));
   INVX1 U265 (.Y(n6394), 
	.A(\ram[22][5] ));
   OAI22X1 U266 (.Y(n938), 
	.B1(n6395), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6334));
   INVX1 U267 (.Y(n6395), 
	.A(\ram[22][4] ));
   OAI22X1 U268 (.Y(n937), 
	.B1(n6396), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6336));
   INVX1 U269 (.Y(n6396), 
	.A(\ram[22][3] ));
   OAI22X1 U270 (.Y(n936), 
	.B1(n6397), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6338));
   INVX1 U271 (.Y(n6397), 
	.A(\ram[22][2] ));
   OAI22X1 U272 (.Y(n935), 
	.B1(n6398), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6306));
   INVX1 U273 (.Y(n6398), 
	.A(\ram[22][1] ));
   OAI22X1 U274 (.Y(n934), 
	.B1(n6399), 
	.B0(n6383), 
	.A1(n6382), 
	.A0(n6309));
   INVX1 U275 (.Y(n6399), 
	.A(\ram[22][0] ));
   NOR2BX1 U276 (.Y(n6383), 
	.B(n6382), 
	.AN(mem_write_en));
   NAND2X1 U277 (.Y(n6382), 
	.B(n6343), 
	.A(n6400));
   OAI22X1 U278 (.Y(n933), 
	.B1(n6403), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6311));
   INVX1 U279 (.Y(n6403), 
	.A(\ram[21][15] ));
   OAI22X1 U280 (.Y(n932), 
	.B1(n6404), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6314));
   INVX1 U281 (.Y(n6404), 
	.A(\ram[21][14] ));
   OAI22X1 U282 (.Y(n931), 
	.B1(n6405), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6316));
   INVX1 U283 (.Y(n6405), 
	.A(\ram[21][13] ));
   OAI22X1 U284 (.Y(n930), 
	.B1(n6406), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6318));
   INVX1 U285 (.Y(n6406), 
	.A(\ram[21][12] ));
   OAI22X1 U286 (.Y(n929), 
	.B1(n6407), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6320));
   INVX1 U287 (.Y(n6407), 
	.A(\ram[21][11] ));
   OAI22X1 U288 (.Y(n928), 
	.B1(n6408), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6322));
   INVX1 U289 (.Y(n6408), 
	.A(\ram[21][10] ));
   OAI22X1 U290 (.Y(n927), 
	.B1(n6409), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6324));
   INVX1 U291 (.Y(n6409), 
	.A(\ram[21][9] ));
   OAI22X1 U292 (.Y(n926), 
	.B1(n6410), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6326));
   INVX1 U293 (.Y(n6410), 
	.A(\ram[21][8] ));
   OAI22X1 U294 (.Y(n925), 
	.B1(n6411), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6328));
   INVX1 U295 (.Y(n6411), 
	.A(\ram[21][7] ));
   OAI22X1 U296 (.Y(n924), 
	.B1(n6412), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6330));
   INVX1 U297 (.Y(n6412), 
	.A(\ram[21][6] ));
   OAI22X1 U298 (.Y(n923), 
	.B1(n6413), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6332));
   INVX1 U299 (.Y(n6413), 
	.A(\ram[21][5] ));
   OAI22X1 U300 (.Y(n922), 
	.B1(n6414), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6334));
   INVX1 U301 (.Y(n6414), 
	.A(\ram[21][4] ));
   OAI22X1 U302 (.Y(n921), 
	.B1(n6415), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6336));
   INVX1 U303 (.Y(n6415), 
	.A(\ram[21][3] ));
   OAI22X1 U304 (.Y(n920), 
	.B1(n6416), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6338));
   INVX1 U305 (.Y(n6416), 
	.A(\ram[21][2] ));
   OAI22X1 U306 (.Y(n919), 
	.B1(n6417), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6306));
   INVX1 U307 (.Y(n6417), 
	.A(\ram[21][1] ));
   OAI22X1 U308 (.Y(n918), 
	.B1(n6418), 
	.B0(n6402), 
	.A1(n6401), 
	.A0(n6309));
   INVX1 U309 (.Y(n6418), 
	.A(\ram[21][0] ));
   NOR2BX1 U310 (.Y(n6402), 
	.B(n6401), 
	.AN(mem_write_en));
   NAND2X1 U311 (.Y(n6401), 
	.B(n6343), 
	.A(n6419));
   OAI22X1 U312 (.Y(n917), 
	.B1(n6422), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6311));
   INVX1 U313 (.Y(n6422), 
	.A(\ram[20][15] ));
   OAI22X1 U314 (.Y(n916), 
	.B1(n6423), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6314));
   INVX1 U315 (.Y(n6423), 
	.A(\ram[20][14] ));
   OAI22X1 U316 (.Y(n915), 
	.B1(n6424), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6316));
   INVX1 U317 (.Y(n6424), 
	.A(\ram[20][13] ));
   OAI22X1 U318 (.Y(n914), 
	.B1(n6425), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6318));
   INVX1 U319 (.Y(n6425), 
	.A(\ram[20][12] ));
   OAI22X1 U320 (.Y(n913), 
	.B1(n6426), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6320));
   INVX1 U321 (.Y(n6426), 
	.A(\ram[20][11] ));
   OAI22X1 U322 (.Y(n912), 
	.B1(n6427), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6322));
   INVX1 U323 (.Y(n6427), 
	.A(\ram[20][10] ));
   OAI22X1 U324 (.Y(n911), 
	.B1(n6428), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6324));
   INVX1 U325 (.Y(n6428), 
	.A(\ram[20][9] ));
   OAI22X1 U326 (.Y(n910), 
	.B1(n6429), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6326));
   INVX1 U327 (.Y(n6429), 
	.A(\ram[20][8] ));
   OAI22X1 U328 (.Y(n909), 
	.B1(n6430), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6328));
   INVX1 U329 (.Y(n6430), 
	.A(\ram[20][7] ));
   OAI22X1 U330 (.Y(n908), 
	.B1(n6431), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6330));
   INVX1 U331 (.Y(n6431), 
	.A(\ram[20][6] ));
   OAI22X1 U332 (.Y(n907), 
	.B1(n6432), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6332));
   INVX1 U333 (.Y(n6432), 
	.A(\ram[20][5] ));
   OAI22X1 U334 (.Y(n906), 
	.B1(n6433), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6334));
   INVX1 U335 (.Y(n6433), 
	.A(\ram[20][4] ));
   OAI22X1 U336 (.Y(n905), 
	.B1(n6434), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6336));
   INVX1 U337 (.Y(n6434), 
	.A(\ram[20][3] ));
   OAI22X1 U338 (.Y(n904), 
	.B1(n6435), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6338));
   INVX1 U339 (.Y(n6435), 
	.A(\ram[20][2] ));
   OAI22X1 U340 (.Y(n903), 
	.B1(n6436), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6306));
   INVX1 U341 (.Y(n6436), 
	.A(\ram[20][1] ));
   OAI22X1 U342 (.Y(n902), 
	.B1(n6437), 
	.B0(n6421), 
	.A1(n6420), 
	.A0(n6309));
   INVX1 U343 (.Y(n6437), 
	.A(\ram[20][0] ));
   NOR2BX1 U344 (.Y(n6421), 
	.B(n6420), 
	.AN(mem_write_en));
   NAND2X1 U345 (.Y(n6420), 
	.B(n6343), 
	.A(n6438));
   OAI22X1 U346 (.Y(n901), 
	.B1(n6441), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6311));
   INVX1 U347 (.Y(n6441), 
	.A(\ram[19][15] ));
   OAI22X1 U348 (.Y(n900), 
	.B1(n6442), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6314));
   INVX1 U349 (.Y(n6442), 
	.A(\ram[19][14] ));
   OAI22X1 U350 (.Y(n899), 
	.B1(n6443), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6316));
   INVX1 U351 (.Y(n6443), 
	.A(\ram[19][13] ));
   OAI22X1 U352 (.Y(n898), 
	.B1(n6444), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6318));
   INVX1 U353 (.Y(n6444), 
	.A(\ram[19][12] ));
   OAI22X1 U354 (.Y(n897), 
	.B1(n6445), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6320));
   INVX1 U355 (.Y(n6445), 
	.A(\ram[19][11] ));
   OAI22X1 U356 (.Y(n896), 
	.B1(n6446), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6322));
   INVX1 U357 (.Y(n6446), 
	.A(\ram[19][10] ));
   OAI22X1 U358 (.Y(n895), 
	.B1(n6447), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6324));
   INVX1 U359 (.Y(n6447), 
	.A(\ram[19][9] ));
   OAI22X1 U360 (.Y(n894), 
	.B1(n6448), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6326));
   INVX1 U361 (.Y(n6448), 
	.A(\ram[19][8] ));
   OAI22X1 U362 (.Y(n893), 
	.B1(n6449), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6328));
   INVX1 U363 (.Y(n6449), 
	.A(\ram[19][7] ));
   OAI22X1 U364 (.Y(n892), 
	.B1(n6450), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6330));
   INVX1 U365 (.Y(n6450), 
	.A(\ram[19][6] ));
   OAI22X1 U366 (.Y(n891), 
	.B1(n6451), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6332));
   INVX1 U367 (.Y(n6451), 
	.A(\ram[19][5] ));
   OAI22X1 U368 (.Y(n890), 
	.B1(n6452), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6334));
   INVX1 U369 (.Y(n6452), 
	.A(\ram[19][4] ));
   OAI22X1 U370 (.Y(n889), 
	.B1(n6453), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6336));
   INVX1 U371 (.Y(n6453), 
	.A(\ram[19][3] ));
   OAI22X1 U372 (.Y(n888), 
	.B1(n6454), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6338));
   INVX1 U373 (.Y(n6454), 
	.A(\ram[19][2] ));
   OAI22X1 U374 (.Y(n887), 
	.B1(n6455), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6306));
   INVX1 U375 (.Y(n6455), 
	.A(\ram[19][1] ));
   OAI22X1 U376 (.Y(n886), 
	.B1(n6456), 
	.B0(n6440), 
	.A1(n6439), 
	.A0(n6309));
   INVX1 U377 (.Y(n6456), 
	.A(\ram[19][0] ));
   NOR2BX1 U378 (.Y(n6440), 
	.B(n6439), 
	.AN(mem_write_en));
   NAND2X1 U379 (.Y(n6439), 
	.B(n6343), 
	.A(n6457));
   OAI22X1 U380 (.Y(n885), 
	.B1(n6460), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6311));
   INVX1 U381 (.Y(n6460), 
	.A(\ram[18][15] ));
   OAI22X1 U382 (.Y(n884), 
	.B1(n6461), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6314));
   INVX1 U383 (.Y(n6461), 
	.A(\ram[18][14] ));
   OAI22X1 U384 (.Y(n883), 
	.B1(n6462), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6316));
   INVX1 U385 (.Y(n6462), 
	.A(\ram[18][13] ));
   OAI22X1 U386 (.Y(n882), 
	.B1(n6463), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6318));
   INVX1 U387 (.Y(n6463), 
	.A(\ram[18][12] ));
   OAI22X1 U388 (.Y(n881), 
	.B1(n6464), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6320));
   INVX1 U389 (.Y(n6464), 
	.A(\ram[18][11] ));
   OAI22X1 U390 (.Y(n880), 
	.B1(n6465), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6322));
   INVX1 U391 (.Y(n6465), 
	.A(\ram[18][10] ));
   OAI22X1 U392 (.Y(n879), 
	.B1(n6466), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6324));
   INVX1 U393 (.Y(n6466), 
	.A(\ram[18][9] ));
   OAI22X1 U394 (.Y(n878), 
	.B1(n6467), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6326));
   INVX1 U395 (.Y(n6467), 
	.A(\ram[18][8] ));
   OAI22X1 U396 (.Y(n877), 
	.B1(n6468), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6328));
   INVX1 U397 (.Y(n6468), 
	.A(\ram[18][7] ));
   OAI22X1 U398 (.Y(n876), 
	.B1(n6469), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6330));
   INVX1 U399 (.Y(n6469), 
	.A(\ram[18][6] ));
   OAI22X1 U400 (.Y(n875), 
	.B1(n6470), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6332));
   INVX1 U401 (.Y(n6470), 
	.A(\ram[18][5] ));
   OAI22X1 U402 (.Y(n874), 
	.B1(n6471), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6334));
   INVX1 U403 (.Y(n6471), 
	.A(\ram[18][4] ));
   OAI22X1 U404 (.Y(n873), 
	.B1(n6472), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6336));
   INVX1 U405 (.Y(n6472), 
	.A(\ram[18][3] ));
   OAI22X1 U406 (.Y(n872), 
	.B1(n6473), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6338));
   INVX1 U407 (.Y(n6473), 
	.A(\ram[18][2] ));
   OAI22X1 U408 (.Y(n871), 
	.B1(n6474), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6306));
   INVX1 U409 (.Y(n6474), 
	.A(\ram[18][1] ));
   OAI22X1 U410 (.Y(n870), 
	.B1(n6475), 
	.B0(n6459), 
	.A1(n6458), 
	.A0(n6309));
   INVX1 U411 (.Y(n6475), 
	.A(\ram[18][0] ));
   NOR2BX1 U412 (.Y(n6459), 
	.B(n6458), 
	.AN(mem_write_en));
   NAND2X1 U413 (.Y(n6458), 
	.B(n6343), 
	.A(n6476));
   OAI22X1 U414 (.Y(n869), 
	.B1(n6479), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6311));
   INVX1 U415 (.Y(n6479), 
	.A(\ram[17][15] ));
   OAI22X1 U416 (.Y(n868), 
	.B1(n6480), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6314));
   INVX1 U417 (.Y(n6480), 
	.A(\ram[17][14] ));
   OAI22X1 U418 (.Y(n867), 
	.B1(n6481), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6316));
   INVX1 U419 (.Y(n6481), 
	.A(\ram[17][13] ));
   OAI22X1 U420 (.Y(n866), 
	.B1(n6482), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6318));
   INVX1 U421 (.Y(n6482), 
	.A(\ram[17][12] ));
   OAI22X1 U422 (.Y(n865), 
	.B1(n6483), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6320));
   INVX1 U423 (.Y(n6483), 
	.A(\ram[17][11] ));
   OAI22X1 U424 (.Y(n864), 
	.B1(n6484), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6322));
   INVX1 U425 (.Y(n6484), 
	.A(\ram[17][10] ));
   OAI22X1 U426 (.Y(n863), 
	.B1(n6485), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6324));
   INVX1 U427 (.Y(n6485), 
	.A(\ram[17][9] ));
   OAI22X1 U428 (.Y(n862), 
	.B1(n6486), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6326));
   INVX1 U429 (.Y(n6486), 
	.A(\ram[17][8] ));
   OAI22X1 U430 (.Y(n861), 
	.B1(n6487), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6328));
   INVX1 U431 (.Y(n6487), 
	.A(\ram[17][7] ));
   OAI22X1 U432 (.Y(n860), 
	.B1(n6488), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6330));
   INVX1 U433 (.Y(n6488), 
	.A(\ram[17][6] ));
   OAI22X1 U434 (.Y(n859), 
	.B1(n6489), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6332));
   INVX1 U435 (.Y(n6489), 
	.A(\ram[17][5] ));
   OAI22X1 U436 (.Y(n858), 
	.B1(n6490), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6334));
   INVX1 U437 (.Y(n6490), 
	.A(\ram[17][4] ));
   OAI22X1 U438 (.Y(n857), 
	.B1(n6491), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6336));
   INVX1 U439 (.Y(n6491), 
	.A(\ram[17][3] ));
   OAI22X1 U440 (.Y(n856), 
	.B1(n6492), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6338));
   INVX1 U441 (.Y(n6492), 
	.A(\ram[17][2] ));
   OAI22X1 U442 (.Y(n855), 
	.B1(n6493), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6306));
   INVX1 U443 (.Y(n6493), 
	.A(\ram[17][1] ));
   OAI22X1 U444 (.Y(n854), 
	.B1(n6494), 
	.B0(n6478), 
	.A1(n6477), 
	.A0(n6309));
   INVX1 U445 (.Y(n6494), 
	.A(\ram[17][0] ));
   NOR2BX1 U446 (.Y(n6478), 
	.B(n6477), 
	.AN(mem_write_en));
   NAND2X1 U447 (.Y(n6477), 
	.B(n6343), 
	.A(n6495));
   OAI22X1 U448 (.Y(n853), 
	.B1(n6498), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6311));
   INVX1 U449 (.Y(n6498), 
	.A(\ram[16][15] ));
   OAI22X1 U450 (.Y(n852), 
	.B1(n6499), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6314));
   INVX1 U451 (.Y(n6499), 
	.A(\ram[16][14] ));
   OAI22X1 U452 (.Y(n851), 
	.B1(n6500), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6316));
   INVX1 U453 (.Y(n6500), 
	.A(\ram[16][13] ));
   OAI22X1 U454 (.Y(n850), 
	.B1(n6501), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6318));
   INVX1 U455 (.Y(n6501), 
	.A(\ram[16][12] ));
   OAI22X1 U456 (.Y(n849), 
	.B1(n6502), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6320));
   INVX1 U457 (.Y(n6502), 
	.A(\ram[16][11] ));
   OAI22X1 U458 (.Y(n848), 
	.B1(n6503), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6322));
   INVX1 U459 (.Y(n6503), 
	.A(\ram[16][10] ));
   OAI22X1 U460 (.Y(n847), 
	.B1(n6504), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6324));
   INVX1 U461 (.Y(n6504), 
	.A(\ram[16][9] ));
   OAI22X1 U462 (.Y(n846), 
	.B1(n6505), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6326));
   INVX1 U463 (.Y(n6505), 
	.A(\ram[16][8] ));
   OAI22X1 U464 (.Y(n845), 
	.B1(n6506), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6328));
   INVX1 U465 (.Y(n6506), 
	.A(\ram[16][7] ));
   OAI22X1 U466 (.Y(n844), 
	.B1(n6507), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6330));
   INVX1 U467 (.Y(n6507), 
	.A(\ram[16][6] ));
   OAI22X1 U468 (.Y(n843), 
	.B1(n6508), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6332));
   INVX1 U469 (.Y(n6508), 
	.A(\ram[16][5] ));
   OAI22X1 U470 (.Y(n842), 
	.B1(n6509), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6334));
   INVX1 U471 (.Y(n6509), 
	.A(\ram[16][4] ));
   OAI22X1 U472 (.Y(n841), 
	.B1(n6510), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6336));
   INVX1 U473 (.Y(n6510), 
	.A(\ram[16][3] ));
   OAI22X1 U474 (.Y(n840), 
	.B1(n6511), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6338));
   INVX1 U475 (.Y(n6511), 
	.A(\ram[16][2] ));
   OAI22X1 U476 (.Y(n839), 
	.B1(n6512), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6306));
   INVX1 U477 (.Y(n6512), 
	.A(\ram[16][1] ));
   OAI22X1 U478 (.Y(n838), 
	.B1(n6513), 
	.B0(n6497), 
	.A1(n6496), 
	.A0(n6309));
   INVX1 U479 (.Y(n6513), 
	.A(\ram[16][0] ));
   NOR2BX1 U480 (.Y(n6497), 
	.B(n6496), 
	.AN(mem_write_en));
   NAND2X1 U481 (.Y(n6496), 
	.B(n6343), 
	.A(n6514));
   OAI22X1 U482 (.Y(n837), 
	.B1(n6517), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6311));
   INVX1 U483 (.Y(n6517), 
	.A(\ram[15][15] ));
   OAI22X1 U484 (.Y(n836), 
	.B1(n6518), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6314));
   INVX1 U485 (.Y(n6518), 
	.A(\ram[15][14] ));
   OAI22X1 U486 (.Y(n835), 
	.B1(n6519), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6316));
   INVX1 U487 (.Y(n6519), 
	.A(\ram[15][13] ));
   OAI22X1 U488 (.Y(n834), 
	.B1(n6520), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6318));
   INVX1 U489 (.Y(n6520), 
	.A(\ram[15][12] ));
   OAI22X1 U490 (.Y(n833), 
	.B1(n6521), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6320));
   INVX1 U491 (.Y(n6521), 
	.A(\ram[15][11] ));
   OAI22X1 U492 (.Y(n832), 
	.B1(n6522), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6322));
   INVX1 U493 (.Y(n6522), 
	.A(\ram[15][10] ));
   OAI22X1 U494 (.Y(n831), 
	.B1(n6523), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6324));
   INVX1 U495 (.Y(n6523), 
	.A(\ram[15][9] ));
   OAI22X1 U496 (.Y(n830), 
	.B1(n6524), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6326));
   INVX1 U497 (.Y(n6524), 
	.A(\ram[15][8] ));
   OAI22X1 U498 (.Y(n829), 
	.B1(n6525), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6328));
   INVX1 U499 (.Y(n6525), 
	.A(\ram[15][7] ));
   OAI22X1 U500 (.Y(n828), 
	.B1(n6526), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6330));
   INVX1 U501 (.Y(n6526), 
	.A(\ram[15][6] ));
   OAI22X1 U502 (.Y(n827), 
	.B1(n6527), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6332));
   INVX1 U503 (.Y(n6527), 
	.A(\ram[15][5] ));
   OAI22X1 U504 (.Y(n826), 
	.B1(n6528), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6334));
   INVX1 U505 (.Y(n6528), 
	.A(\ram[15][4] ));
   OAI22X1 U506 (.Y(n825), 
	.B1(n6529), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6336));
   INVX1 U507 (.Y(n6529), 
	.A(\ram[15][3] ));
   OAI22X1 U508 (.Y(n824), 
	.B1(n6530), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6338));
   INVX1 U509 (.Y(n6530), 
	.A(\ram[15][2] ));
   OAI22X1 U510 (.Y(n823), 
	.B1(n6531), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6306));
   INVX1 U511 (.Y(n6531), 
	.A(\ram[15][1] ));
   OAI22X1 U512 (.Y(n822), 
	.B1(n6532), 
	.B0(n6516), 
	.A1(n6515), 
	.A0(n6309));
   INVX1 U513 (.Y(n6532), 
	.A(\ram[15][0] ));
   NOR2BX1 U514 (.Y(n6516), 
	.B(n6515), 
	.AN(mem_write_en));
   NAND2X1 U515 (.Y(n6515), 
	.B(n6534), 
	.A(n6533));
   OAI22X1 U516 (.Y(n821), 
	.B1(n6537), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6311));
   INVX1 U517 (.Y(n6537), 
	.A(\ram[14][15] ));
   OAI22X1 U518 (.Y(n820), 
	.B1(n6538), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6314));
   INVX1 U519 (.Y(n6538), 
	.A(\ram[14][14] ));
   OAI22X1 U520 (.Y(n819), 
	.B1(n6539), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6316));
   INVX1 U521 (.Y(n6539), 
	.A(\ram[14][13] ));
   OAI22X1 U522 (.Y(n818), 
	.B1(n6540), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6318));
   INVX1 U523 (.Y(n6540), 
	.A(\ram[14][12] ));
   OAI22X1 U524 (.Y(n817), 
	.B1(n6541), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6320));
   INVX1 U525 (.Y(n6541), 
	.A(\ram[14][11] ));
   OAI22X1 U526 (.Y(n816), 
	.B1(n6542), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6322));
   INVX1 U527 (.Y(n6542), 
	.A(\ram[14][10] ));
   OAI22X1 U528 (.Y(n815), 
	.B1(n6543), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6324));
   INVX1 U529 (.Y(n6543), 
	.A(\ram[14][9] ));
   OAI22X1 U530 (.Y(n814), 
	.B1(n6544), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6326));
   INVX1 U531 (.Y(n6544), 
	.A(\ram[14][8] ));
   OAI22X1 U532 (.Y(n813), 
	.B1(n6545), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6328));
   INVX1 U533 (.Y(n6545), 
	.A(\ram[14][7] ));
   OAI22X1 U534 (.Y(n812), 
	.B1(n6546), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6330));
   INVX1 U535 (.Y(n6546), 
	.A(\ram[14][6] ));
   OAI22X1 U536 (.Y(n811), 
	.B1(n6547), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6332));
   INVX1 U537 (.Y(n6547), 
	.A(\ram[14][5] ));
   OAI22X1 U538 (.Y(n810), 
	.B1(n6548), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6334));
   INVX1 U539 (.Y(n6548), 
	.A(\ram[14][4] ));
   OAI22X1 U540 (.Y(n809), 
	.B1(n6549), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6336));
   INVX1 U541 (.Y(n6549), 
	.A(\ram[14][3] ));
   OAI22X1 U542 (.Y(n808), 
	.B1(n6550), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6338));
   INVX1 U543 (.Y(n6550), 
	.A(\ram[14][2] ));
   OAI22X1 U544 (.Y(n807), 
	.B1(n6551), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6306));
   INVX1 U545 (.Y(n6551), 
	.A(\ram[14][1] ));
   OAI22X1 U546 (.Y(n806), 
	.B1(n6552), 
	.B0(n6536), 
	.A1(n6535), 
	.A0(n6309));
   INVX1 U547 (.Y(n6552), 
	.A(\ram[14][0] ));
   NOR2BX1 U548 (.Y(n6536), 
	.B(n6535), 
	.AN(mem_write_en));
   NAND2X1 U549 (.Y(n6535), 
	.B(n6534), 
	.A(n6553));
   OAI22X1 U550 (.Y(n805), 
	.B1(n6556), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6311));
   INVX1 U551 (.Y(n6556), 
	.A(\ram[13][15] ));
   OAI22X1 U552 (.Y(n804), 
	.B1(n6557), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6314));
   INVX1 U553 (.Y(n6557), 
	.A(\ram[13][14] ));
   OAI22X1 U554 (.Y(n803), 
	.B1(n6558), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6316));
   INVX1 U555 (.Y(n6558), 
	.A(\ram[13][13] ));
   OAI22X1 U556 (.Y(n802), 
	.B1(n6559), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6318));
   INVX1 U557 (.Y(n6559), 
	.A(\ram[13][12] ));
   OAI22X1 U558 (.Y(n801), 
	.B1(n6560), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6320));
   INVX1 U559 (.Y(n6560), 
	.A(\ram[13][11] ));
   OAI22X1 U560 (.Y(n800), 
	.B1(n6561), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6322));
   INVX1 U561 (.Y(n6561), 
	.A(\ram[13][10] ));
   OAI22X1 U562 (.Y(n799), 
	.B1(n6562), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6324));
   INVX1 U563 (.Y(n6562), 
	.A(\ram[13][9] ));
   OAI22X1 U564 (.Y(n798), 
	.B1(n6563), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6326));
   INVX1 U565 (.Y(n6563), 
	.A(\ram[13][8] ));
   OAI22X1 U566 (.Y(n797), 
	.B1(n6564), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6328));
   INVX1 U567 (.Y(n6564), 
	.A(\ram[13][7] ));
   OAI22X1 U568 (.Y(n796), 
	.B1(n6565), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6330));
   INVX1 U569 (.Y(n6565), 
	.A(\ram[13][6] ));
   OAI22X1 U570 (.Y(n795), 
	.B1(n6566), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6332));
   INVX1 U571 (.Y(n6566), 
	.A(\ram[13][5] ));
   OAI22X1 U572 (.Y(n794), 
	.B1(n6567), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6334));
   INVX1 U573 (.Y(n6567), 
	.A(\ram[13][4] ));
   OAI22X1 U574 (.Y(n793), 
	.B1(n6568), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6336));
   INVX1 U575 (.Y(n6568), 
	.A(\ram[13][3] ));
   OAI22X1 U576 (.Y(n792), 
	.B1(n6569), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6338));
   INVX1 U577 (.Y(n6569), 
	.A(\ram[13][2] ));
   OAI22X1 U578 (.Y(n791), 
	.B1(n6570), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6306));
   INVX1 U579 (.Y(n6570), 
	.A(\ram[13][1] ));
   OAI22X1 U580 (.Y(n790), 
	.B1(n6571), 
	.B0(n6555), 
	.A1(n6554), 
	.A0(n6309));
   INVX1 U581 (.Y(n6571), 
	.A(\ram[13][0] ));
   NOR2BX1 U582 (.Y(n6555), 
	.B(n6554), 
	.AN(mem_write_en));
   NAND2X1 U583 (.Y(n6554), 
	.B(n6534), 
	.A(n6572));
   OAI22X1 U584 (.Y(n789), 
	.B1(n6575), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6311));
   INVX1 U585 (.Y(n6575), 
	.A(\ram[12][15] ));
   OAI22X1 U586 (.Y(n788), 
	.B1(n6576), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6314));
   INVX1 U587 (.Y(n6576), 
	.A(\ram[12][14] ));
   OAI22X1 U588 (.Y(n787), 
	.B1(n6577), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6316));
   INVX1 U589 (.Y(n6577), 
	.A(\ram[12][13] ));
   OAI22X1 U590 (.Y(n786), 
	.B1(n6578), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6318));
   INVX1 U591 (.Y(n6578), 
	.A(\ram[12][12] ));
   OAI22X1 U592 (.Y(n785), 
	.B1(n6579), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6320));
   INVX1 U593 (.Y(n6579), 
	.A(\ram[12][11] ));
   OAI22X1 U594 (.Y(n784), 
	.B1(n6580), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6322));
   INVX1 U595 (.Y(n6580), 
	.A(\ram[12][10] ));
   OAI22X1 U596 (.Y(n783), 
	.B1(n6581), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6324));
   INVX1 U597 (.Y(n6581), 
	.A(\ram[12][9] ));
   OAI22X1 U598 (.Y(n782), 
	.B1(n6582), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6326));
   INVX1 U599 (.Y(n6582), 
	.A(\ram[12][8] ));
   OAI22X1 U600 (.Y(n781), 
	.B1(n6583), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6328));
   INVX1 U601 (.Y(n6583), 
	.A(\ram[12][7] ));
   OAI22X1 U602 (.Y(n780), 
	.B1(n6584), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6330));
   INVX1 U603 (.Y(n6584), 
	.A(\ram[12][6] ));
   OAI22X1 U604 (.Y(n779), 
	.B1(n6585), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6332));
   INVX1 U605 (.Y(n6585), 
	.A(\ram[12][5] ));
   OAI22X1 U606 (.Y(n778), 
	.B1(n6586), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6334));
   INVX1 U607 (.Y(n6586), 
	.A(\ram[12][4] ));
   OAI22X1 U608 (.Y(n777), 
	.B1(n6587), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6336));
   INVX1 U609 (.Y(n6587), 
	.A(\ram[12][3] ));
   OAI22X1 U610 (.Y(n776), 
	.B1(n6588), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6338));
   INVX1 U611 (.Y(n6588), 
	.A(\ram[12][2] ));
   OAI22X1 U612 (.Y(n775), 
	.B1(n6589), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6306));
   INVX1 U613 (.Y(n6589), 
	.A(\ram[12][1] ));
   OAI22X1 U614 (.Y(n774), 
	.B1(n6590), 
	.B0(n6574), 
	.A1(n6573), 
	.A0(n6309));
   INVX1 U615 (.Y(n6590), 
	.A(\ram[12][0] ));
   NOR2BX1 U616 (.Y(n6574), 
	.B(n6573), 
	.AN(mem_write_en));
   NAND2X1 U617 (.Y(n6573), 
	.B(n6534), 
	.A(n6591));
   OAI22X1 U618 (.Y(n773), 
	.B1(n6594), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6311));
   INVX1 U619 (.Y(n6594), 
	.A(\ram[11][15] ));
   OAI22X1 U620 (.Y(n772), 
	.B1(n6595), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6314));
   INVX1 U621 (.Y(n6595), 
	.A(\ram[11][14] ));
   OAI22X1 U622 (.Y(n771), 
	.B1(n6596), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6316));
   INVX1 U623 (.Y(n6596), 
	.A(\ram[11][13] ));
   OAI22X1 U624 (.Y(n770), 
	.B1(n6597), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6318));
   INVX1 U625 (.Y(n6597), 
	.A(\ram[11][12] ));
   OAI22X1 U626 (.Y(n769), 
	.B1(n6598), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6320));
   INVX1 U627 (.Y(n6598), 
	.A(\ram[11][11] ));
   OAI22X1 U628 (.Y(n768), 
	.B1(n6599), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6322));
   INVX1 U629 (.Y(n6599), 
	.A(\ram[11][10] ));
   OAI22X1 U630 (.Y(n767), 
	.B1(n6600), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6324));
   INVX1 U631 (.Y(n6600), 
	.A(\ram[11][9] ));
   OAI22X1 U632 (.Y(n766), 
	.B1(n6601), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6326));
   INVX1 U633 (.Y(n6601), 
	.A(\ram[11][8] ));
   OAI22X1 U634 (.Y(n765), 
	.B1(n6602), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6328));
   INVX1 U635 (.Y(n6602), 
	.A(\ram[11][7] ));
   OAI22X1 U636 (.Y(n764), 
	.B1(n6603), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6330));
   INVX1 U637 (.Y(n6603), 
	.A(\ram[11][6] ));
   OAI22X1 U638 (.Y(n763), 
	.B1(n6604), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6332));
   INVX1 U639 (.Y(n6604), 
	.A(\ram[11][5] ));
   OAI22X1 U640 (.Y(n762), 
	.B1(n6605), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6334));
   INVX1 U641 (.Y(n6605), 
	.A(\ram[11][4] ));
   OAI22X1 U642 (.Y(n761), 
	.B1(n6606), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6336));
   INVX1 U643 (.Y(n6606), 
	.A(\ram[11][3] ));
   OAI22X1 U644 (.Y(n760), 
	.B1(n6607), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6338));
   INVX1 U645 (.Y(n6607), 
	.A(\ram[11][2] ));
   OAI22X1 U646 (.Y(n759), 
	.B1(n6608), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6306));
   INVX1 U647 (.Y(n6608), 
	.A(\ram[11][1] ));
   OAI22X1 U648 (.Y(n758), 
	.B1(n6609), 
	.B0(n6593), 
	.A1(n6592), 
	.A0(n6309));
   INVX1 U649 (.Y(n6609), 
	.A(\ram[11][0] ));
   NOR2BX1 U650 (.Y(n6593), 
	.B(n6592), 
	.AN(mem_write_en));
   NAND2X1 U651 (.Y(n6592), 
	.B(n6534), 
	.A(n6610));
   OAI22X1 U652 (.Y(n757), 
	.B1(n6613), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6311));
   INVX1 U653 (.Y(n6613), 
	.A(\ram[10][15] ));
   OAI22X1 U654 (.Y(n756), 
	.B1(n6614), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6314));
   INVX1 U655 (.Y(n6614), 
	.A(\ram[10][14] ));
   OAI22X1 U656 (.Y(n755), 
	.B1(n6615), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6316));
   INVX1 U657 (.Y(n6615), 
	.A(\ram[10][13] ));
   OAI22X1 U658 (.Y(n754), 
	.B1(n6616), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6318));
   INVX1 U659 (.Y(n6616), 
	.A(\ram[10][12] ));
   OAI22X1 U660 (.Y(n753), 
	.B1(n6617), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6320));
   INVX1 U661 (.Y(n6617), 
	.A(\ram[10][11] ));
   OAI22X1 U662 (.Y(n752), 
	.B1(n6618), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6322));
   INVX1 U663 (.Y(n6618), 
	.A(\ram[10][10] ));
   OAI22X1 U664 (.Y(n751), 
	.B1(n6619), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6324));
   INVX1 U665 (.Y(n6619), 
	.A(\ram[10][9] ));
   OAI22X1 U666 (.Y(n750), 
	.B1(n6620), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6326));
   INVX1 U667 (.Y(n6620), 
	.A(\ram[10][8] ));
   OAI22X1 U668 (.Y(n749), 
	.B1(n6621), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6328));
   INVX1 U669 (.Y(n6621), 
	.A(\ram[10][7] ));
   OAI22X1 U670 (.Y(n748), 
	.B1(n6622), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6330));
   INVX1 U671 (.Y(n6622), 
	.A(\ram[10][6] ));
   OAI22X1 U672 (.Y(n747), 
	.B1(n6623), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6332));
   INVX1 U673 (.Y(n6623), 
	.A(\ram[10][5] ));
   OAI22X1 U674 (.Y(n746), 
	.B1(n6624), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6334));
   INVX1 U675 (.Y(n6624), 
	.A(\ram[10][4] ));
   OAI22X1 U676 (.Y(n745), 
	.B1(n6625), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6336));
   INVX1 U677 (.Y(n6625), 
	.A(\ram[10][3] ));
   OAI22X1 U678 (.Y(n744), 
	.B1(n6626), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6338));
   INVX1 U679 (.Y(n6626), 
	.A(\ram[10][2] ));
   OAI22X1 U680 (.Y(n743), 
	.B1(n6627), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6306));
   INVX1 U681 (.Y(n6627), 
	.A(\ram[10][1] ));
   OAI22X1 U682 (.Y(n742), 
	.B1(n6628), 
	.B0(n6612), 
	.A1(n6611), 
	.A0(n6309));
   INVX1 U683 (.Y(n6628), 
	.A(\ram[10][0] ));
   NOR2BX1 U684 (.Y(n6612), 
	.B(n6611), 
	.AN(mem_write_en));
   NAND2X1 U685 (.Y(n6611), 
	.B(n6629), 
	.A(n6534));
   OAI22X1 U686 (.Y(n741), 
	.B1(n6632), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6311));
   INVX1 U687 (.Y(n6632), 
	.A(\ram[9][15] ));
   OAI22X1 U688 (.Y(n740), 
	.B1(n6633), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6314));
   INVX1 U689 (.Y(n6633), 
	.A(\ram[9][14] ));
   OAI22X1 U690 (.Y(n739), 
	.B1(n6634), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6316));
   INVX1 U691 (.Y(n6634), 
	.A(\ram[9][13] ));
   OAI22X1 U692 (.Y(n738), 
	.B1(n6635), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6318));
   INVX1 U693 (.Y(n6635), 
	.A(\ram[9][12] ));
   OAI22X1 U694 (.Y(n737), 
	.B1(n6636), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6320));
   INVX1 U695 (.Y(n6636), 
	.A(\ram[9][11] ));
   OAI22X1 U696 (.Y(n736), 
	.B1(n6637), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6322));
   INVX1 U697 (.Y(n6637), 
	.A(\ram[9][10] ));
   OAI22X1 U698 (.Y(n735), 
	.B1(n6638), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6324));
   INVX1 U699 (.Y(n6638), 
	.A(\ram[9][9] ));
   OAI22X1 U700 (.Y(n734), 
	.B1(n6639), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6326));
   INVX1 U701 (.Y(n6639), 
	.A(\ram[9][8] ));
   OAI22X1 U702 (.Y(n733), 
	.B1(n6640), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6328));
   INVX1 U703 (.Y(n6640), 
	.A(\ram[9][7] ));
   OAI22X1 U704 (.Y(n732), 
	.B1(n6641), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6330));
   INVX1 U705 (.Y(n6641), 
	.A(\ram[9][6] ));
   OAI22X1 U706 (.Y(n731), 
	.B1(n6642), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6332));
   INVX1 U707 (.Y(n6642), 
	.A(\ram[9][5] ));
   OAI22X1 U708 (.Y(n730), 
	.B1(n6643), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6334));
   INVX1 U709 (.Y(n6643), 
	.A(\ram[9][4] ));
   OAI22X1 U710 (.Y(n729), 
	.B1(n6644), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6336));
   INVX1 U711 (.Y(n6644), 
	.A(\ram[9][3] ));
   OAI22X1 U712 (.Y(n728), 
	.B1(n6645), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6338));
   INVX1 U713 (.Y(n6645), 
	.A(\ram[9][2] ));
   OAI22X1 U714 (.Y(n727), 
	.B1(n6646), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6306));
   INVX1 U715 (.Y(n6646), 
	.A(\ram[9][1] ));
   OAI22X1 U716 (.Y(n726), 
	.B1(n6647), 
	.B0(n6631), 
	.A1(n6630), 
	.A0(n6309));
   INVX1 U717 (.Y(n6647), 
	.A(\ram[9][0] ));
   NOR2BX1 U718 (.Y(n6631), 
	.B(n6630), 
	.AN(mem_write_en));
   NAND2X1 U719 (.Y(n6630), 
	.B(n6342), 
	.A(n6534));
   OAI22X1 U720 (.Y(n725), 
	.B1(n6650), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6311));
   INVX1 U721 (.Y(n6650), 
	.A(\ram[8][15] ));
   OAI22X1 U722 (.Y(n724), 
	.B1(n6651), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6314));
   INVX1 U723 (.Y(n6651), 
	.A(\ram[8][14] ));
   OAI22X1 U724 (.Y(n723), 
	.B1(n6652), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6316));
   INVX1 U725 (.Y(n6652), 
	.A(\ram[8][13] ));
   OAI22X1 U726 (.Y(n722), 
	.B1(n6653), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6318));
   INVX1 U727 (.Y(n6653), 
	.A(\ram[8][12] ));
   OAI22X1 U728 (.Y(n721), 
	.B1(n6654), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6320));
   INVX1 U729 (.Y(n6654), 
	.A(\ram[8][11] ));
   OAI22X1 U730 (.Y(n720), 
	.B1(n6655), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6322));
   INVX1 U731 (.Y(n6655), 
	.A(\ram[8][10] ));
   OAI22X1 U732 (.Y(n719), 
	.B1(n6656), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6324));
   INVX1 U733 (.Y(n6656), 
	.A(\ram[8][9] ));
   OAI22X1 U734 (.Y(n718), 
	.B1(n6657), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6326));
   INVX1 U735 (.Y(n6657), 
	.A(\ram[8][8] ));
   OAI22X1 U736 (.Y(n717), 
	.B1(n6658), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6328));
   INVX1 U737 (.Y(n6658), 
	.A(\ram[8][7] ));
   OAI22X1 U738 (.Y(n716), 
	.B1(n6659), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6330));
   INVX1 U739 (.Y(n6659), 
	.A(\ram[8][6] ));
   OAI22X1 U740 (.Y(n715), 
	.B1(n6660), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6332));
   INVX1 U741 (.Y(n6660), 
	.A(\ram[8][5] ));
   OAI22X1 U742 (.Y(n714), 
	.B1(n6661), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6334));
   INVX1 U743 (.Y(n6661), 
	.A(\ram[8][4] ));
   OAI22X1 U744 (.Y(n713), 
	.B1(n6662), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6336));
   INVX1 U745 (.Y(n6662), 
	.A(\ram[8][3] ));
   OAI22X1 U746 (.Y(n712), 
	.B1(n6663), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6338));
   INVX1 U747 (.Y(n6663), 
	.A(\ram[8][2] ));
   OAI22X1 U748 (.Y(n711), 
	.B1(n6664), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6306));
   INVX1 U749 (.Y(n6664), 
	.A(\ram[8][1] ));
   OAI22X1 U750 (.Y(n710), 
	.B1(n6665), 
	.B0(n6649), 
	.A1(n6648), 
	.A0(n6309));
   INVX1 U751 (.Y(n6665), 
	.A(\ram[8][0] ));
   NOR2BX1 U752 (.Y(n6649), 
	.B(n6648), 
	.AN(mem_write_en));
   NAND2X1 U753 (.Y(n6648), 
	.B(n6362), 
	.A(n6534));
   OAI22X1 U754 (.Y(n709), 
	.B1(n6668), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6311));
   INVX1 U755 (.Y(n6668), 
	.A(\ram[7][15] ));
   OAI22X1 U756 (.Y(n708), 
	.B1(n6669), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6314));
   INVX1 U757 (.Y(n6669), 
	.A(\ram[7][14] ));
   OAI22X1 U758 (.Y(n707), 
	.B1(n6670), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6316));
   INVX1 U759 (.Y(n6670), 
	.A(\ram[7][13] ));
   OAI22X1 U760 (.Y(n706), 
	.B1(n6671), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6318));
   INVX1 U761 (.Y(n6671), 
	.A(\ram[7][12] ));
   OAI22X1 U762 (.Y(n705), 
	.B1(n6672), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6320));
   INVX1 U763 (.Y(n6672), 
	.A(\ram[7][11] ));
   OAI22X1 U764 (.Y(n704), 
	.B1(n6673), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6322));
   INVX1 U765 (.Y(n6673), 
	.A(\ram[7][10] ));
   OAI22X1 U766 (.Y(n703), 
	.B1(n6674), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6324));
   INVX1 U767 (.Y(n6674), 
	.A(\ram[7][9] ));
   OAI22X1 U768 (.Y(n702), 
	.B1(n6675), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6326));
   INVX1 U769 (.Y(n6675), 
	.A(\ram[7][8] ));
   OAI22X1 U770 (.Y(n701), 
	.B1(n6676), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6328));
   INVX1 U771 (.Y(n6676), 
	.A(\ram[7][7] ));
   OAI22X1 U772 (.Y(n700), 
	.B1(n6677), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6330));
   INVX1 U773 (.Y(n6677), 
	.A(\ram[7][6] ));
   OAI22X1 U774 (.Y(n699), 
	.B1(n6678), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6332));
   INVX1 U775 (.Y(n6678), 
	.A(\ram[7][5] ));
   OAI22X1 U776 (.Y(n698), 
	.B1(n6679), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6334));
   INVX1 U777 (.Y(n6679), 
	.A(\ram[7][4] ));
   OAI22X1 U778 (.Y(n697), 
	.B1(n6680), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6336));
   INVX1 U779 (.Y(n6680), 
	.A(\ram[7][3] ));
   OAI22X1 U780 (.Y(n696), 
	.B1(n6681), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6338));
   INVX1 U781 (.Y(n6681), 
	.A(\ram[7][2] ));
   OAI22X1 U782 (.Y(n695), 
	.B1(n6682), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6306));
   INVX1 U783 (.Y(n6682), 
	.A(\ram[7][1] ));
   OAI22X1 U784 (.Y(n694), 
	.B1(n6683), 
	.B0(n6667), 
	.A1(n6666), 
	.A0(n6309));
   INVX1 U785 (.Y(n6683), 
	.A(\ram[7][0] ));
   NOR2BX1 U786 (.Y(n6667), 
	.B(n6666), 
	.AN(mem_write_en));
   NAND2X1 U787 (.Y(n6666), 
	.B(n6381), 
	.A(n6534));
   OAI22X1 U788 (.Y(n693), 
	.B1(n6686), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6311));
   INVX1 U789 (.Y(n6686), 
	.A(\ram[6][15] ));
   OAI22X1 U790 (.Y(n692), 
	.B1(n6687), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6314));
   INVX1 U791 (.Y(n6687), 
	.A(\ram[6][14] ));
   OAI22X1 U792 (.Y(n691), 
	.B1(n6688), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6316));
   INVX1 U793 (.Y(n6688), 
	.A(\ram[6][13] ));
   OAI22X1 U794 (.Y(n690), 
	.B1(n6689), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6318));
   INVX1 U795 (.Y(n6689), 
	.A(\ram[6][12] ));
   OAI22X1 U796 (.Y(n689), 
	.B1(n6690), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6320));
   INVX1 U797 (.Y(n6690), 
	.A(\ram[6][11] ));
   OAI22X1 U798 (.Y(n688), 
	.B1(n6691), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6322));
   INVX1 U799 (.Y(n6691), 
	.A(\ram[6][10] ));
   OAI22X1 U800 (.Y(n687), 
	.B1(n6692), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6324));
   INVX1 U801 (.Y(n6692), 
	.A(\ram[6][9] ));
   OAI22X1 U802 (.Y(n686), 
	.B1(n6693), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6326));
   INVX1 U803 (.Y(n6693), 
	.A(\ram[6][8] ));
   OAI22X1 U804 (.Y(n685), 
	.B1(n6694), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6328));
   INVX1 U805 (.Y(n6694), 
	.A(\ram[6][7] ));
   OAI22X1 U806 (.Y(n684), 
	.B1(n6695), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6330));
   INVX1 U807 (.Y(n6695), 
	.A(\ram[6][6] ));
   OAI22X1 U808 (.Y(n683), 
	.B1(n6696), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6332));
   INVX1 U809 (.Y(n6696), 
	.A(\ram[6][5] ));
   OAI22X1 U810 (.Y(n682), 
	.B1(n6697), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6334));
   INVX1 U811 (.Y(n6697), 
	.A(\ram[6][4] ));
   OAI22X1 U812 (.Y(n681), 
	.B1(n6698), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6336));
   INVX1 U813 (.Y(n6698), 
	.A(\ram[6][3] ));
   OAI22X1 U814 (.Y(n680), 
	.B1(n6699), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6338));
   INVX1 U815 (.Y(n6699), 
	.A(\ram[6][2] ));
   OAI22X1 U816 (.Y(n679), 
	.B1(n6700), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6306));
   INVX1 U817 (.Y(n6700), 
	.A(\ram[6][1] ));
   OAI22X1 U818 (.Y(n678), 
	.B1(n6701), 
	.B0(n6685), 
	.A1(n6684), 
	.A0(n6309));
   INVX1 U819 (.Y(n6701), 
	.A(\ram[6][0] ));
   NOR2BX1 U820 (.Y(n6685), 
	.B(n6684), 
	.AN(mem_write_en));
   NAND2X1 U821 (.Y(n6684), 
	.B(n6400), 
	.A(n6534));
   OAI22X1 U822 (.Y(n677), 
	.B1(n6704), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6311));
   INVX1 U823 (.Y(n6704), 
	.A(\ram[5][15] ));
   OAI22X1 U824 (.Y(n676), 
	.B1(n6705), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6314));
   INVX1 U825 (.Y(n6705), 
	.A(\ram[5][14] ));
   OAI22X1 U826 (.Y(n675), 
	.B1(n6706), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6316));
   INVX1 U827 (.Y(n6706), 
	.A(\ram[5][13] ));
   OAI22X1 U828 (.Y(n674), 
	.B1(n6707), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6318));
   INVX1 U829 (.Y(n6707), 
	.A(\ram[5][12] ));
   OAI22X1 U830 (.Y(n673), 
	.B1(n6708), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6320));
   INVX1 U831 (.Y(n6708), 
	.A(\ram[5][11] ));
   OAI22X1 U832 (.Y(n672), 
	.B1(n6709), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6322));
   INVX1 U833 (.Y(n6709), 
	.A(\ram[5][10] ));
   OAI22X1 U834 (.Y(n671), 
	.B1(n6710), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6324));
   INVX1 U835 (.Y(n6710), 
	.A(\ram[5][9] ));
   OAI22X1 U836 (.Y(n670), 
	.B1(n6711), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6326));
   INVX1 U837 (.Y(n6711), 
	.A(\ram[5][8] ));
   OAI22X1 U838 (.Y(n669), 
	.B1(n6712), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6328));
   INVX1 U839 (.Y(n6712), 
	.A(\ram[5][7] ));
   OAI22X1 U840 (.Y(n668), 
	.B1(n6713), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6330));
   INVX1 U841 (.Y(n6713), 
	.A(\ram[5][6] ));
   OAI22X1 U842 (.Y(n667), 
	.B1(n6714), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6332));
   INVX1 U843 (.Y(n6714), 
	.A(\ram[5][5] ));
   OAI22X1 U844 (.Y(n666), 
	.B1(n6715), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6334));
   INVX1 U845 (.Y(n6715), 
	.A(\ram[5][4] ));
   OAI22X1 U846 (.Y(n665), 
	.B1(n6716), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6336));
   INVX1 U847 (.Y(n6716), 
	.A(\ram[5][3] ));
   OAI22X1 U848 (.Y(n664), 
	.B1(n6717), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6338));
   INVX1 U849 (.Y(n6717), 
	.A(\ram[5][2] ));
   OAI22X1 U850 (.Y(n663), 
	.B1(n6718), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6306));
   INVX1 U851 (.Y(n6718), 
	.A(\ram[5][1] ));
   OAI22X1 U852 (.Y(n662), 
	.B1(n6719), 
	.B0(n6703), 
	.A1(n6702), 
	.A0(n6309));
   INVX1 U853 (.Y(n6719), 
	.A(\ram[5][0] ));
   NOR2BX1 U854 (.Y(n6703), 
	.B(n6702), 
	.AN(mem_write_en));
   NAND2X1 U855 (.Y(n6702), 
	.B(n6419), 
	.A(n6534));
   OAI22X1 U856 (.Y(n661), 
	.B1(n6722), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6311));
   INVX1 U857 (.Y(n6722), 
	.A(\ram[4][15] ));
   OAI22X1 U858 (.Y(n660), 
	.B1(n6723), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6314));
   INVX1 U859 (.Y(n6723), 
	.A(\ram[4][14] ));
   OAI22X1 U860 (.Y(n659), 
	.B1(n6724), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6316));
   INVX1 U861 (.Y(n6724), 
	.A(\ram[4][13] ));
   OAI22X1 U862 (.Y(n658), 
	.B1(n6725), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6318));
   INVX1 U863 (.Y(n6725), 
	.A(\ram[4][12] ));
   OAI22X1 U864 (.Y(n657), 
	.B1(n6726), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6320));
   INVX1 U865 (.Y(n6726), 
	.A(\ram[4][11] ));
   OAI22X1 U866 (.Y(n656), 
	.B1(n6727), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6322));
   INVX1 U867 (.Y(n6727), 
	.A(\ram[4][10] ));
   OAI22X1 U868 (.Y(n655), 
	.B1(n6728), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6324));
   INVX1 U869 (.Y(n6728), 
	.A(\ram[4][9] ));
   OAI22X1 U870 (.Y(n654), 
	.B1(n6729), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6326));
   INVX1 U871 (.Y(n6729), 
	.A(\ram[4][8] ));
   OAI22X1 U872 (.Y(n653), 
	.B1(n6730), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6328));
   INVX1 U873 (.Y(n6730), 
	.A(\ram[4][7] ));
   OAI22X1 U874 (.Y(n652), 
	.B1(n6731), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6330));
   INVX1 U875 (.Y(n6731), 
	.A(\ram[4][6] ));
   OAI22X1 U876 (.Y(n651), 
	.B1(n6732), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6332));
   INVX1 U877 (.Y(n6732), 
	.A(\ram[4][5] ));
   OAI22X1 U878 (.Y(n650), 
	.B1(n6733), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6334));
   INVX1 U879 (.Y(n6733), 
	.A(\ram[4][4] ));
   OAI22X1 U880 (.Y(n649), 
	.B1(n6734), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6336));
   INVX1 U881 (.Y(n6734), 
	.A(\ram[4][3] ));
   OAI22X1 U882 (.Y(n648), 
	.B1(n6735), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6338));
   INVX1 U883 (.Y(n6735), 
	.A(\ram[4][2] ));
   OAI22X1 U884 (.Y(n647), 
	.B1(n6736), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6306));
   INVX1 U885 (.Y(n6736), 
	.A(\ram[4][1] ));
   OAI22X1 U886 (.Y(n646), 
	.B1(n6737), 
	.B0(n6721), 
	.A1(n6720), 
	.A0(n6309));
   INVX1 U887 (.Y(n6737), 
	.A(\ram[4][0] ));
   NOR2BX1 U888 (.Y(n6721), 
	.B(n6720), 
	.AN(mem_write_en));
   NAND2X1 U889 (.Y(n6720), 
	.B(n6438), 
	.A(n6534));
   OAI22X1 U890 (.Y(n645), 
	.B1(n6740), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6311));
   INVX1 U891 (.Y(n6740), 
	.A(\ram[3][15] ));
   OAI22X1 U892 (.Y(n644), 
	.B1(n6741), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6314));
   INVX1 U893 (.Y(n6741), 
	.A(\ram[3][14] ));
   OAI22X1 U894 (.Y(n643), 
	.B1(n6742), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6316));
   INVX1 U895 (.Y(n6742), 
	.A(\ram[3][13] ));
   OAI22X1 U896 (.Y(n642), 
	.B1(n6743), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6318));
   INVX1 U897 (.Y(n6743), 
	.A(\ram[3][12] ));
   OAI22X1 U898 (.Y(n641), 
	.B1(n6744), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6320));
   INVX1 U899 (.Y(n6744), 
	.A(\ram[3][11] ));
   OAI22X1 U900 (.Y(n640), 
	.B1(n6745), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6322));
   INVX1 U901 (.Y(n6745), 
	.A(\ram[3][10] ));
   OAI22X1 U902 (.Y(n639), 
	.B1(n6746), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6324));
   INVX1 U903 (.Y(n6746), 
	.A(\ram[3][9] ));
   OAI22X1 U904 (.Y(n638), 
	.B1(n6747), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6326));
   INVX1 U905 (.Y(n6747), 
	.A(\ram[3][8] ));
   OAI22X1 U906 (.Y(n637), 
	.B1(n6748), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6328));
   INVX1 U907 (.Y(n6748), 
	.A(\ram[3][7] ));
   OAI22X1 U908 (.Y(n636), 
	.B1(n6749), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6330));
   INVX1 U909 (.Y(n6749), 
	.A(\ram[3][6] ));
   OAI22X1 U910 (.Y(n635), 
	.B1(n6750), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6332));
   INVX1 U911 (.Y(n6750), 
	.A(\ram[3][5] ));
   OAI22X1 U912 (.Y(n634), 
	.B1(n6751), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6334));
   INVX1 U913 (.Y(n6751), 
	.A(\ram[3][4] ));
   OAI22X1 U914 (.Y(n633), 
	.B1(n6752), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6336));
   INVX1 U915 (.Y(n6752), 
	.A(\ram[3][3] ));
   OAI22X1 U916 (.Y(n632), 
	.B1(n6753), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6338));
   INVX1 U917 (.Y(n6753), 
	.A(\ram[3][2] ));
   OAI22X1 U918 (.Y(n631), 
	.B1(n6754), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6306));
   INVX1 U919 (.Y(n6754), 
	.A(\ram[3][1] ));
   OAI22X1 U920 (.Y(n630), 
	.B1(n6755), 
	.B0(n6739), 
	.A1(n6738), 
	.A0(n6309));
   INVX1 U921 (.Y(n6755), 
	.A(\ram[3][0] ));
   NOR2BX1 U922 (.Y(n6739), 
	.B(n6738), 
	.AN(mem_write_en));
   NAND2X1 U923 (.Y(n6738), 
	.B(n6457), 
	.A(n6534));
   OAI22X1 U924 (.Y(n629), 
	.B1(n6758), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6311));
   INVX1 U925 (.Y(n6758), 
	.A(\ram[2][15] ));
   OAI22X1 U926 (.Y(n628), 
	.B1(n6759), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6314));
   INVX1 U927 (.Y(n6759), 
	.A(\ram[2][14] ));
   OAI22X1 U928 (.Y(n627), 
	.B1(n6760), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6316));
   INVX1 U929 (.Y(n6760), 
	.A(\ram[2][13] ));
   OAI22X1 U930 (.Y(n626), 
	.B1(n6761), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6318));
   INVX1 U931 (.Y(n6761), 
	.A(\ram[2][12] ));
   OAI22X1 U932 (.Y(n625), 
	.B1(n6762), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6320));
   INVX1 U933 (.Y(n6762), 
	.A(\ram[2][11] ));
   OAI22X1 U934 (.Y(n624), 
	.B1(n6763), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6322));
   INVX1 U935 (.Y(n6763), 
	.A(\ram[2][10] ));
   OAI22X1 U936 (.Y(n623), 
	.B1(n6764), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6324));
   INVX1 U937 (.Y(n6764), 
	.A(\ram[2][9] ));
   OAI22X1 U938 (.Y(n622), 
	.B1(n6765), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6326));
   INVX1 U939 (.Y(n6765), 
	.A(\ram[2][8] ));
   OAI22X1 U940 (.Y(n621), 
	.B1(n6766), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6328));
   INVX1 U941 (.Y(n6766), 
	.A(\ram[2][7] ));
   OAI22X1 U942 (.Y(n620), 
	.B1(n6767), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6330));
   INVX1 U943 (.Y(n6767), 
	.A(\ram[2][6] ));
   OAI22X1 U944 (.Y(n619), 
	.B1(n6768), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6332));
   INVX1 U945 (.Y(n6768), 
	.A(\ram[2][5] ));
   OAI22X1 U946 (.Y(n618), 
	.B1(n6769), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6334));
   INVX1 U947 (.Y(n6769), 
	.A(\ram[2][4] ));
   OAI22X1 U948 (.Y(n617), 
	.B1(n6770), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6336));
   INVX1 U949 (.Y(n6770), 
	.A(\ram[2][3] ));
   OAI22X1 U950 (.Y(n616), 
	.B1(n6771), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6338));
   INVX1 U951 (.Y(n6771), 
	.A(\ram[2][2] ));
   OAI22X1 U952 (.Y(n615), 
	.B1(n6772), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6306));
   INVX1 U953 (.Y(n6772), 
	.A(\ram[2][1] ));
   OAI22X1 U954 (.Y(n614), 
	.B1(n6773), 
	.B0(n6757), 
	.A1(n6756), 
	.A0(n6309));
   INVX1 U955 (.Y(n6773), 
	.A(\ram[2][0] ));
   NOR2BX1 U956 (.Y(n6757), 
	.B(n6756), 
	.AN(mem_write_en));
   NAND2X1 U957 (.Y(n6756), 
	.B(n6476), 
	.A(n6534));
   OAI22X1 U958 (.Y(n613), 
	.B1(n6776), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6311));
   INVX1 U959 (.Y(n6776), 
	.A(\ram[1][15] ));
   OAI22X1 U960 (.Y(n612), 
	.B1(n6777), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6314));
   INVX1 U961 (.Y(n6777), 
	.A(\ram[1][14] ));
   OAI22X1 U962 (.Y(n611), 
	.B1(n6778), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6316));
   INVX1 U963 (.Y(n6778), 
	.A(\ram[1][13] ));
   OAI22X1 U964 (.Y(n610), 
	.B1(n6779), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6318));
   INVX1 U965 (.Y(n6779), 
	.A(\ram[1][12] ));
   OAI22X1 U966 (.Y(n609), 
	.B1(n6780), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6320));
   INVX1 U967 (.Y(n6780), 
	.A(\ram[1][11] ));
   OAI22X1 U968 (.Y(n608), 
	.B1(n6781), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6322));
   INVX1 U969 (.Y(n6781), 
	.A(\ram[1][10] ));
   OAI22X1 U970 (.Y(n607), 
	.B1(n6782), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6324));
   INVX1 U971 (.Y(n6782), 
	.A(\ram[1][9] ));
   OAI22X1 U972 (.Y(n606), 
	.B1(n6783), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6326));
   INVX1 U973 (.Y(n6783), 
	.A(\ram[1][8] ));
   OAI22X1 U974 (.Y(n605), 
	.B1(n6784), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6328));
   INVX1 U975 (.Y(n6784), 
	.A(\ram[1][7] ));
   OAI22X1 U976 (.Y(n604), 
	.B1(n6785), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6330));
   INVX1 U977 (.Y(n6785), 
	.A(\ram[1][6] ));
   OAI22X1 U978 (.Y(n603), 
	.B1(n6786), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6332));
   INVX1 U979 (.Y(n6786), 
	.A(\ram[1][5] ));
   OAI22X1 U980 (.Y(n602), 
	.B1(n6787), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6334));
   INVX1 U981 (.Y(n6787), 
	.A(\ram[1][4] ));
   OAI22X1 U982 (.Y(n601), 
	.B1(n6788), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6336));
   INVX1 U983 (.Y(n6788), 
	.A(\ram[1][3] ));
   OAI22X1 U984 (.Y(n600), 
	.B1(n6789), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6338));
   INVX1 U985 (.Y(n6789), 
	.A(\ram[1][2] ));
   OAI22X1 U986 (.Y(n599), 
	.B1(n6790), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6306));
   INVX1 U987 (.Y(n6790), 
	.A(\ram[1][1] ));
   OAI22X1 U988 (.Y(n598), 
	.B1(n6791), 
	.B0(n6775), 
	.A1(n6774), 
	.A0(n6309));
   INVX1 U989 (.Y(n6791), 
	.A(\ram[1][0] ));
   NOR2BX1 U990 (.Y(n6775), 
	.B(n6774), 
	.AN(mem_write_en));
   NAND2X1 U991 (.Y(n6774), 
	.B(n6495), 
	.A(n6534));
   OAI22X1 U992 (.Y(n597), 
	.B1(n6794), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6311));
   INVX1 U993 (.Y(n6794), 
	.A(\ram[0][15] ));
   OAI22X1 U994 (.Y(n596), 
	.B1(n6795), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6314));
   INVX1 U995 (.Y(n6795), 
	.A(\ram[0][14] ));
   OAI22X1 U996 (.Y(n595), 
	.B1(n6796), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6316));
   INVX1 U997 (.Y(n6796), 
	.A(\ram[0][13] ));
   OAI22X1 U998 (.Y(n594), 
	.B1(n6797), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6318));
   INVX1 U999 (.Y(n6797), 
	.A(\ram[0][12] ));
   OAI22X1 U1000 (.Y(n593), 
	.B1(n6798), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6320));
   INVX1 U1001 (.Y(n6798), 
	.A(\ram[0][11] ));
   OAI22X1 U1002 (.Y(n592), 
	.B1(n6799), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6322));
   INVX1 U1003 (.Y(n6799), 
	.A(\ram[0][10] ));
   OAI22X1 U1004 (.Y(n591), 
	.B1(n6800), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6324));
   INVX1 U1005 (.Y(n6800), 
	.A(\ram[0][9] ));
   OAI22X1 U1006 (.Y(n590), 
	.B1(n6801), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6326));
   INVX1 U1007 (.Y(n6801), 
	.A(\ram[0][8] ));
   OAI22X1 U1008 (.Y(n589), 
	.B1(n6802), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6328));
   INVX1 U1009 (.Y(n6802), 
	.A(\ram[0][7] ));
   OAI22X1 U1010 (.Y(n588), 
	.B1(n6803), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6330));
   INVX1 U1011 (.Y(n6803), 
	.A(\ram[0][6] ));
   OAI22X1 U1012 (.Y(n587), 
	.B1(n6804), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6332));
   INVX1 U1013 (.Y(n6804), 
	.A(\ram[0][5] ));
   OAI22X1 U1014 (.Y(n586), 
	.B1(n6805), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6334));
   INVX1 U1015 (.Y(n6805), 
	.A(\ram[0][4] ));
   OAI22X1 U1016 (.Y(n585), 
	.B1(n6806), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6336));
   INVX1 U1017 (.Y(n6806), 
	.A(\ram[0][3] ));
   OAI22X1 U1018 (.Y(n584), 
	.B1(n6807), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6338));
   INVX1 U1019 (.Y(n6807), 
	.A(\ram[0][2] ));
   OAI22X1 U1020 (.Y(n583), 
	.B1(n6808), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6306));
   INVX1 U1021 (.Y(n6808), 
	.A(\ram[0][1] ));
   OAI22X1 U1022 (.Y(n582), 
	.B1(n6809), 
	.B0(n6793), 
	.A1(n6792), 
	.A0(n6309));
   INVX1 U1023 (.Y(n6809), 
	.A(\ram[0][0] ));
   NOR2BX1 U1024 (.Y(n6793), 
	.B(n6792), 
	.AN(mem_write_en));
   NAND2X1 U1025 (.Y(n6792), 
	.B(n6514), 
	.A(n6534));
   OAI22X1 U1026 (.Y(n4677), 
	.B1(n6812), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6311));
   INVX1 U1027 (.Y(n6812), 
	.A(\ram[255][15] ));
   OAI22X1 U1028 (.Y(n4676), 
	.B1(n6813), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6314));
   INVX1 U1029 (.Y(n6813), 
	.A(\ram[255][14] ));
   OAI22X1 U1030 (.Y(n4675), 
	.B1(n6814), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6316));
   INVX1 U1031 (.Y(n6814), 
	.A(\ram[255][13] ));
   OAI22X1 U1032 (.Y(n4674), 
	.B1(n6815), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6318));
   INVX1 U1033 (.Y(n6815), 
	.A(\ram[255][12] ));
   OAI22X1 U1034 (.Y(n4673), 
	.B1(n6816), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6320));
   INVX1 U1035 (.Y(n6816), 
	.A(\ram[255][11] ));
   OAI22X1 U1036 (.Y(n4672), 
	.B1(n6817), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6322));
   INVX1 U1037 (.Y(n6817), 
	.A(\ram[255][10] ));
   OAI22X1 U1038 (.Y(n4671), 
	.B1(n6818), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6324));
   INVX1 U1039 (.Y(n6818), 
	.A(\ram[255][9] ));
   OAI22X1 U1040 (.Y(n4670), 
	.B1(n6819), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6326));
   INVX1 U1041 (.Y(n6819), 
	.A(\ram[255][8] ));
   OAI22X1 U1042 (.Y(n4669), 
	.B1(n6820), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6328));
   INVX1 U1043 (.Y(n6820), 
	.A(\ram[255][7] ));
   OAI22X1 U1044 (.Y(n4668), 
	.B1(n6821), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6330));
   INVX1 U1045 (.Y(n6821), 
	.A(\ram[255][6] ));
   OAI22X1 U1046 (.Y(n4667), 
	.B1(n6822), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6332));
   INVX1 U1047 (.Y(n6822), 
	.A(\ram[255][5] ));
   OAI22X1 U1048 (.Y(n4666), 
	.B1(n6823), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6334));
   INVX1 U1049 (.Y(n6823), 
	.A(\ram[255][4] ));
   OAI22X1 U1050 (.Y(n4665), 
	.B1(n6824), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6336));
   INVX1 U1051 (.Y(n6824), 
	.A(\ram[255][3] ));
   OAI22X1 U1052 (.Y(n4664), 
	.B1(n6825), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6338));
   INVX1 U1053 (.Y(n6825), 
	.A(\ram[255][2] ));
   OAI22X1 U1054 (.Y(n4663), 
	.B1(n6826), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6306));
   INVX1 U1055 (.Y(n6826), 
	.A(\ram[255][1] ));
   OAI22X1 U1056 (.Y(n4662), 
	.B1(n6827), 
	.B0(n6811), 
	.A1(n6810), 
	.A0(n6309));
   INVX1 U1057 (.Y(n6827), 
	.A(\ram[255][0] ));
   NOR2BX1 U1058 (.Y(n6811), 
	.B(n6810), 
	.AN(mem_write_en));
   NAND2X1 U1059 (.Y(n6810), 
	.B(n6533), 
	.A(n6828));
   OAI22X1 U1060 (.Y(n4661), 
	.B1(n6831), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6311));
   INVX1 U1061 (.Y(n6831), 
	.A(\ram[254][15] ));
   OAI22X1 U1062 (.Y(n4660), 
	.B1(n6832), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6314));
   INVX1 U1063 (.Y(n6832), 
	.A(\ram[254][14] ));
   OAI22X1 U1064 (.Y(n4659), 
	.B1(n6833), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6316));
   INVX1 U1065 (.Y(n6833), 
	.A(\ram[254][13] ));
   OAI22X1 U1066 (.Y(n4658), 
	.B1(n6834), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6318));
   INVX1 U1067 (.Y(n6834), 
	.A(\ram[254][12] ));
   OAI22X1 U1068 (.Y(n4657), 
	.B1(n6835), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6320));
   INVX1 U1069 (.Y(n6835), 
	.A(\ram[254][11] ));
   OAI22X1 U1070 (.Y(n4656), 
	.B1(n6836), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6322));
   INVX1 U1071 (.Y(n6836), 
	.A(\ram[254][10] ));
   OAI22X1 U1072 (.Y(n4655), 
	.B1(n6837), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6324));
   INVX1 U1073 (.Y(n6837), 
	.A(\ram[254][9] ));
   OAI22X1 U1074 (.Y(n4654), 
	.B1(n6838), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6326));
   INVX1 U1075 (.Y(n6838), 
	.A(\ram[254][8] ));
   OAI22X1 U1076 (.Y(n4653), 
	.B1(n6839), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6328));
   INVX1 U1077 (.Y(n6839), 
	.A(\ram[254][7] ));
   OAI22X1 U1078 (.Y(n4652), 
	.B1(n6840), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6330));
   INVX1 U1079 (.Y(n6840), 
	.A(\ram[254][6] ));
   OAI22X1 U1080 (.Y(n4651), 
	.B1(n6841), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6332));
   INVX1 U1081 (.Y(n6841), 
	.A(\ram[254][5] ));
   OAI22X1 U1082 (.Y(n4650), 
	.B1(n6842), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6334));
   INVX1 U1083 (.Y(n6842), 
	.A(\ram[254][4] ));
   OAI22X1 U1084 (.Y(n4649), 
	.B1(n6843), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6336));
   INVX1 U1085 (.Y(n6843), 
	.A(\ram[254][3] ));
   OAI22X1 U1086 (.Y(n4648), 
	.B1(n6844), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6338));
   INVX1 U1087 (.Y(n6844), 
	.A(\ram[254][2] ));
   OAI22X1 U1088 (.Y(n4647), 
	.B1(n6845), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6306));
   INVX1 U1089 (.Y(n6845), 
	.A(\ram[254][1] ));
   OAI22X1 U1090 (.Y(n4646), 
	.B1(n6846), 
	.B0(n6830), 
	.A1(n6829), 
	.A0(n6309));
   INVX1 U1091 (.Y(n6846), 
	.A(\ram[254][0] ));
   NOR2BX1 U1092 (.Y(n6830), 
	.B(n6829), 
	.AN(mem_write_en));
   NAND2X1 U1093 (.Y(n6829), 
	.B(n6553), 
	.A(n6828));
   OAI22X1 U1094 (.Y(n4645), 
	.B1(n6849), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6311));
   INVX1 U1095 (.Y(n6849), 
	.A(\ram[253][15] ));
   OAI22X1 U1096 (.Y(n4644), 
	.B1(n6850), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6314));
   INVX1 U1097 (.Y(n6850), 
	.A(\ram[253][14] ));
   OAI22X1 U1098 (.Y(n4643), 
	.B1(n6851), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6316));
   INVX1 U1099 (.Y(n6851), 
	.A(\ram[253][13] ));
   OAI22X1 U1100 (.Y(n4642), 
	.B1(n6852), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6318));
   INVX1 U1101 (.Y(n6852), 
	.A(\ram[253][12] ));
   OAI22X1 U1102 (.Y(n4641), 
	.B1(n6853), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6320));
   INVX1 U1103 (.Y(n6853), 
	.A(\ram[253][11] ));
   OAI22X1 U1104 (.Y(n4640), 
	.B1(n6854), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6322));
   INVX1 U1105 (.Y(n6854), 
	.A(\ram[253][10] ));
   OAI22X1 U1106 (.Y(n4639), 
	.B1(n6855), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6324));
   INVX1 U1107 (.Y(n6855), 
	.A(\ram[253][9] ));
   OAI22X1 U1108 (.Y(n4638), 
	.B1(n6856), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6326));
   INVX1 U1109 (.Y(n6856), 
	.A(\ram[253][8] ));
   OAI22X1 U1110 (.Y(n4637), 
	.B1(n6857), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6328));
   INVX1 U1111 (.Y(n6857), 
	.A(\ram[253][7] ));
   OAI22X1 U1112 (.Y(n4636), 
	.B1(n6858), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6330));
   INVX1 U1113 (.Y(n6858), 
	.A(\ram[253][6] ));
   OAI22X1 U1114 (.Y(n4635), 
	.B1(n6859), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6332));
   INVX1 U1115 (.Y(n6859), 
	.A(\ram[253][5] ));
   OAI22X1 U1116 (.Y(n4634), 
	.B1(n6860), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6334));
   INVX1 U1117 (.Y(n6860), 
	.A(\ram[253][4] ));
   OAI22X1 U1118 (.Y(n4633), 
	.B1(n6861), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6336));
   INVX1 U1119 (.Y(n6861), 
	.A(\ram[253][3] ));
   OAI22X1 U1120 (.Y(n4632), 
	.B1(n6862), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6338));
   INVX1 U1121 (.Y(n6862), 
	.A(\ram[253][2] ));
   OAI22X1 U1122 (.Y(n4631), 
	.B1(n6863), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6306));
   INVX1 U1123 (.Y(n6863), 
	.A(\ram[253][1] ));
   OAI22X1 U1124 (.Y(n4630), 
	.B1(n6864), 
	.B0(n6848), 
	.A1(n6847), 
	.A0(n6309));
   INVX1 U1125 (.Y(n6864), 
	.A(\ram[253][0] ));
   NOR2BX1 U1126 (.Y(n6848), 
	.B(n6847), 
	.AN(mem_write_en));
   NAND2X1 U1127 (.Y(n6847), 
	.B(n6572), 
	.A(n6828));
   OAI22X1 U1128 (.Y(n4629), 
	.B1(n6867), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6311));
   INVX1 U1129 (.Y(n6867), 
	.A(\ram[252][15] ));
   OAI22X1 U1130 (.Y(n4628), 
	.B1(n6868), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6314));
   INVX1 U1131 (.Y(n6868), 
	.A(\ram[252][14] ));
   OAI22X1 U1132 (.Y(n4627), 
	.B1(n6869), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6316));
   INVX1 U1133 (.Y(n6869), 
	.A(\ram[252][13] ));
   OAI22X1 U1134 (.Y(n4626), 
	.B1(n6870), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6318));
   INVX1 U1135 (.Y(n6870), 
	.A(\ram[252][12] ));
   OAI22X1 U1136 (.Y(n4625), 
	.B1(n6871), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6320));
   INVX1 U1137 (.Y(n6871), 
	.A(\ram[252][11] ));
   OAI22X1 U1138 (.Y(n4624), 
	.B1(n6872), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6322));
   INVX1 U1139 (.Y(n6872), 
	.A(\ram[252][10] ));
   OAI22X1 U1140 (.Y(n4623), 
	.B1(n6873), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6324));
   INVX1 U1141 (.Y(n6873), 
	.A(\ram[252][9] ));
   OAI22X1 U1142 (.Y(n4622), 
	.B1(n6874), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6326));
   INVX1 U1143 (.Y(n6874), 
	.A(\ram[252][8] ));
   OAI22X1 U1144 (.Y(n4621), 
	.B1(n6875), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6328));
   INVX1 U1145 (.Y(n6875), 
	.A(\ram[252][7] ));
   OAI22X1 U1146 (.Y(n4620), 
	.B1(n6876), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6330));
   INVX1 U1147 (.Y(n6876), 
	.A(\ram[252][6] ));
   OAI22X1 U1148 (.Y(n4619), 
	.B1(n6877), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6332));
   INVX1 U1149 (.Y(n6877), 
	.A(\ram[252][5] ));
   OAI22X1 U1150 (.Y(n4618), 
	.B1(n6878), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6334));
   INVX1 U1151 (.Y(n6878), 
	.A(\ram[252][4] ));
   OAI22X1 U1152 (.Y(n4617), 
	.B1(n6879), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6336));
   INVX1 U1153 (.Y(n6879), 
	.A(\ram[252][3] ));
   OAI22X1 U1154 (.Y(n4616), 
	.B1(n6880), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6338));
   INVX1 U1155 (.Y(n6880), 
	.A(\ram[252][2] ));
   OAI22X1 U1156 (.Y(n4615), 
	.B1(n6881), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6306));
   INVX1 U1157 (.Y(n6881), 
	.A(\ram[252][1] ));
   OAI22X1 U1158 (.Y(n4614), 
	.B1(n6882), 
	.B0(n6866), 
	.A1(n6865), 
	.A0(n6309));
   INVX1 U1159 (.Y(n6882), 
	.A(\ram[252][0] ));
   NOR2BX1 U1160 (.Y(n6866), 
	.B(n6865), 
	.AN(mem_write_en));
   NAND2X1 U1161 (.Y(n6865), 
	.B(n6591), 
	.A(n6828));
   OAI22X1 U1162 (.Y(n4613), 
	.B1(n6885), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6311));
   INVX1 U1163 (.Y(n6885), 
	.A(\ram[251][15] ));
   OAI22X1 U1164 (.Y(n4612), 
	.B1(n6886), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6314));
   INVX1 U1165 (.Y(n6886), 
	.A(\ram[251][14] ));
   OAI22X1 U1166 (.Y(n4611), 
	.B1(n6887), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6316));
   INVX1 U1167 (.Y(n6887), 
	.A(\ram[251][13] ));
   OAI22X1 U1168 (.Y(n4610), 
	.B1(n6888), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6318));
   INVX1 U1169 (.Y(n6888), 
	.A(\ram[251][12] ));
   OAI22X1 U1170 (.Y(n4609), 
	.B1(n6889), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6320));
   INVX1 U1171 (.Y(n6889), 
	.A(\ram[251][11] ));
   OAI22X1 U1172 (.Y(n4608), 
	.B1(n6890), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6322));
   INVX1 U1173 (.Y(n6890), 
	.A(\ram[251][10] ));
   OAI22X1 U1174 (.Y(n4607), 
	.B1(n6891), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6324));
   INVX1 U1175 (.Y(n6891), 
	.A(\ram[251][9] ));
   OAI22X1 U1176 (.Y(n4606), 
	.B1(n6892), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6326));
   INVX1 U1177 (.Y(n6892), 
	.A(\ram[251][8] ));
   OAI22X1 U1178 (.Y(n4605), 
	.B1(n6893), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6328));
   INVX1 U1179 (.Y(n6893), 
	.A(\ram[251][7] ));
   OAI22X1 U1180 (.Y(n4604), 
	.B1(n6894), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6330));
   INVX1 U1181 (.Y(n6894), 
	.A(\ram[251][6] ));
   OAI22X1 U1182 (.Y(n4603), 
	.B1(n6895), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6332));
   INVX1 U1183 (.Y(n6895), 
	.A(\ram[251][5] ));
   OAI22X1 U1184 (.Y(n4602), 
	.B1(n6896), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6334));
   INVX1 U1185 (.Y(n6896), 
	.A(\ram[251][4] ));
   OAI22X1 U1186 (.Y(n4601), 
	.B1(n6897), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6336));
   INVX1 U1187 (.Y(n6897), 
	.A(\ram[251][3] ));
   OAI22X1 U1188 (.Y(n4600), 
	.B1(n6898), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6338));
   INVX1 U1189 (.Y(n6898), 
	.A(\ram[251][2] ));
   OAI22X1 U1190 (.Y(n4599), 
	.B1(n6899), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6306));
   INVX1 U1191 (.Y(n6899), 
	.A(\ram[251][1] ));
   OAI22X1 U1192 (.Y(n4598), 
	.B1(n6900), 
	.B0(n6884), 
	.A1(n6883), 
	.A0(n6309));
   INVX1 U1193 (.Y(n6900), 
	.A(\ram[251][0] ));
   NOR2BX1 U1194 (.Y(n6884), 
	.B(n6883), 
	.AN(mem_write_en));
   NAND2X1 U1195 (.Y(n6883), 
	.B(n6610), 
	.A(n6828));
   OAI22X1 U1196 (.Y(n4597), 
	.B1(n6903), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6311));
   INVX1 U1197 (.Y(n6903), 
	.A(\ram[250][15] ));
   OAI22X1 U1198 (.Y(n4596), 
	.B1(n6904), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6314));
   INVX1 U1199 (.Y(n6904), 
	.A(\ram[250][14] ));
   OAI22X1 U1200 (.Y(n4595), 
	.B1(n6905), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6316));
   INVX1 U1201 (.Y(n6905), 
	.A(\ram[250][13] ));
   OAI22X1 U1202 (.Y(n4594), 
	.B1(n6906), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6318));
   INVX1 U1203 (.Y(n6906), 
	.A(\ram[250][12] ));
   OAI22X1 U1204 (.Y(n4593), 
	.B1(n6907), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6320));
   INVX1 U1205 (.Y(n6907), 
	.A(\ram[250][11] ));
   OAI22X1 U1206 (.Y(n4592), 
	.B1(n6908), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6322));
   INVX1 U1207 (.Y(n6908), 
	.A(\ram[250][10] ));
   OAI22X1 U1208 (.Y(n4591), 
	.B1(n6909), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6324));
   INVX1 U1209 (.Y(n6909), 
	.A(\ram[250][9] ));
   OAI22X1 U1210 (.Y(n4590), 
	.B1(n6910), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6326));
   INVX1 U1211 (.Y(n6910), 
	.A(\ram[250][8] ));
   OAI22X1 U1212 (.Y(n4589), 
	.B1(n6911), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6328));
   INVX1 U1213 (.Y(n6911), 
	.A(\ram[250][7] ));
   OAI22X1 U1214 (.Y(n4588), 
	.B1(n6912), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6330));
   INVX1 U1215 (.Y(n6912), 
	.A(\ram[250][6] ));
   OAI22X1 U1216 (.Y(n4587), 
	.B1(n6913), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6332));
   INVX1 U1217 (.Y(n6913), 
	.A(\ram[250][5] ));
   OAI22X1 U1218 (.Y(n4586), 
	.B1(n6914), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6334));
   INVX1 U1219 (.Y(n6914), 
	.A(\ram[250][4] ));
   OAI22X1 U1220 (.Y(n4585), 
	.B1(n6915), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6336));
   INVX1 U1221 (.Y(n6915), 
	.A(\ram[250][3] ));
   OAI22X1 U1222 (.Y(n4584), 
	.B1(n6916), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6338));
   INVX1 U1223 (.Y(n6916), 
	.A(\ram[250][2] ));
   OAI22X1 U1224 (.Y(n4583), 
	.B1(n6917), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6306));
   INVX1 U1225 (.Y(n6917), 
	.A(\ram[250][1] ));
   OAI22X1 U1226 (.Y(n4582), 
	.B1(n6918), 
	.B0(n6902), 
	.A1(n6901), 
	.A0(n6309));
   INVX1 U1227 (.Y(n6918), 
	.A(\ram[250][0] ));
   NOR2BX1 U1228 (.Y(n6902), 
	.B(n6901), 
	.AN(mem_write_en));
   NAND2X1 U1229 (.Y(n6901), 
	.B(n6629), 
	.A(n6828));
   OAI22X1 U1230 (.Y(n4581), 
	.B1(n6921), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6311));
   INVX1 U1231 (.Y(n6921), 
	.A(\ram[249][15] ));
   OAI22X1 U1232 (.Y(n4580), 
	.B1(n6922), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6314));
   INVX1 U1233 (.Y(n6922), 
	.A(\ram[249][14] ));
   OAI22X1 U1234 (.Y(n4579), 
	.B1(n6923), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6316));
   INVX1 U1235 (.Y(n6923), 
	.A(\ram[249][13] ));
   OAI22X1 U1236 (.Y(n4578), 
	.B1(n6924), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6318));
   INVX1 U1237 (.Y(n6924), 
	.A(\ram[249][12] ));
   OAI22X1 U1238 (.Y(n4577), 
	.B1(n6925), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6320));
   INVX1 U1239 (.Y(n6925), 
	.A(\ram[249][11] ));
   OAI22X1 U1240 (.Y(n4576), 
	.B1(n6926), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6322));
   INVX1 U1241 (.Y(n6926), 
	.A(\ram[249][10] ));
   OAI22X1 U1242 (.Y(n4575), 
	.B1(n6927), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6324));
   INVX1 U1243 (.Y(n6927), 
	.A(\ram[249][9] ));
   OAI22X1 U1244 (.Y(n4574), 
	.B1(n6928), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6326));
   INVX1 U1245 (.Y(n6928), 
	.A(\ram[249][8] ));
   OAI22X1 U1246 (.Y(n4573), 
	.B1(n6929), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6328));
   INVX1 U1247 (.Y(n6929), 
	.A(\ram[249][7] ));
   OAI22X1 U1248 (.Y(n4572), 
	.B1(n6930), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6330));
   INVX1 U1249 (.Y(n6930), 
	.A(\ram[249][6] ));
   OAI22X1 U1250 (.Y(n4571), 
	.B1(n6931), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6332));
   INVX1 U1251 (.Y(n6931), 
	.A(\ram[249][5] ));
   OAI22X1 U1252 (.Y(n4570), 
	.B1(n6932), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6334));
   INVX1 U1253 (.Y(n6932), 
	.A(\ram[249][4] ));
   OAI22X1 U1254 (.Y(n4569), 
	.B1(n6933), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6336));
   INVX1 U1255 (.Y(n6933), 
	.A(\ram[249][3] ));
   OAI22X1 U1256 (.Y(n4568), 
	.B1(n6934), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6338));
   INVX1 U1257 (.Y(n6934), 
	.A(\ram[249][2] ));
   OAI22X1 U1258 (.Y(n4567), 
	.B1(n6935), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6306));
   INVX1 U1259 (.Y(n6935), 
	.A(\ram[249][1] ));
   OAI22X1 U1260 (.Y(n4566), 
	.B1(n6936), 
	.B0(n6920), 
	.A1(n6919), 
	.A0(n6309));
   INVX1 U1261 (.Y(n6936), 
	.A(\ram[249][0] ));
   NOR2BX1 U1262 (.Y(n6920), 
	.B(n6919), 
	.AN(mem_write_en));
   NAND2X1 U1263 (.Y(n6919), 
	.B(n6342), 
	.A(n6828));
   OAI22X1 U1264 (.Y(n4565), 
	.B1(n6939), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6311));
   INVX1 U1265 (.Y(n6939), 
	.A(\ram[248][15] ));
   OAI22X1 U1266 (.Y(n4564), 
	.B1(n6940), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6314));
   INVX1 U1267 (.Y(n6940), 
	.A(\ram[248][14] ));
   OAI22X1 U1268 (.Y(n4563), 
	.B1(n6941), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6316));
   INVX1 U1269 (.Y(n6941), 
	.A(\ram[248][13] ));
   OAI22X1 U1270 (.Y(n4562), 
	.B1(n6942), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6318));
   INVX1 U1271 (.Y(n6942), 
	.A(\ram[248][12] ));
   OAI22X1 U1272 (.Y(n4561), 
	.B1(n6943), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6320));
   INVX1 U1273 (.Y(n6943), 
	.A(\ram[248][11] ));
   OAI22X1 U1274 (.Y(n4560), 
	.B1(n6944), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6322));
   INVX1 U1275 (.Y(n6944), 
	.A(\ram[248][10] ));
   OAI22X1 U1276 (.Y(n4559), 
	.B1(n6945), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6324));
   INVX1 U1277 (.Y(n6945), 
	.A(\ram[248][9] ));
   OAI22X1 U1278 (.Y(n4558), 
	.B1(n6946), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6326));
   INVX1 U1279 (.Y(n6946), 
	.A(\ram[248][8] ));
   OAI22X1 U1280 (.Y(n4557), 
	.B1(n6947), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6328));
   INVX1 U1281 (.Y(n6947), 
	.A(\ram[248][7] ));
   OAI22X1 U1282 (.Y(n4556), 
	.B1(n6948), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6330));
   INVX1 U1283 (.Y(n6948), 
	.A(\ram[248][6] ));
   OAI22X1 U1284 (.Y(n4555), 
	.B1(n6949), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6332));
   INVX1 U1285 (.Y(n6949), 
	.A(\ram[248][5] ));
   OAI22X1 U1286 (.Y(n4554), 
	.B1(n6950), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6334));
   INVX1 U1287 (.Y(n6950), 
	.A(\ram[248][4] ));
   OAI22X1 U1288 (.Y(n4553), 
	.B1(n6951), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6336));
   INVX1 U1289 (.Y(n6951), 
	.A(\ram[248][3] ));
   OAI22X1 U1290 (.Y(n4552), 
	.B1(n6952), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6338));
   INVX1 U1291 (.Y(n6952), 
	.A(\ram[248][2] ));
   OAI22X1 U1292 (.Y(n4551), 
	.B1(n6953), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6306));
   INVX1 U1293 (.Y(n6953), 
	.A(\ram[248][1] ));
   OAI22X1 U1294 (.Y(n4550), 
	.B1(n6954), 
	.B0(n6938), 
	.A1(n6937), 
	.A0(n6309));
   INVX1 U1295 (.Y(n6954), 
	.A(\ram[248][0] ));
   NOR2BX1 U1296 (.Y(n6938), 
	.B(n6937), 
	.AN(mem_write_en));
   NAND2X1 U1297 (.Y(n6937), 
	.B(n6362), 
	.A(n6828));
   OAI22X1 U1298 (.Y(n4549), 
	.B1(n6957), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6311));
   INVX1 U1299 (.Y(n6957), 
	.A(\ram[247][15] ));
   OAI22X1 U1300 (.Y(n4548), 
	.B1(n6958), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6314));
   INVX1 U1301 (.Y(n6958), 
	.A(\ram[247][14] ));
   OAI22X1 U1302 (.Y(n4547), 
	.B1(n6959), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6316));
   INVX1 U1303 (.Y(n6959), 
	.A(\ram[247][13] ));
   OAI22X1 U1304 (.Y(n4546), 
	.B1(n6960), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6318));
   INVX1 U1305 (.Y(n6960), 
	.A(\ram[247][12] ));
   OAI22X1 U1306 (.Y(n4545), 
	.B1(n6961), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6320));
   INVX1 U1307 (.Y(n6961), 
	.A(\ram[247][11] ));
   OAI22X1 U1308 (.Y(n4544), 
	.B1(n6962), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6322));
   INVX1 U1309 (.Y(n6962), 
	.A(\ram[247][10] ));
   OAI22X1 U1310 (.Y(n4543), 
	.B1(n6963), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6324));
   INVX1 U1311 (.Y(n6963), 
	.A(\ram[247][9] ));
   OAI22X1 U1312 (.Y(n4542), 
	.B1(n6964), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6326));
   INVX1 U1313 (.Y(n6964), 
	.A(\ram[247][8] ));
   OAI22X1 U1314 (.Y(n4541), 
	.B1(n6965), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6328));
   INVX1 U1315 (.Y(n6965), 
	.A(\ram[247][7] ));
   OAI22X1 U1316 (.Y(n4540), 
	.B1(n6966), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6330));
   INVX1 U1317 (.Y(n6966), 
	.A(\ram[247][6] ));
   OAI22X1 U1318 (.Y(n4539), 
	.B1(n6967), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6332));
   INVX1 U1319 (.Y(n6967), 
	.A(\ram[247][5] ));
   OAI22X1 U1320 (.Y(n4538), 
	.B1(n6968), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6334));
   INVX1 U1321 (.Y(n6968), 
	.A(\ram[247][4] ));
   OAI22X1 U1322 (.Y(n4537), 
	.B1(n6969), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6336));
   INVX1 U1323 (.Y(n6969), 
	.A(\ram[247][3] ));
   OAI22X1 U1324 (.Y(n4536), 
	.B1(n6970), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6338));
   INVX1 U1325 (.Y(n6970), 
	.A(\ram[247][2] ));
   OAI22X1 U1326 (.Y(n4535), 
	.B1(n6971), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6306));
   INVX1 U1327 (.Y(n6971), 
	.A(\ram[247][1] ));
   OAI22X1 U1328 (.Y(n4534), 
	.B1(n6972), 
	.B0(n6956), 
	.A1(n6955), 
	.A0(n6309));
   INVX1 U1329 (.Y(n6972), 
	.A(\ram[247][0] ));
   NOR2BX1 U1330 (.Y(n6956), 
	.B(n6955), 
	.AN(mem_write_en));
   NAND2X1 U1331 (.Y(n6955), 
	.B(n6381), 
	.A(n6828));
   OAI22X1 U1332 (.Y(n4533), 
	.B1(n6975), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6311));
   INVX1 U1333 (.Y(n6975), 
	.A(\ram[246][15] ));
   OAI22X1 U1334 (.Y(n4532), 
	.B1(n6976), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6314));
   INVX1 U1335 (.Y(n6976), 
	.A(\ram[246][14] ));
   OAI22X1 U1336 (.Y(n4531), 
	.B1(n6977), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6316));
   INVX1 U1337 (.Y(n6977), 
	.A(\ram[246][13] ));
   OAI22X1 U1338 (.Y(n4530), 
	.B1(n6978), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6318));
   INVX1 U1339 (.Y(n6978), 
	.A(\ram[246][12] ));
   OAI22X1 U1340 (.Y(n4529), 
	.B1(n6979), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6320));
   INVX1 U1341 (.Y(n6979), 
	.A(\ram[246][11] ));
   OAI22X1 U1342 (.Y(n4528), 
	.B1(n6980), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6322));
   INVX1 U1343 (.Y(n6980), 
	.A(\ram[246][10] ));
   OAI22X1 U1344 (.Y(n4527), 
	.B1(n6981), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6324));
   INVX1 U1345 (.Y(n6981), 
	.A(\ram[246][9] ));
   OAI22X1 U1346 (.Y(n4526), 
	.B1(n6982), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6326));
   INVX1 U1347 (.Y(n6982), 
	.A(\ram[246][8] ));
   OAI22X1 U1348 (.Y(n4525), 
	.B1(n6983), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6328));
   INVX1 U1349 (.Y(n6983), 
	.A(\ram[246][7] ));
   OAI22X1 U1350 (.Y(n4524), 
	.B1(n6984), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6330));
   INVX1 U1351 (.Y(n6984), 
	.A(\ram[246][6] ));
   OAI22X1 U1352 (.Y(n4523), 
	.B1(n6985), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6332));
   INVX1 U1353 (.Y(n6985), 
	.A(\ram[246][5] ));
   OAI22X1 U1354 (.Y(n4522), 
	.B1(n6986), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6334));
   INVX1 U1355 (.Y(n6986), 
	.A(\ram[246][4] ));
   OAI22X1 U1356 (.Y(n4521), 
	.B1(n6987), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6336));
   INVX1 U1357 (.Y(n6987), 
	.A(\ram[246][3] ));
   OAI22X1 U1358 (.Y(n4520), 
	.B1(n6988), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6338));
   INVX1 U1359 (.Y(n6988), 
	.A(\ram[246][2] ));
   OAI22X1 U1360 (.Y(n4519), 
	.B1(n6989), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6306));
   INVX1 U1361 (.Y(n6989), 
	.A(\ram[246][1] ));
   OAI22X1 U1362 (.Y(n4518), 
	.B1(n6990), 
	.B0(n6974), 
	.A1(n6973), 
	.A0(n6309));
   INVX1 U1363 (.Y(n6990), 
	.A(\ram[246][0] ));
   NOR2BX1 U1364 (.Y(n6974), 
	.B(n6973), 
	.AN(mem_write_en));
   NAND2X1 U1365 (.Y(n6973), 
	.B(n6400), 
	.A(n6828));
   OAI22X1 U1366 (.Y(n4517), 
	.B1(n6993), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6311));
   INVX1 U1367 (.Y(n6993), 
	.A(\ram[245][15] ));
   OAI22X1 U1368 (.Y(n4516), 
	.B1(n6994), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6314));
   INVX1 U1369 (.Y(n6994), 
	.A(\ram[245][14] ));
   OAI22X1 U1370 (.Y(n4515), 
	.B1(n6995), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6316));
   INVX1 U1371 (.Y(n6995), 
	.A(\ram[245][13] ));
   OAI22X1 U1372 (.Y(n4514), 
	.B1(n6996), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6318));
   INVX1 U1373 (.Y(n6996), 
	.A(\ram[245][12] ));
   OAI22X1 U1374 (.Y(n4513), 
	.B1(n6997), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6320));
   INVX1 U1375 (.Y(n6997), 
	.A(\ram[245][11] ));
   OAI22X1 U1376 (.Y(n4512), 
	.B1(n6998), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6322));
   INVX1 U1377 (.Y(n6998), 
	.A(\ram[245][10] ));
   OAI22X1 U1378 (.Y(n4511), 
	.B1(n6999), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6324));
   INVX1 U1379 (.Y(n6999), 
	.A(\ram[245][9] ));
   OAI22X1 U1380 (.Y(n4510), 
	.B1(n7000), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6326));
   INVX1 U1381 (.Y(n7000), 
	.A(\ram[245][8] ));
   OAI22X1 U1382 (.Y(n4509), 
	.B1(n7001), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6328));
   INVX1 U1383 (.Y(n7001), 
	.A(\ram[245][7] ));
   OAI22X1 U1384 (.Y(n4508), 
	.B1(n7002), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6330));
   INVX1 U1385 (.Y(n7002), 
	.A(\ram[245][6] ));
   OAI22X1 U1386 (.Y(n4507), 
	.B1(n7003), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6332));
   INVX1 U1387 (.Y(n7003), 
	.A(\ram[245][5] ));
   OAI22X1 U1388 (.Y(n4506), 
	.B1(n7004), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6334));
   INVX1 U1389 (.Y(n7004), 
	.A(\ram[245][4] ));
   OAI22X1 U1390 (.Y(n4505), 
	.B1(n7005), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6336));
   INVX1 U1391 (.Y(n7005), 
	.A(\ram[245][3] ));
   OAI22X1 U1392 (.Y(n4504), 
	.B1(n7006), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6338));
   INVX1 U1393 (.Y(n7006), 
	.A(\ram[245][2] ));
   OAI22X1 U1394 (.Y(n4503), 
	.B1(n7007), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6306));
   INVX1 U1395 (.Y(n7007), 
	.A(\ram[245][1] ));
   OAI22X1 U1396 (.Y(n4502), 
	.B1(n7008), 
	.B0(n6992), 
	.A1(n6991), 
	.A0(n6309));
   INVX1 U1397 (.Y(n7008), 
	.A(\ram[245][0] ));
   NOR2BX1 U1398 (.Y(n6992), 
	.B(n6991), 
	.AN(mem_write_en));
   NAND2X1 U1399 (.Y(n6991), 
	.B(n6419), 
	.A(n6828));
   OAI22X1 U1400 (.Y(n4501), 
	.B1(n7011), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6311));
   INVX1 U1401 (.Y(n7011), 
	.A(\ram[244][15] ));
   OAI22X1 U1402 (.Y(n4500), 
	.B1(n7012), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6314));
   INVX1 U1403 (.Y(n7012), 
	.A(\ram[244][14] ));
   OAI22X1 U1404 (.Y(n4499), 
	.B1(n7013), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6316));
   INVX1 U1405 (.Y(n7013), 
	.A(\ram[244][13] ));
   OAI22X1 U1406 (.Y(n4498), 
	.B1(n7014), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6318));
   INVX1 U1407 (.Y(n7014), 
	.A(\ram[244][12] ));
   OAI22X1 U1408 (.Y(n4497), 
	.B1(n7015), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6320));
   INVX1 U1409 (.Y(n7015), 
	.A(\ram[244][11] ));
   OAI22X1 U1410 (.Y(n4496), 
	.B1(n7016), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6322));
   INVX1 U1411 (.Y(n7016), 
	.A(\ram[244][10] ));
   OAI22X1 U1412 (.Y(n4495), 
	.B1(n7017), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6324));
   INVX1 U1413 (.Y(n7017), 
	.A(\ram[244][9] ));
   OAI22X1 U1414 (.Y(n4494), 
	.B1(n7018), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6326));
   INVX1 U1415 (.Y(n7018), 
	.A(\ram[244][8] ));
   OAI22X1 U1416 (.Y(n4493), 
	.B1(n7019), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6328));
   INVX1 U1417 (.Y(n7019), 
	.A(\ram[244][7] ));
   OAI22X1 U1418 (.Y(n4492), 
	.B1(n7020), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6330));
   INVX1 U1419 (.Y(n7020), 
	.A(\ram[244][6] ));
   OAI22X1 U1420 (.Y(n4491), 
	.B1(n7021), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6332));
   INVX1 U1421 (.Y(n7021), 
	.A(\ram[244][5] ));
   OAI22X1 U1422 (.Y(n4490), 
	.B1(n7022), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6334));
   INVX1 U1423 (.Y(n7022), 
	.A(\ram[244][4] ));
   OAI22X1 U1424 (.Y(n4489), 
	.B1(n7023), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6336));
   INVX1 U1425 (.Y(n7023), 
	.A(\ram[244][3] ));
   OAI22X1 U1426 (.Y(n4488), 
	.B1(n7024), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6338));
   INVX1 U1427 (.Y(n7024), 
	.A(\ram[244][2] ));
   OAI22X1 U1428 (.Y(n4487), 
	.B1(n7025), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6306));
   INVX1 U1429 (.Y(n7025), 
	.A(\ram[244][1] ));
   OAI22X1 U1430 (.Y(n4486), 
	.B1(n7026), 
	.B0(n7010), 
	.A1(n7009), 
	.A0(n6309));
   INVX1 U1431 (.Y(n7026), 
	.A(\ram[244][0] ));
   NOR2BX1 U1432 (.Y(n7010), 
	.B(n7009), 
	.AN(mem_write_en));
   NAND2X1 U1433 (.Y(n7009), 
	.B(n6438), 
	.A(n6828));
   OAI22X1 U1434 (.Y(n4485), 
	.B1(n7029), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6311));
   INVX1 U1435 (.Y(n7029), 
	.A(\ram[243][15] ));
   OAI22X1 U1436 (.Y(n4484), 
	.B1(n7030), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6314));
   INVX1 U1437 (.Y(n7030), 
	.A(\ram[243][14] ));
   OAI22X1 U1438 (.Y(n4483), 
	.B1(n7031), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6316));
   INVX1 U1439 (.Y(n7031), 
	.A(\ram[243][13] ));
   OAI22X1 U1440 (.Y(n4482), 
	.B1(n7032), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6318));
   INVX1 U1441 (.Y(n7032), 
	.A(\ram[243][12] ));
   OAI22X1 U1442 (.Y(n4481), 
	.B1(n7033), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6320));
   INVX1 U1443 (.Y(n7033), 
	.A(\ram[243][11] ));
   OAI22X1 U1444 (.Y(n4480), 
	.B1(n7034), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6322));
   INVX1 U1445 (.Y(n7034), 
	.A(\ram[243][10] ));
   OAI22X1 U1446 (.Y(n4479), 
	.B1(n7035), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6324));
   INVX1 U1447 (.Y(n7035), 
	.A(\ram[243][9] ));
   OAI22X1 U1448 (.Y(n4478), 
	.B1(n7036), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6326));
   INVX1 U1449 (.Y(n7036), 
	.A(\ram[243][8] ));
   OAI22X1 U1450 (.Y(n4477), 
	.B1(n7037), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6328));
   INVX1 U1451 (.Y(n7037), 
	.A(\ram[243][7] ));
   OAI22X1 U1452 (.Y(n4476), 
	.B1(n7038), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6330));
   INVX1 U1453 (.Y(n7038), 
	.A(\ram[243][6] ));
   OAI22X1 U1454 (.Y(n4475), 
	.B1(n7039), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6332));
   INVX1 U1455 (.Y(n7039), 
	.A(\ram[243][5] ));
   OAI22X1 U1456 (.Y(n4474), 
	.B1(n7040), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6334));
   INVX1 U1457 (.Y(n7040), 
	.A(\ram[243][4] ));
   OAI22X1 U1458 (.Y(n4473), 
	.B1(n7041), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6336));
   INVX1 U1459 (.Y(n7041), 
	.A(\ram[243][3] ));
   OAI22X1 U1460 (.Y(n4472), 
	.B1(n7042), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6338));
   INVX1 U1461 (.Y(n7042), 
	.A(\ram[243][2] ));
   OAI22X1 U1462 (.Y(n4471), 
	.B1(n7043), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6306));
   INVX1 U1463 (.Y(n7043), 
	.A(\ram[243][1] ));
   OAI22X1 U1464 (.Y(n4470), 
	.B1(n7044), 
	.B0(n7028), 
	.A1(n7027), 
	.A0(n6309));
   INVX1 U1465 (.Y(n7044), 
	.A(\ram[243][0] ));
   NOR2BX1 U1466 (.Y(n7028), 
	.B(n7027), 
	.AN(mem_write_en));
   NAND2X1 U1467 (.Y(n7027), 
	.B(n6457), 
	.A(n6828));
   OAI22X1 U1468 (.Y(n4469), 
	.B1(n7047), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6311));
   INVX1 U1469 (.Y(n7047), 
	.A(\ram[242][15] ));
   OAI22X1 U1470 (.Y(n4468), 
	.B1(n7048), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6314));
   INVX1 U1471 (.Y(n7048), 
	.A(\ram[242][14] ));
   OAI22X1 U1472 (.Y(n4467), 
	.B1(n7049), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6316));
   INVX1 U1473 (.Y(n7049), 
	.A(\ram[242][13] ));
   OAI22X1 U1474 (.Y(n4466), 
	.B1(n7050), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6318));
   INVX1 U1475 (.Y(n7050), 
	.A(\ram[242][12] ));
   OAI22X1 U1476 (.Y(n4465), 
	.B1(n7051), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6320));
   INVX1 U1477 (.Y(n7051), 
	.A(\ram[242][11] ));
   OAI22X1 U1478 (.Y(n4464), 
	.B1(n7052), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6322));
   INVX1 U1479 (.Y(n7052), 
	.A(\ram[242][10] ));
   OAI22X1 U1480 (.Y(n4463), 
	.B1(n7053), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6324));
   INVX1 U1481 (.Y(n7053), 
	.A(\ram[242][9] ));
   OAI22X1 U1482 (.Y(n4462), 
	.B1(n7054), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6326));
   INVX1 U1483 (.Y(n7054), 
	.A(\ram[242][8] ));
   OAI22X1 U1484 (.Y(n4461), 
	.B1(n7055), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6328));
   INVX1 U1485 (.Y(n7055), 
	.A(\ram[242][7] ));
   OAI22X1 U1486 (.Y(n4460), 
	.B1(n7056), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6330));
   INVX1 U1487 (.Y(n7056), 
	.A(\ram[242][6] ));
   OAI22X1 U1488 (.Y(n4459), 
	.B1(n7057), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6332));
   INVX1 U1489 (.Y(n7057), 
	.A(\ram[242][5] ));
   OAI22X1 U1490 (.Y(n4458), 
	.B1(n7058), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6334));
   INVX1 U1491 (.Y(n7058), 
	.A(\ram[242][4] ));
   OAI22X1 U1492 (.Y(n4457), 
	.B1(n7059), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6336));
   INVX1 U1493 (.Y(n7059), 
	.A(\ram[242][3] ));
   OAI22X1 U1494 (.Y(n4456), 
	.B1(n7060), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6338));
   INVX1 U1495 (.Y(n7060), 
	.A(\ram[242][2] ));
   OAI22X1 U1496 (.Y(n4455), 
	.B1(n7061), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6306));
   INVX1 U1497 (.Y(n7061), 
	.A(\ram[242][1] ));
   OAI22X1 U1498 (.Y(n4454), 
	.B1(n7062), 
	.B0(n7046), 
	.A1(n7045), 
	.A0(n6309));
   INVX1 U1499 (.Y(n7062), 
	.A(\ram[242][0] ));
   NOR2BX1 U1500 (.Y(n7046), 
	.B(n7045), 
	.AN(mem_write_en));
   NAND2X1 U1501 (.Y(n7045), 
	.B(n6476), 
	.A(n6828));
   OAI22X1 U1502 (.Y(n4453), 
	.B1(n7065), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6311));
   INVX1 U1503 (.Y(n7065), 
	.A(\ram[241][15] ));
   OAI22X1 U1504 (.Y(n4452), 
	.B1(n7066), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6314));
   INVX1 U1505 (.Y(n7066), 
	.A(\ram[241][14] ));
   OAI22X1 U1506 (.Y(n4451), 
	.B1(n7067), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6316));
   INVX1 U1507 (.Y(n7067), 
	.A(\ram[241][13] ));
   OAI22X1 U1508 (.Y(n4450), 
	.B1(n7068), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6318));
   INVX1 U1509 (.Y(n7068), 
	.A(\ram[241][12] ));
   OAI22X1 U1510 (.Y(n4449), 
	.B1(n7069), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6320));
   INVX1 U1511 (.Y(n7069), 
	.A(\ram[241][11] ));
   OAI22X1 U1512 (.Y(n4448), 
	.B1(n7070), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6322));
   INVX1 U1513 (.Y(n7070), 
	.A(\ram[241][10] ));
   OAI22X1 U1514 (.Y(n4447), 
	.B1(n7071), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6324));
   INVX1 U1515 (.Y(n7071), 
	.A(\ram[241][9] ));
   OAI22X1 U1516 (.Y(n4446), 
	.B1(n7072), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6326));
   INVX1 U1517 (.Y(n7072), 
	.A(\ram[241][8] ));
   OAI22X1 U1518 (.Y(n4445), 
	.B1(n7073), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6328));
   INVX1 U1519 (.Y(n7073), 
	.A(\ram[241][7] ));
   OAI22X1 U1520 (.Y(n4444), 
	.B1(n7074), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6330));
   INVX1 U1521 (.Y(n7074), 
	.A(\ram[241][6] ));
   OAI22X1 U1522 (.Y(n4443), 
	.B1(n7075), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6332));
   INVX1 U1523 (.Y(n7075), 
	.A(\ram[241][5] ));
   OAI22X1 U1524 (.Y(n4442), 
	.B1(n7076), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6334));
   INVX1 U1525 (.Y(n7076), 
	.A(\ram[241][4] ));
   OAI22X1 U1526 (.Y(n4441), 
	.B1(n7077), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6336));
   INVX1 U1527 (.Y(n7077), 
	.A(\ram[241][3] ));
   OAI22X1 U1528 (.Y(n4440), 
	.B1(n7078), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6338));
   INVX1 U1529 (.Y(n7078), 
	.A(\ram[241][2] ));
   OAI22X1 U1530 (.Y(n4439), 
	.B1(n7079), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6306));
   INVX1 U1531 (.Y(n7079), 
	.A(\ram[241][1] ));
   OAI22X1 U1532 (.Y(n4438), 
	.B1(n7080), 
	.B0(n7064), 
	.A1(n7063), 
	.A0(n6309));
   INVX1 U1533 (.Y(n7080), 
	.A(\ram[241][0] ));
   NOR2BX1 U1534 (.Y(n7064), 
	.B(n7063), 
	.AN(mem_write_en));
   NAND2X1 U1535 (.Y(n7063), 
	.B(n6495), 
	.A(n6828));
   OAI22X1 U1536 (.Y(n4437), 
	.B1(n7083), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6311));
   INVX1 U1537 (.Y(n7083), 
	.A(\ram[240][15] ));
   OAI22X1 U1538 (.Y(n4436), 
	.B1(n7084), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6314));
   INVX1 U1539 (.Y(n7084), 
	.A(\ram[240][14] ));
   OAI22X1 U1540 (.Y(n4435), 
	.B1(n7085), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6316));
   INVX1 U1541 (.Y(n7085), 
	.A(\ram[240][13] ));
   OAI22X1 U1542 (.Y(n4434), 
	.B1(n7086), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6318));
   INVX1 U1543 (.Y(n7086), 
	.A(\ram[240][12] ));
   OAI22X1 U1544 (.Y(n4433), 
	.B1(n7087), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6320));
   INVX1 U1545 (.Y(n7087), 
	.A(\ram[240][11] ));
   OAI22X1 U1546 (.Y(n4432), 
	.B1(n7088), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6322));
   INVX1 U1547 (.Y(n7088), 
	.A(\ram[240][10] ));
   OAI22X1 U1548 (.Y(n4431), 
	.B1(n7089), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6324));
   INVX1 U1549 (.Y(n7089), 
	.A(\ram[240][9] ));
   OAI22X1 U1550 (.Y(n4430), 
	.B1(n7090), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6326));
   INVX1 U1551 (.Y(n7090), 
	.A(\ram[240][8] ));
   OAI22X1 U1552 (.Y(n4429), 
	.B1(n7091), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6328));
   INVX1 U1553 (.Y(n7091), 
	.A(\ram[240][7] ));
   OAI22X1 U1554 (.Y(n4428), 
	.B1(n7092), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6330));
   INVX1 U1555 (.Y(n7092), 
	.A(\ram[240][6] ));
   OAI22X1 U1556 (.Y(n4427), 
	.B1(n7093), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6332));
   INVX1 U1557 (.Y(n7093), 
	.A(\ram[240][5] ));
   OAI22X1 U1558 (.Y(n4426), 
	.B1(n7094), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6334));
   INVX1 U1559 (.Y(n7094), 
	.A(\ram[240][4] ));
   OAI22X1 U1560 (.Y(n4425), 
	.B1(n7095), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6336));
   INVX1 U1561 (.Y(n7095), 
	.A(\ram[240][3] ));
   OAI22X1 U1562 (.Y(n4424), 
	.B1(n7096), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6338));
   INVX1 U1563 (.Y(n7096), 
	.A(\ram[240][2] ));
   OAI22X1 U1564 (.Y(n4423), 
	.B1(n7097), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6306));
   INVX1 U1565 (.Y(n7097), 
	.A(\ram[240][1] ));
   OAI22X1 U1566 (.Y(n4422), 
	.B1(n7098), 
	.B0(n7082), 
	.A1(n7081), 
	.A0(n6309));
   INVX1 U1567 (.Y(n7098), 
	.A(\ram[240][0] ));
   NOR2BX1 U1568 (.Y(n7082), 
	.B(n7081), 
	.AN(mem_write_en));
   NAND2X1 U1569 (.Y(n7081), 
	.B(n6514), 
	.A(n6828));
   OAI22X1 U1570 (.Y(n4421), 
	.B1(n7101), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6311));
   INVX1 U1571 (.Y(n7101), 
	.A(\ram[239][15] ));
   OAI22X1 U1572 (.Y(n4420), 
	.B1(n7102), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6314));
   INVX1 U1573 (.Y(n7102), 
	.A(\ram[239][14] ));
   OAI22X1 U1574 (.Y(n4419), 
	.B1(n7103), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6316));
   INVX1 U1575 (.Y(n7103), 
	.A(\ram[239][13] ));
   OAI22X1 U1576 (.Y(n4418), 
	.B1(n7104), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6318));
   INVX1 U1577 (.Y(n7104), 
	.A(\ram[239][12] ));
   OAI22X1 U1578 (.Y(n4417), 
	.B1(n7105), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6320));
   INVX1 U1579 (.Y(n7105), 
	.A(\ram[239][11] ));
   OAI22X1 U1580 (.Y(n4416), 
	.B1(n7106), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6322));
   INVX1 U1581 (.Y(n7106), 
	.A(\ram[239][10] ));
   OAI22X1 U1582 (.Y(n4415), 
	.B1(n7107), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6324));
   INVX1 U1583 (.Y(n7107), 
	.A(\ram[239][9] ));
   OAI22X1 U1584 (.Y(n4414), 
	.B1(n7108), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6326));
   INVX1 U1585 (.Y(n7108), 
	.A(\ram[239][8] ));
   OAI22X1 U1586 (.Y(n4413), 
	.B1(n7109), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6328));
   INVX1 U1587 (.Y(n7109), 
	.A(\ram[239][7] ));
   OAI22X1 U1588 (.Y(n4412), 
	.B1(n7110), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6330));
   INVX1 U1589 (.Y(n7110), 
	.A(\ram[239][6] ));
   OAI22X1 U1590 (.Y(n4411), 
	.B1(n7111), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6332));
   INVX1 U1591 (.Y(n7111), 
	.A(\ram[239][5] ));
   OAI22X1 U1592 (.Y(n4410), 
	.B1(n7112), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6334));
   INVX1 U1593 (.Y(n7112), 
	.A(\ram[239][4] ));
   OAI22X1 U1594 (.Y(n4409), 
	.B1(n7113), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6336));
   INVX1 U1595 (.Y(n7113), 
	.A(\ram[239][3] ));
   OAI22X1 U1596 (.Y(n4408), 
	.B1(n7114), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6338));
   INVX1 U1597 (.Y(n7114), 
	.A(\ram[239][2] ));
   OAI22X1 U1598 (.Y(n4407), 
	.B1(n7115), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6306));
   INVX1 U1599 (.Y(n7115), 
	.A(\ram[239][1] ));
   OAI22X1 U1600 (.Y(n4406), 
	.B1(n7116), 
	.B0(n7100), 
	.A1(n7099), 
	.A0(n6309));
   INVX1 U1601 (.Y(n7116), 
	.A(\ram[239][0] ));
   NOR2BX1 U1602 (.Y(n7100), 
	.B(n7099), 
	.AN(mem_write_en));
   NAND2X1 U1603 (.Y(n7099), 
	.B(n6533), 
	.A(n7117));
   OAI22X1 U1604 (.Y(n4405), 
	.B1(n7120), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6311));
   INVX1 U1605 (.Y(n7120), 
	.A(\ram[238][15] ));
   OAI22X1 U1606 (.Y(n4404), 
	.B1(n7121), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6314));
   INVX1 U1607 (.Y(n7121), 
	.A(\ram[238][14] ));
   OAI22X1 U1608 (.Y(n4403), 
	.B1(n7122), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6316));
   INVX1 U1609 (.Y(n7122), 
	.A(\ram[238][13] ));
   OAI22X1 U1610 (.Y(n4402), 
	.B1(n7123), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6318));
   INVX1 U1611 (.Y(n7123), 
	.A(\ram[238][12] ));
   OAI22X1 U1612 (.Y(n4401), 
	.B1(n7124), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6320));
   INVX1 U1613 (.Y(n7124), 
	.A(\ram[238][11] ));
   OAI22X1 U1614 (.Y(n4400), 
	.B1(n7125), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6322));
   INVX1 U1615 (.Y(n7125), 
	.A(\ram[238][10] ));
   OAI22X1 U1616 (.Y(n4399), 
	.B1(n7126), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6324));
   INVX1 U1617 (.Y(n7126), 
	.A(\ram[238][9] ));
   OAI22X1 U1618 (.Y(n4398), 
	.B1(n7127), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6326));
   INVX1 U1619 (.Y(n7127), 
	.A(\ram[238][8] ));
   OAI22X1 U1620 (.Y(n4397), 
	.B1(n7128), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6328));
   INVX1 U1621 (.Y(n7128), 
	.A(\ram[238][7] ));
   OAI22X1 U1622 (.Y(n4396), 
	.B1(n7129), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6330));
   INVX1 U1623 (.Y(n7129), 
	.A(\ram[238][6] ));
   OAI22X1 U1624 (.Y(n4395), 
	.B1(n7130), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6332));
   INVX1 U1625 (.Y(n7130), 
	.A(\ram[238][5] ));
   OAI22X1 U1626 (.Y(n4394), 
	.B1(n7131), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6334));
   INVX1 U1627 (.Y(n7131), 
	.A(\ram[238][4] ));
   OAI22X1 U1628 (.Y(n4393), 
	.B1(n7132), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6336));
   INVX1 U1629 (.Y(n7132), 
	.A(\ram[238][3] ));
   OAI22X1 U1630 (.Y(n4392), 
	.B1(n7133), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6338));
   INVX1 U1631 (.Y(n7133), 
	.A(\ram[238][2] ));
   OAI22X1 U1632 (.Y(n4391), 
	.B1(n7134), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6306));
   INVX1 U1633 (.Y(n7134), 
	.A(\ram[238][1] ));
   OAI22X1 U1634 (.Y(n4390), 
	.B1(n7135), 
	.B0(n7119), 
	.A1(n7118), 
	.A0(n6309));
   INVX1 U1635 (.Y(n7135), 
	.A(\ram[238][0] ));
   NOR2BX1 U1636 (.Y(n7119), 
	.B(n7118), 
	.AN(mem_write_en));
   NAND2X1 U1637 (.Y(n7118), 
	.B(n6553), 
	.A(n7117));
   OAI22X1 U1638 (.Y(n4389), 
	.B1(n7138), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6311));
   INVX1 U1639 (.Y(n7138), 
	.A(\ram[237][15] ));
   OAI22X1 U1640 (.Y(n4388), 
	.B1(n7139), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6314));
   INVX1 U1641 (.Y(n7139), 
	.A(\ram[237][14] ));
   OAI22X1 U1642 (.Y(n4387), 
	.B1(n7140), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6316));
   INVX1 U1643 (.Y(n7140), 
	.A(\ram[237][13] ));
   OAI22X1 U1644 (.Y(n4386), 
	.B1(n7141), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6318));
   INVX1 U1645 (.Y(n7141), 
	.A(\ram[237][12] ));
   OAI22X1 U1646 (.Y(n4385), 
	.B1(n7142), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6320));
   INVX1 U1647 (.Y(n7142), 
	.A(\ram[237][11] ));
   OAI22X1 U1648 (.Y(n4384), 
	.B1(n7143), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6322));
   INVX1 U1649 (.Y(n7143), 
	.A(\ram[237][10] ));
   OAI22X1 U1650 (.Y(n4383), 
	.B1(n7144), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6324));
   INVX1 U1651 (.Y(n7144), 
	.A(\ram[237][9] ));
   OAI22X1 U1652 (.Y(n4382), 
	.B1(n7145), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6326));
   INVX1 U1653 (.Y(n7145), 
	.A(\ram[237][8] ));
   OAI22X1 U1654 (.Y(n4381), 
	.B1(n7146), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6328));
   INVX1 U1655 (.Y(n7146), 
	.A(\ram[237][7] ));
   OAI22X1 U1656 (.Y(n4380), 
	.B1(n7147), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6330));
   INVX1 U1657 (.Y(n7147), 
	.A(\ram[237][6] ));
   OAI22X1 U1658 (.Y(n4379), 
	.B1(n7148), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6332));
   INVX1 U1659 (.Y(n7148), 
	.A(\ram[237][5] ));
   OAI22X1 U1660 (.Y(n4378), 
	.B1(n7149), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6334));
   INVX1 U1661 (.Y(n7149), 
	.A(\ram[237][4] ));
   OAI22X1 U1662 (.Y(n4377), 
	.B1(n7150), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6336));
   INVX1 U1663 (.Y(n7150), 
	.A(\ram[237][3] ));
   OAI22X1 U1664 (.Y(n4376), 
	.B1(n7151), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6338));
   INVX1 U1665 (.Y(n7151), 
	.A(\ram[237][2] ));
   OAI22X1 U1666 (.Y(n4375), 
	.B1(n7152), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6306));
   INVX1 U1667 (.Y(n7152), 
	.A(\ram[237][1] ));
   OAI22X1 U1668 (.Y(n4374), 
	.B1(n7153), 
	.B0(n7137), 
	.A1(n7136), 
	.A0(n6309));
   INVX1 U1669 (.Y(n7153), 
	.A(\ram[237][0] ));
   NOR2BX1 U1670 (.Y(n7137), 
	.B(n7136), 
	.AN(mem_write_en));
   NAND2X1 U1671 (.Y(n7136), 
	.B(n6572), 
	.A(n7117));
   OAI22X1 U1672 (.Y(n4373), 
	.B1(n7156), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6311));
   INVX1 U1673 (.Y(n7156), 
	.A(\ram[236][15] ));
   OAI22X1 U1674 (.Y(n4372), 
	.B1(n7157), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6314));
   INVX1 U1675 (.Y(n7157), 
	.A(\ram[236][14] ));
   OAI22X1 U1676 (.Y(n4371), 
	.B1(n7158), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6316));
   INVX1 U1677 (.Y(n7158), 
	.A(\ram[236][13] ));
   OAI22X1 U1678 (.Y(n4370), 
	.B1(n7159), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6318));
   INVX1 U1679 (.Y(n7159), 
	.A(\ram[236][12] ));
   OAI22X1 U1680 (.Y(n4369), 
	.B1(n7160), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6320));
   INVX1 U1681 (.Y(n7160), 
	.A(\ram[236][11] ));
   OAI22X1 U1682 (.Y(n4368), 
	.B1(n7161), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6322));
   INVX1 U1683 (.Y(n7161), 
	.A(\ram[236][10] ));
   OAI22X1 U1684 (.Y(n4367), 
	.B1(n7162), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6324));
   INVX1 U1685 (.Y(n7162), 
	.A(\ram[236][9] ));
   OAI22X1 U1686 (.Y(n4366), 
	.B1(n7163), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6326));
   INVX1 U1687 (.Y(n7163), 
	.A(\ram[236][8] ));
   OAI22X1 U1688 (.Y(n4365), 
	.B1(n7164), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6328));
   INVX1 U1689 (.Y(n7164), 
	.A(\ram[236][7] ));
   OAI22X1 U1690 (.Y(n4364), 
	.B1(n7165), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6330));
   INVX1 U1691 (.Y(n7165), 
	.A(\ram[236][6] ));
   OAI22X1 U1692 (.Y(n4363), 
	.B1(n7166), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6332));
   INVX1 U1693 (.Y(n7166), 
	.A(\ram[236][5] ));
   OAI22X1 U1694 (.Y(n4362), 
	.B1(n7167), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6334));
   INVX1 U1695 (.Y(n7167), 
	.A(\ram[236][4] ));
   OAI22X1 U1696 (.Y(n4361), 
	.B1(n7168), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6336));
   INVX1 U1697 (.Y(n7168), 
	.A(\ram[236][3] ));
   OAI22X1 U1698 (.Y(n4360), 
	.B1(n7169), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6338));
   INVX1 U1699 (.Y(n7169), 
	.A(\ram[236][2] ));
   OAI22X1 U1700 (.Y(n4359), 
	.B1(n7170), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6306));
   INVX1 U1701 (.Y(n7170), 
	.A(\ram[236][1] ));
   OAI22X1 U1702 (.Y(n4358), 
	.B1(n7171), 
	.B0(n7155), 
	.A1(n7154), 
	.A0(n6309));
   INVX1 U1703 (.Y(n7171), 
	.A(\ram[236][0] ));
   NOR2BX1 U1704 (.Y(n7155), 
	.B(n7154), 
	.AN(mem_write_en));
   NAND2X1 U1705 (.Y(n7154), 
	.B(n6591), 
	.A(n7117));
   OAI22X1 U1706 (.Y(n4357), 
	.B1(n7174), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6311));
   INVX1 U1707 (.Y(n7174), 
	.A(\ram[235][15] ));
   OAI22X1 U1708 (.Y(n4356), 
	.B1(n7175), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6314));
   INVX1 U1709 (.Y(n7175), 
	.A(\ram[235][14] ));
   OAI22X1 U1710 (.Y(n4355), 
	.B1(n7176), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6316));
   INVX1 U1711 (.Y(n7176), 
	.A(\ram[235][13] ));
   OAI22X1 U1712 (.Y(n4354), 
	.B1(n7177), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6318));
   INVX1 U1713 (.Y(n7177), 
	.A(\ram[235][12] ));
   OAI22X1 U1714 (.Y(n4353), 
	.B1(n7178), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6320));
   INVX1 U1715 (.Y(n7178), 
	.A(\ram[235][11] ));
   OAI22X1 U1716 (.Y(n4352), 
	.B1(n7179), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6322));
   INVX1 U1717 (.Y(n7179), 
	.A(\ram[235][10] ));
   OAI22X1 U1718 (.Y(n4351), 
	.B1(n7180), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6324));
   INVX1 U1719 (.Y(n7180), 
	.A(\ram[235][9] ));
   OAI22X1 U1720 (.Y(n4350), 
	.B1(n7181), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6326));
   INVX1 U1721 (.Y(n7181), 
	.A(\ram[235][8] ));
   OAI22X1 U1722 (.Y(n4349), 
	.B1(n7182), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6328));
   INVX1 U1723 (.Y(n7182), 
	.A(\ram[235][7] ));
   OAI22X1 U1724 (.Y(n4348), 
	.B1(n7183), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6330));
   INVX1 U1725 (.Y(n7183), 
	.A(\ram[235][6] ));
   OAI22X1 U1726 (.Y(n4347), 
	.B1(n7184), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6332));
   INVX1 U1727 (.Y(n7184), 
	.A(\ram[235][5] ));
   OAI22X1 U1728 (.Y(n4346), 
	.B1(n7185), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6334));
   INVX1 U1729 (.Y(n7185), 
	.A(\ram[235][4] ));
   OAI22X1 U1730 (.Y(n4345), 
	.B1(n7186), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6336));
   INVX1 U1731 (.Y(n7186), 
	.A(\ram[235][3] ));
   OAI22X1 U1732 (.Y(n4344), 
	.B1(n7187), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6338));
   INVX1 U1733 (.Y(n7187), 
	.A(\ram[235][2] ));
   OAI22X1 U1734 (.Y(n4343), 
	.B1(n7188), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6306));
   INVX1 U1735 (.Y(n7188), 
	.A(\ram[235][1] ));
   OAI22X1 U1736 (.Y(n4342), 
	.B1(n7189), 
	.B0(n7173), 
	.A1(n7172), 
	.A0(n6309));
   INVX1 U1737 (.Y(n7189), 
	.A(\ram[235][0] ));
   NOR2BX1 U1738 (.Y(n7173), 
	.B(n7172), 
	.AN(mem_write_en));
   NAND2X1 U1739 (.Y(n7172), 
	.B(n6610), 
	.A(n7117));
   OAI22X1 U1740 (.Y(n4341), 
	.B1(n7192), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6311));
   INVX1 U1741 (.Y(n7192), 
	.A(\ram[234][15] ));
   OAI22X1 U1742 (.Y(n4340), 
	.B1(n7193), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6314));
   INVX1 U1743 (.Y(n7193), 
	.A(\ram[234][14] ));
   OAI22X1 U1744 (.Y(n4339), 
	.B1(n7194), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6316));
   INVX1 U1745 (.Y(n7194), 
	.A(\ram[234][13] ));
   OAI22X1 U1746 (.Y(n4338), 
	.B1(n7195), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6318));
   INVX1 U1747 (.Y(n7195), 
	.A(\ram[234][12] ));
   OAI22X1 U1748 (.Y(n4337), 
	.B1(n7196), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6320));
   INVX1 U1749 (.Y(n7196), 
	.A(\ram[234][11] ));
   OAI22X1 U1750 (.Y(n4336), 
	.B1(n7197), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6322));
   INVX1 U1751 (.Y(n7197), 
	.A(\ram[234][10] ));
   OAI22X1 U1752 (.Y(n4335), 
	.B1(n7198), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6324));
   INVX1 U1753 (.Y(n7198), 
	.A(\ram[234][9] ));
   OAI22X1 U1754 (.Y(n4334), 
	.B1(n7199), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6326));
   INVX1 U1755 (.Y(n7199), 
	.A(\ram[234][8] ));
   OAI22X1 U1756 (.Y(n4333), 
	.B1(n7200), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6328));
   INVX1 U1757 (.Y(n7200), 
	.A(\ram[234][7] ));
   OAI22X1 U1758 (.Y(n4332), 
	.B1(n7201), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6330));
   INVX1 U1759 (.Y(n7201), 
	.A(\ram[234][6] ));
   OAI22X1 U1760 (.Y(n4331), 
	.B1(n7202), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6332));
   INVX1 U1761 (.Y(n7202), 
	.A(\ram[234][5] ));
   OAI22X1 U1762 (.Y(n4330), 
	.B1(n7203), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6334));
   INVX1 U1763 (.Y(n7203), 
	.A(\ram[234][4] ));
   OAI22X1 U1764 (.Y(n4329), 
	.B1(n7204), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6336));
   INVX1 U1765 (.Y(n7204), 
	.A(\ram[234][3] ));
   OAI22X1 U1766 (.Y(n4328), 
	.B1(n7205), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6338));
   INVX1 U1767 (.Y(n7205), 
	.A(\ram[234][2] ));
   OAI22X1 U1768 (.Y(n4327), 
	.B1(n7206), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6306));
   INVX1 U1769 (.Y(n7206), 
	.A(\ram[234][1] ));
   OAI22X1 U1770 (.Y(n4326), 
	.B1(n7207), 
	.B0(n7191), 
	.A1(n7190), 
	.A0(n6309));
   INVX1 U1771 (.Y(n7207), 
	.A(\ram[234][0] ));
   NOR2BX1 U1772 (.Y(n7191), 
	.B(n7190), 
	.AN(mem_write_en));
   NAND2X1 U1773 (.Y(n7190), 
	.B(n6629), 
	.A(n7117));
   OAI22X1 U1774 (.Y(n4325), 
	.B1(n7210), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6311));
   INVX1 U1775 (.Y(n7210), 
	.A(\ram[233][15] ));
   OAI22X1 U1776 (.Y(n4324), 
	.B1(n7211), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6314));
   INVX1 U1777 (.Y(n7211), 
	.A(\ram[233][14] ));
   OAI22X1 U1778 (.Y(n4323), 
	.B1(n7212), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6316));
   INVX1 U1779 (.Y(n7212), 
	.A(\ram[233][13] ));
   OAI22X1 U1780 (.Y(n4322), 
	.B1(n7213), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6318));
   INVX1 U1781 (.Y(n7213), 
	.A(\ram[233][12] ));
   OAI22X1 U1782 (.Y(n4321), 
	.B1(n7214), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6320));
   INVX1 U1783 (.Y(n7214), 
	.A(\ram[233][11] ));
   OAI22X1 U1784 (.Y(n4320), 
	.B1(n7215), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6322));
   INVX1 U1785 (.Y(n7215), 
	.A(\ram[233][10] ));
   OAI22X1 U1786 (.Y(n4319), 
	.B1(n7216), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6324));
   INVX1 U1787 (.Y(n7216), 
	.A(\ram[233][9] ));
   OAI22X1 U1788 (.Y(n4318), 
	.B1(n7217), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6326));
   INVX1 U1789 (.Y(n7217), 
	.A(\ram[233][8] ));
   OAI22X1 U1790 (.Y(n4317), 
	.B1(n7218), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6328));
   INVX1 U1791 (.Y(n7218), 
	.A(\ram[233][7] ));
   OAI22X1 U1792 (.Y(n4316), 
	.B1(n7219), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6330));
   INVX1 U1793 (.Y(n7219), 
	.A(\ram[233][6] ));
   OAI22X1 U1794 (.Y(n4315), 
	.B1(n7220), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6332));
   INVX1 U1795 (.Y(n7220), 
	.A(\ram[233][5] ));
   OAI22X1 U1796 (.Y(n4314), 
	.B1(n7221), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6334));
   INVX1 U1797 (.Y(n7221), 
	.A(\ram[233][4] ));
   OAI22X1 U1798 (.Y(n4313), 
	.B1(n7222), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6336));
   INVX1 U1799 (.Y(n7222), 
	.A(\ram[233][3] ));
   OAI22X1 U1800 (.Y(n4312), 
	.B1(n7223), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6338));
   INVX1 U1801 (.Y(n7223), 
	.A(\ram[233][2] ));
   OAI22X1 U1802 (.Y(n4311), 
	.B1(n7224), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6306));
   INVX1 U1803 (.Y(n7224), 
	.A(\ram[233][1] ));
   OAI22X1 U1804 (.Y(n4310), 
	.B1(n7225), 
	.B0(n7209), 
	.A1(n7208), 
	.A0(n6309));
   INVX1 U1805 (.Y(n7225), 
	.A(\ram[233][0] ));
   NOR2BX1 U1806 (.Y(n7209), 
	.B(n7208), 
	.AN(mem_write_en));
   NAND2X1 U1807 (.Y(n7208), 
	.B(n6342), 
	.A(n7117));
   OAI22X1 U1808 (.Y(n4309), 
	.B1(n7228), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6311));
   INVX1 U1809 (.Y(n7228), 
	.A(\ram[232][15] ));
   OAI22X1 U1810 (.Y(n4308), 
	.B1(n7229), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6314));
   INVX1 U1811 (.Y(n7229), 
	.A(\ram[232][14] ));
   OAI22X1 U1812 (.Y(n4307), 
	.B1(n7230), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6316));
   INVX1 U1813 (.Y(n7230), 
	.A(\ram[232][13] ));
   OAI22X1 U1814 (.Y(n4306), 
	.B1(n7231), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6318));
   INVX1 U1815 (.Y(n7231), 
	.A(\ram[232][12] ));
   OAI22X1 U1816 (.Y(n4305), 
	.B1(n7232), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6320));
   INVX1 U1817 (.Y(n7232), 
	.A(\ram[232][11] ));
   OAI22X1 U1818 (.Y(n4304), 
	.B1(n7233), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6322));
   INVX1 U1819 (.Y(n7233), 
	.A(\ram[232][10] ));
   OAI22X1 U1820 (.Y(n4303), 
	.B1(n7234), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6324));
   INVX1 U1821 (.Y(n7234), 
	.A(\ram[232][9] ));
   OAI22X1 U1822 (.Y(n4302), 
	.B1(n7235), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6326));
   INVX1 U1823 (.Y(n7235), 
	.A(\ram[232][8] ));
   OAI22X1 U1824 (.Y(n4301), 
	.B1(n7236), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6328));
   INVX1 U1825 (.Y(n7236), 
	.A(\ram[232][7] ));
   OAI22X1 U1826 (.Y(n4300), 
	.B1(n7237), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6330));
   INVX1 U1827 (.Y(n7237), 
	.A(\ram[232][6] ));
   OAI22X1 U1828 (.Y(n4299), 
	.B1(n7238), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6332));
   INVX1 U1829 (.Y(n7238), 
	.A(\ram[232][5] ));
   OAI22X1 U1830 (.Y(n4298), 
	.B1(n7239), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6334));
   INVX1 U1831 (.Y(n7239), 
	.A(\ram[232][4] ));
   OAI22X1 U1832 (.Y(n4297), 
	.B1(n7240), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6336));
   INVX1 U1833 (.Y(n7240), 
	.A(\ram[232][3] ));
   OAI22X1 U1834 (.Y(n4296), 
	.B1(n7241), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6338));
   INVX1 U1835 (.Y(n7241), 
	.A(\ram[232][2] ));
   OAI22X1 U1836 (.Y(n4295), 
	.B1(n7242), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6306));
   INVX1 U1837 (.Y(n7242), 
	.A(\ram[232][1] ));
   OAI22X1 U1838 (.Y(n4294), 
	.B1(n7243), 
	.B0(n7227), 
	.A1(n7226), 
	.A0(n6309));
   INVX1 U1839 (.Y(n7243), 
	.A(\ram[232][0] ));
   NOR2BX1 U1840 (.Y(n7227), 
	.B(n7226), 
	.AN(mem_write_en));
   NAND2X1 U1841 (.Y(n7226), 
	.B(n6362), 
	.A(n7117));
   OAI22X1 U1842 (.Y(n4293), 
	.B1(n7246), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6311));
   INVX1 U1843 (.Y(n7246), 
	.A(\ram[231][15] ));
   OAI22X1 U1844 (.Y(n4292), 
	.B1(n7247), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6314));
   INVX1 U1845 (.Y(n7247), 
	.A(\ram[231][14] ));
   OAI22X1 U1846 (.Y(n4291), 
	.B1(n7248), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6316));
   INVX1 U1847 (.Y(n7248), 
	.A(\ram[231][13] ));
   OAI22X1 U1848 (.Y(n4290), 
	.B1(n7249), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6318));
   INVX1 U1849 (.Y(n7249), 
	.A(\ram[231][12] ));
   OAI22X1 U1850 (.Y(n4289), 
	.B1(n7250), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6320));
   INVX1 U1851 (.Y(n7250), 
	.A(\ram[231][11] ));
   OAI22X1 U1852 (.Y(n4288), 
	.B1(n7251), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6322));
   INVX1 U1853 (.Y(n7251), 
	.A(\ram[231][10] ));
   OAI22X1 U1854 (.Y(n4287), 
	.B1(n7252), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6324));
   INVX1 U1855 (.Y(n7252), 
	.A(\ram[231][9] ));
   OAI22X1 U1856 (.Y(n4286), 
	.B1(n7253), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6326));
   INVX1 U1857 (.Y(n7253), 
	.A(\ram[231][8] ));
   OAI22X1 U1858 (.Y(n4285), 
	.B1(n7254), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6328));
   INVX1 U1859 (.Y(n7254), 
	.A(\ram[231][7] ));
   OAI22X1 U1860 (.Y(n4284), 
	.B1(n7255), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6330));
   INVX1 U1861 (.Y(n7255), 
	.A(\ram[231][6] ));
   OAI22X1 U1862 (.Y(n4283), 
	.B1(n7256), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6332));
   INVX1 U1863 (.Y(n7256), 
	.A(\ram[231][5] ));
   OAI22X1 U1864 (.Y(n4282), 
	.B1(n7257), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6334));
   INVX1 U1865 (.Y(n7257), 
	.A(\ram[231][4] ));
   OAI22X1 U1866 (.Y(n4281), 
	.B1(n7258), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6336));
   INVX1 U1867 (.Y(n7258), 
	.A(\ram[231][3] ));
   OAI22X1 U1868 (.Y(n4280), 
	.B1(n7259), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6338));
   INVX1 U1869 (.Y(n7259), 
	.A(\ram[231][2] ));
   OAI22X1 U1870 (.Y(n4279), 
	.B1(n7260), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6306));
   INVX1 U1871 (.Y(n7260), 
	.A(\ram[231][1] ));
   OAI22X1 U1872 (.Y(n4278), 
	.B1(n7261), 
	.B0(n7245), 
	.A1(n7244), 
	.A0(n6309));
   INVX1 U1873 (.Y(n7261), 
	.A(\ram[231][0] ));
   NOR2BX1 U1874 (.Y(n7245), 
	.B(n7244), 
	.AN(mem_write_en));
   NAND2X1 U1875 (.Y(n7244), 
	.B(n6381), 
	.A(n7117));
   OAI22X1 U1876 (.Y(n4277), 
	.B1(n7264), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6311));
   INVX1 U1877 (.Y(n7264), 
	.A(\ram[230][15] ));
   OAI22X1 U1878 (.Y(n4276), 
	.B1(n7265), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6314));
   INVX1 U1879 (.Y(n7265), 
	.A(\ram[230][14] ));
   OAI22X1 U1880 (.Y(n4275), 
	.B1(n7266), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6316));
   INVX1 U1881 (.Y(n7266), 
	.A(\ram[230][13] ));
   OAI22X1 U1882 (.Y(n4274), 
	.B1(n7267), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6318));
   INVX1 U1883 (.Y(n7267), 
	.A(\ram[230][12] ));
   OAI22X1 U1884 (.Y(n4273), 
	.B1(n7268), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6320));
   INVX1 U1885 (.Y(n7268), 
	.A(\ram[230][11] ));
   OAI22X1 U1886 (.Y(n4272), 
	.B1(n7269), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6322));
   INVX1 U1887 (.Y(n7269), 
	.A(\ram[230][10] ));
   OAI22X1 U1888 (.Y(n4271), 
	.B1(n7270), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6324));
   INVX1 U1889 (.Y(n7270), 
	.A(\ram[230][9] ));
   OAI22X1 U1890 (.Y(n4270), 
	.B1(n7271), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6326));
   INVX1 U1891 (.Y(n7271), 
	.A(\ram[230][8] ));
   OAI22X1 U1892 (.Y(n4269), 
	.B1(n7272), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6328));
   INVX1 U1893 (.Y(n7272), 
	.A(\ram[230][7] ));
   OAI22X1 U1894 (.Y(n4268), 
	.B1(n7273), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6330));
   INVX1 U1895 (.Y(n7273), 
	.A(\ram[230][6] ));
   OAI22X1 U1896 (.Y(n4267), 
	.B1(n7274), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6332));
   INVX1 U1897 (.Y(n7274), 
	.A(\ram[230][5] ));
   OAI22X1 U1898 (.Y(n4266), 
	.B1(n7275), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6334));
   INVX1 U1899 (.Y(n7275), 
	.A(\ram[230][4] ));
   OAI22X1 U1900 (.Y(n4265), 
	.B1(n7276), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6336));
   INVX1 U1901 (.Y(n7276), 
	.A(\ram[230][3] ));
   OAI22X1 U1902 (.Y(n4264), 
	.B1(n7277), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6338));
   INVX1 U1903 (.Y(n7277), 
	.A(\ram[230][2] ));
   OAI22X1 U1904 (.Y(n4263), 
	.B1(n7278), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6306));
   INVX1 U1905 (.Y(n7278), 
	.A(\ram[230][1] ));
   OAI22X1 U1906 (.Y(n4262), 
	.B1(n7279), 
	.B0(n7263), 
	.A1(n7262), 
	.A0(n6309));
   INVX1 U1907 (.Y(n7279), 
	.A(\ram[230][0] ));
   NOR2BX1 U1908 (.Y(n7263), 
	.B(n7262), 
	.AN(mem_write_en));
   NAND2X1 U1909 (.Y(n7262), 
	.B(n6400), 
	.A(n7117));
   OAI22X1 U1910 (.Y(n4261), 
	.B1(n7282), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6311));
   INVX1 U1911 (.Y(n7282), 
	.A(\ram[229][15] ));
   OAI22X1 U1912 (.Y(n4260), 
	.B1(n7283), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6314));
   INVX1 U1913 (.Y(n7283), 
	.A(\ram[229][14] ));
   OAI22X1 U1914 (.Y(n4259), 
	.B1(n7284), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6316));
   INVX1 U1915 (.Y(n7284), 
	.A(\ram[229][13] ));
   OAI22X1 U1916 (.Y(n4258), 
	.B1(n7285), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6318));
   INVX1 U1917 (.Y(n7285), 
	.A(\ram[229][12] ));
   OAI22X1 U1918 (.Y(n4257), 
	.B1(n7286), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6320));
   INVX1 U1919 (.Y(n7286), 
	.A(\ram[229][11] ));
   OAI22X1 U1920 (.Y(n4256), 
	.B1(n7287), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6322));
   INVX1 U1921 (.Y(n7287), 
	.A(\ram[229][10] ));
   OAI22X1 U1922 (.Y(n4255), 
	.B1(n7288), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6324));
   INVX1 U1923 (.Y(n7288), 
	.A(\ram[229][9] ));
   OAI22X1 U1924 (.Y(n4254), 
	.B1(n7289), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6326));
   INVX1 U1925 (.Y(n7289), 
	.A(\ram[229][8] ));
   OAI22X1 U1926 (.Y(n4253), 
	.B1(n7290), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6328));
   INVX1 U1927 (.Y(n7290), 
	.A(\ram[229][7] ));
   OAI22X1 U1928 (.Y(n4252), 
	.B1(n7291), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6330));
   INVX1 U1929 (.Y(n7291), 
	.A(\ram[229][6] ));
   OAI22X1 U1930 (.Y(n4251), 
	.B1(n7292), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6332));
   INVX1 U1931 (.Y(n7292), 
	.A(\ram[229][5] ));
   OAI22X1 U1932 (.Y(n4250), 
	.B1(n7293), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6334));
   INVX1 U1933 (.Y(n7293), 
	.A(\ram[229][4] ));
   OAI22X1 U1934 (.Y(n4249), 
	.B1(n7294), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6336));
   INVX1 U1935 (.Y(n7294), 
	.A(\ram[229][3] ));
   OAI22X1 U1936 (.Y(n4248), 
	.B1(n7295), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6338));
   INVX1 U1937 (.Y(n7295), 
	.A(\ram[229][2] ));
   OAI22X1 U1938 (.Y(n4247), 
	.B1(n7296), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6306));
   INVX1 U1939 (.Y(n7296), 
	.A(\ram[229][1] ));
   OAI22X1 U1940 (.Y(n4246), 
	.B1(n7297), 
	.B0(n7281), 
	.A1(n7280), 
	.A0(n6309));
   INVX1 U1941 (.Y(n7297), 
	.A(\ram[229][0] ));
   NOR2BX1 U1942 (.Y(n7281), 
	.B(n7280), 
	.AN(mem_write_en));
   NAND2X1 U1943 (.Y(n7280), 
	.B(n6419), 
	.A(n7117));
   OAI22X1 U1944 (.Y(n4245), 
	.B1(n7300), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6311));
   INVX1 U1945 (.Y(n7300), 
	.A(\ram[228][15] ));
   OAI22X1 U1946 (.Y(n4244), 
	.B1(n7301), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6314));
   INVX1 U1947 (.Y(n7301), 
	.A(\ram[228][14] ));
   OAI22X1 U1948 (.Y(n4243), 
	.B1(n7302), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6316));
   INVX1 U1949 (.Y(n7302), 
	.A(\ram[228][13] ));
   OAI22X1 U1950 (.Y(n4242), 
	.B1(n7303), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6318));
   INVX1 U1951 (.Y(n7303), 
	.A(\ram[228][12] ));
   OAI22X1 U1952 (.Y(n4241), 
	.B1(n7304), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6320));
   INVX1 U1953 (.Y(n7304), 
	.A(\ram[228][11] ));
   OAI22X1 U1954 (.Y(n4240), 
	.B1(n7305), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6322));
   INVX1 U1955 (.Y(n7305), 
	.A(\ram[228][10] ));
   OAI22X1 U1956 (.Y(n4239), 
	.B1(n7306), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6324));
   INVX1 U1957 (.Y(n7306), 
	.A(\ram[228][9] ));
   OAI22X1 U1958 (.Y(n4238), 
	.B1(n7307), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6326));
   INVX1 U1959 (.Y(n7307), 
	.A(\ram[228][8] ));
   OAI22X1 U1960 (.Y(n4237), 
	.B1(n7308), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6328));
   INVX1 U1961 (.Y(n7308), 
	.A(\ram[228][7] ));
   OAI22X1 U1962 (.Y(n4236), 
	.B1(n7309), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6330));
   INVX1 U1963 (.Y(n7309), 
	.A(\ram[228][6] ));
   OAI22X1 U1964 (.Y(n4235), 
	.B1(n7310), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6332));
   INVX1 U1965 (.Y(n7310), 
	.A(\ram[228][5] ));
   OAI22X1 U1966 (.Y(n4234), 
	.B1(n7311), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6334));
   INVX1 U1967 (.Y(n7311), 
	.A(\ram[228][4] ));
   OAI22X1 U1968 (.Y(n4233), 
	.B1(n7312), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6336));
   INVX1 U1969 (.Y(n7312), 
	.A(\ram[228][3] ));
   OAI22X1 U1970 (.Y(n4232), 
	.B1(n7313), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6338));
   INVX1 U1971 (.Y(n7313), 
	.A(\ram[228][2] ));
   OAI22X1 U1972 (.Y(n4231), 
	.B1(n7314), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6306));
   INVX1 U1973 (.Y(n7314), 
	.A(\ram[228][1] ));
   OAI22X1 U1974 (.Y(n4230), 
	.B1(n7315), 
	.B0(n7299), 
	.A1(n7298), 
	.A0(n6309));
   INVX1 U1975 (.Y(n7315), 
	.A(\ram[228][0] ));
   NOR2BX1 U1976 (.Y(n7299), 
	.B(n7298), 
	.AN(mem_write_en));
   NAND2X1 U1977 (.Y(n7298), 
	.B(n6438), 
	.A(n7117));
   OAI22X1 U1978 (.Y(n4229), 
	.B1(n7318), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6311));
   INVX1 U1979 (.Y(n7318), 
	.A(\ram[227][15] ));
   OAI22X1 U1980 (.Y(n4228), 
	.B1(n7319), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6314));
   INVX1 U1981 (.Y(n7319), 
	.A(\ram[227][14] ));
   OAI22X1 U1982 (.Y(n4227), 
	.B1(n7320), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6316));
   INVX1 U1983 (.Y(n7320), 
	.A(\ram[227][13] ));
   OAI22X1 U1984 (.Y(n4226), 
	.B1(n7321), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6318));
   INVX1 U1985 (.Y(n7321), 
	.A(\ram[227][12] ));
   OAI22X1 U1986 (.Y(n4225), 
	.B1(n7322), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6320));
   INVX1 U1987 (.Y(n7322), 
	.A(\ram[227][11] ));
   OAI22X1 U1988 (.Y(n4224), 
	.B1(n7323), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6322));
   INVX1 U1989 (.Y(n7323), 
	.A(\ram[227][10] ));
   OAI22X1 U1990 (.Y(n4223), 
	.B1(n7324), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6324));
   INVX1 U1991 (.Y(n7324), 
	.A(\ram[227][9] ));
   OAI22X1 U1992 (.Y(n4222), 
	.B1(n7325), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6326));
   INVX1 U1993 (.Y(n7325), 
	.A(\ram[227][8] ));
   OAI22X1 U1994 (.Y(n4221), 
	.B1(n7326), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6328));
   INVX1 U1995 (.Y(n7326), 
	.A(\ram[227][7] ));
   OAI22X1 U1996 (.Y(n4220), 
	.B1(n7327), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6330));
   INVX1 U1997 (.Y(n7327), 
	.A(\ram[227][6] ));
   OAI22X1 U1998 (.Y(n4219), 
	.B1(n7328), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6332));
   INVX1 U1999 (.Y(n7328), 
	.A(\ram[227][5] ));
   OAI22X1 U2000 (.Y(n4218), 
	.B1(n7329), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6334));
   INVX1 U2001 (.Y(n7329), 
	.A(\ram[227][4] ));
   OAI22X1 U2002 (.Y(n4217), 
	.B1(n7330), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6336));
   INVX1 U2003 (.Y(n7330), 
	.A(\ram[227][3] ));
   OAI22X1 U2004 (.Y(n4216), 
	.B1(n7331), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6338));
   INVX1 U2005 (.Y(n7331), 
	.A(\ram[227][2] ));
   OAI22X1 U2006 (.Y(n4215), 
	.B1(n7332), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6306));
   INVX1 U2007 (.Y(n7332), 
	.A(\ram[227][1] ));
   OAI22X1 U2008 (.Y(n4214), 
	.B1(n7333), 
	.B0(n7317), 
	.A1(n7316), 
	.A0(n6309));
   INVX1 U2009 (.Y(n7333), 
	.A(\ram[227][0] ));
   NOR2BX1 U2010 (.Y(n7317), 
	.B(n7316), 
	.AN(mem_write_en));
   NAND2X1 U2011 (.Y(n7316), 
	.B(n6457), 
	.A(n7117));
   OAI22X1 U2012 (.Y(n4213), 
	.B1(n7336), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6311));
   INVX1 U2013 (.Y(n7336), 
	.A(\ram[226][15] ));
   OAI22X1 U2014 (.Y(n4212), 
	.B1(n7337), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6314));
   INVX1 U2015 (.Y(n7337), 
	.A(\ram[226][14] ));
   OAI22X1 U2016 (.Y(n4211), 
	.B1(n7338), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6316));
   INVX1 U2017 (.Y(n7338), 
	.A(\ram[226][13] ));
   OAI22X1 U2018 (.Y(n4210), 
	.B1(n7339), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6318));
   INVX1 U2019 (.Y(n7339), 
	.A(\ram[226][12] ));
   OAI22X1 U2020 (.Y(n4209), 
	.B1(n7340), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6320));
   INVX1 U2021 (.Y(n7340), 
	.A(\ram[226][11] ));
   OAI22X1 U2022 (.Y(n4208), 
	.B1(n7341), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6322));
   INVX1 U2023 (.Y(n7341), 
	.A(\ram[226][10] ));
   OAI22X1 U2024 (.Y(n4207), 
	.B1(n7342), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6324));
   INVX1 U2025 (.Y(n7342), 
	.A(\ram[226][9] ));
   OAI22X1 U2026 (.Y(n4206), 
	.B1(n7343), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6326));
   INVX1 U2027 (.Y(n7343), 
	.A(\ram[226][8] ));
   OAI22X1 U2028 (.Y(n4205), 
	.B1(n7344), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6328));
   INVX1 U2029 (.Y(n7344), 
	.A(\ram[226][7] ));
   OAI22X1 U2030 (.Y(n4204), 
	.B1(n7345), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6330));
   INVX1 U2031 (.Y(n7345), 
	.A(\ram[226][6] ));
   OAI22X1 U2032 (.Y(n4203), 
	.B1(n7346), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6332));
   INVX1 U2033 (.Y(n7346), 
	.A(\ram[226][5] ));
   OAI22X1 U2034 (.Y(n4202), 
	.B1(n7347), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6334));
   INVX1 U2035 (.Y(n7347), 
	.A(\ram[226][4] ));
   OAI22X1 U2036 (.Y(n4201), 
	.B1(n7348), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6336));
   INVX1 U2037 (.Y(n7348), 
	.A(\ram[226][3] ));
   OAI22X1 U2038 (.Y(n4200), 
	.B1(n7349), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6338));
   INVX1 U2039 (.Y(n7349), 
	.A(\ram[226][2] ));
   OAI22X1 U2040 (.Y(n4199), 
	.B1(n7350), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6306));
   INVX1 U2041 (.Y(n7350), 
	.A(\ram[226][1] ));
   OAI22X1 U2042 (.Y(n4198), 
	.B1(n7351), 
	.B0(n7335), 
	.A1(n7334), 
	.A0(n6309));
   INVX1 U2043 (.Y(n7351), 
	.A(\ram[226][0] ));
   NOR2BX1 U2044 (.Y(n7335), 
	.B(n7334), 
	.AN(mem_write_en));
   NAND2X1 U2045 (.Y(n7334), 
	.B(n6476), 
	.A(n7117));
   OAI22X1 U2046 (.Y(n4197), 
	.B1(n7354), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6311));
   INVX1 U2047 (.Y(n7354), 
	.A(\ram[225][15] ));
   OAI22X1 U2048 (.Y(n4196), 
	.B1(n7355), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6314));
   INVX1 U2049 (.Y(n7355), 
	.A(\ram[225][14] ));
   OAI22X1 U2050 (.Y(n4195), 
	.B1(n7356), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6316));
   INVX1 U2051 (.Y(n7356), 
	.A(\ram[225][13] ));
   OAI22X1 U2052 (.Y(n4194), 
	.B1(n7357), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6318));
   INVX1 U2053 (.Y(n7357), 
	.A(\ram[225][12] ));
   OAI22X1 U2054 (.Y(n4193), 
	.B1(n7358), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6320));
   INVX1 U2055 (.Y(n7358), 
	.A(\ram[225][11] ));
   OAI22X1 U2056 (.Y(n4192), 
	.B1(n7359), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6322));
   INVX1 U2057 (.Y(n7359), 
	.A(\ram[225][10] ));
   OAI22X1 U2058 (.Y(n4191), 
	.B1(n7360), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6324));
   INVX1 U2059 (.Y(n7360), 
	.A(\ram[225][9] ));
   OAI22X1 U2060 (.Y(n4190), 
	.B1(n7361), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6326));
   INVX1 U2061 (.Y(n7361), 
	.A(\ram[225][8] ));
   OAI22X1 U2062 (.Y(n4189), 
	.B1(n7362), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6328));
   INVX1 U2063 (.Y(n7362), 
	.A(\ram[225][7] ));
   OAI22X1 U2064 (.Y(n4188), 
	.B1(n7363), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6330));
   INVX1 U2065 (.Y(n7363), 
	.A(\ram[225][6] ));
   OAI22X1 U2066 (.Y(n4187), 
	.B1(n7364), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6332));
   INVX1 U2067 (.Y(n7364), 
	.A(\ram[225][5] ));
   OAI22X1 U2068 (.Y(n4186), 
	.B1(n7365), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6334));
   INVX1 U2069 (.Y(n7365), 
	.A(\ram[225][4] ));
   OAI22X1 U2070 (.Y(n4185), 
	.B1(n7366), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6336));
   INVX1 U2071 (.Y(n7366), 
	.A(\ram[225][3] ));
   OAI22X1 U2072 (.Y(n4184), 
	.B1(n7367), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6338));
   INVX1 U2073 (.Y(n7367), 
	.A(\ram[225][2] ));
   OAI22X1 U2074 (.Y(n4183), 
	.B1(n7368), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6306));
   INVX1 U2075 (.Y(n7368), 
	.A(\ram[225][1] ));
   OAI22X1 U2076 (.Y(n4182), 
	.B1(n7369), 
	.B0(n7353), 
	.A1(n7352), 
	.A0(n6309));
   INVX1 U2077 (.Y(n7369), 
	.A(\ram[225][0] ));
   NOR2BX1 U2078 (.Y(n7353), 
	.B(n7352), 
	.AN(mem_write_en));
   NAND2X1 U2079 (.Y(n7352), 
	.B(n6495), 
	.A(n7117));
   OAI22X1 U2080 (.Y(n4181), 
	.B1(n7372), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6311));
   INVX1 U2081 (.Y(n7372), 
	.A(\ram[224][15] ));
   OAI22X1 U2082 (.Y(n4180), 
	.B1(n7373), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6314));
   INVX1 U2083 (.Y(n7373), 
	.A(\ram[224][14] ));
   OAI22X1 U2084 (.Y(n4179), 
	.B1(n7374), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6316));
   INVX1 U2085 (.Y(n7374), 
	.A(\ram[224][13] ));
   OAI22X1 U2086 (.Y(n4178), 
	.B1(n7375), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6318));
   INVX1 U2087 (.Y(n7375), 
	.A(\ram[224][12] ));
   OAI22X1 U2088 (.Y(n4177), 
	.B1(n7376), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6320));
   INVX1 U2089 (.Y(n7376), 
	.A(\ram[224][11] ));
   OAI22X1 U2090 (.Y(n4176), 
	.B1(n7377), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6322));
   INVX1 U2091 (.Y(n7377), 
	.A(\ram[224][10] ));
   OAI22X1 U2092 (.Y(n4175), 
	.B1(n7378), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6324));
   INVX1 U2093 (.Y(n7378), 
	.A(\ram[224][9] ));
   OAI22X1 U2094 (.Y(n4174), 
	.B1(n7379), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6326));
   INVX1 U2095 (.Y(n7379), 
	.A(\ram[224][8] ));
   OAI22X1 U2096 (.Y(n4173), 
	.B1(n7380), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6328));
   INVX1 U2097 (.Y(n7380), 
	.A(\ram[224][7] ));
   OAI22X1 U2098 (.Y(n4172), 
	.B1(n7381), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6330));
   INVX1 U2099 (.Y(n7381), 
	.A(\ram[224][6] ));
   OAI22X1 U2100 (.Y(n4171), 
	.B1(n7382), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6332));
   INVX1 U2101 (.Y(n7382), 
	.A(\ram[224][5] ));
   OAI22X1 U2102 (.Y(n4170), 
	.B1(n7383), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6334));
   INVX1 U2103 (.Y(n7383), 
	.A(\ram[224][4] ));
   OAI22X1 U2104 (.Y(n4169), 
	.B1(n7384), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6336));
   INVX1 U2105 (.Y(n7384), 
	.A(\ram[224][3] ));
   OAI22X1 U2106 (.Y(n4168), 
	.B1(n7385), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6338));
   INVX1 U2107 (.Y(n7385), 
	.A(\ram[224][2] ));
   OAI22X1 U2108 (.Y(n4167), 
	.B1(n7386), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6306));
   INVX1 U2109 (.Y(n7386), 
	.A(\ram[224][1] ));
   OAI22X1 U2110 (.Y(n4166), 
	.B1(n7387), 
	.B0(n7371), 
	.A1(n7370), 
	.A0(n6309));
   INVX1 U2111 (.Y(n7387), 
	.A(\ram[224][0] ));
   NOR2BX1 U2112 (.Y(n7371), 
	.B(n7370), 
	.AN(mem_write_en));
   NAND2X1 U2113 (.Y(n7370), 
	.B(n6514), 
	.A(n7117));
   OAI22X1 U2114 (.Y(n4165), 
	.B1(n7390), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6311));
   INVX1 U2115 (.Y(n7390), 
	.A(\ram[223][15] ));
   OAI22X1 U2116 (.Y(n4164), 
	.B1(n7391), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6314));
   INVX1 U2117 (.Y(n7391), 
	.A(\ram[223][14] ));
   OAI22X1 U2118 (.Y(n4163), 
	.B1(n7392), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6316));
   INVX1 U2119 (.Y(n7392), 
	.A(\ram[223][13] ));
   OAI22X1 U2120 (.Y(n4162), 
	.B1(n7393), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6318));
   INVX1 U2121 (.Y(n7393), 
	.A(\ram[223][12] ));
   OAI22X1 U2122 (.Y(n4161), 
	.B1(n7394), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6320));
   INVX1 U2123 (.Y(n7394), 
	.A(\ram[223][11] ));
   OAI22X1 U2124 (.Y(n4160), 
	.B1(n7395), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6322));
   INVX1 U2125 (.Y(n7395), 
	.A(\ram[223][10] ));
   OAI22X1 U2126 (.Y(n4159), 
	.B1(n7396), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6324));
   INVX1 U2127 (.Y(n7396), 
	.A(\ram[223][9] ));
   OAI22X1 U2128 (.Y(n4158), 
	.B1(n7397), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6326));
   INVX1 U2129 (.Y(n7397), 
	.A(\ram[223][8] ));
   OAI22X1 U2130 (.Y(n4157), 
	.B1(n7398), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6328));
   INVX1 U2131 (.Y(n7398), 
	.A(\ram[223][7] ));
   OAI22X1 U2132 (.Y(n4156), 
	.B1(n7399), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6330));
   INVX1 U2133 (.Y(n7399), 
	.A(\ram[223][6] ));
   OAI22X1 U2134 (.Y(n4155), 
	.B1(n7400), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6332));
   INVX1 U2135 (.Y(n7400), 
	.A(\ram[223][5] ));
   OAI22X1 U2136 (.Y(n4154), 
	.B1(n7401), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6334));
   INVX1 U2137 (.Y(n7401), 
	.A(\ram[223][4] ));
   OAI22X1 U2138 (.Y(n4153), 
	.B1(n7402), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6336));
   INVX1 U2139 (.Y(n7402), 
	.A(\ram[223][3] ));
   OAI22X1 U2140 (.Y(n4152), 
	.B1(n7403), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6338));
   INVX1 U2141 (.Y(n7403), 
	.A(\ram[223][2] ));
   OAI22X1 U2142 (.Y(n4151), 
	.B1(n7404), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6306));
   INVX1 U2143 (.Y(n7404), 
	.A(\ram[223][1] ));
   OAI22X1 U2144 (.Y(n4150), 
	.B1(n7405), 
	.B0(n7389), 
	.A1(n7388), 
	.A0(n6309));
   INVX1 U2145 (.Y(n7405), 
	.A(\ram[223][0] ));
   NOR2BX1 U2146 (.Y(n7389), 
	.B(n7388), 
	.AN(mem_write_en));
   NAND2X1 U2147 (.Y(n7388), 
	.B(n6533), 
	.A(n7406));
   OAI22X1 U2148 (.Y(n4149), 
	.B1(n7409), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6311));
   INVX1 U2149 (.Y(n7409), 
	.A(\ram[222][15] ));
   OAI22X1 U2150 (.Y(n4148), 
	.B1(n7410), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6314));
   INVX1 U2151 (.Y(n7410), 
	.A(\ram[222][14] ));
   OAI22X1 U2152 (.Y(n4147), 
	.B1(n7411), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6316));
   INVX1 U2153 (.Y(n7411), 
	.A(\ram[222][13] ));
   OAI22X1 U2154 (.Y(n4146), 
	.B1(n7412), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6318));
   INVX1 U2155 (.Y(n7412), 
	.A(\ram[222][12] ));
   OAI22X1 U2156 (.Y(n4145), 
	.B1(n7413), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6320));
   INVX1 U2157 (.Y(n7413), 
	.A(\ram[222][11] ));
   OAI22X1 U2158 (.Y(n4144), 
	.B1(n7414), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6322));
   INVX1 U2159 (.Y(n7414), 
	.A(\ram[222][10] ));
   OAI22X1 U2160 (.Y(n4143), 
	.B1(n7415), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6324));
   INVX1 U2161 (.Y(n7415), 
	.A(\ram[222][9] ));
   OAI22X1 U2162 (.Y(n4142), 
	.B1(n7416), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6326));
   INVX1 U2163 (.Y(n7416), 
	.A(\ram[222][8] ));
   OAI22X1 U2164 (.Y(n4141), 
	.B1(n7417), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6328));
   INVX1 U2165 (.Y(n7417), 
	.A(\ram[222][7] ));
   OAI22X1 U2166 (.Y(n4140), 
	.B1(n7418), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6330));
   INVX1 U2167 (.Y(n7418), 
	.A(\ram[222][6] ));
   OAI22X1 U2168 (.Y(n4139), 
	.B1(n7419), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6332));
   INVX1 U2169 (.Y(n7419), 
	.A(\ram[222][5] ));
   OAI22X1 U2170 (.Y(n4138), 
	.B1(n7420), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6334));
   INVX1 U2171 (.Y(n7420), 
	.A(\ram[222][4] ));
   OAI22X1 U2172 (.Y(n4137), 
	.B1(n7421), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6336));
   INVX1 U2173 (.Y(n7421), 
	.A(\ram[222][3] ));
   OAI22X1 U2174 (.Y(n4136), 
	.B1(n7422), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6338));
   INVX1 U2175 (.Y(n7422), 
	.A(\ram[222][2] ));
   OAI22X1 U2176 (.Y(n4135), 
	.B1(n7423), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6306));
   INVX1 U2177 (.Y(n7423), 
	.A(\ram[222][1] ));
   OAI22X1 U2178 (.Y(n4134), 
	.B1(n7424), 
	.B0(n7408), 
	.A1(n7407), 
	.A0(n6309));
   INVX1 U2179 (.Y(n7424), 
	.A(\ram[222][0] ));
   NOR2BX1 U2180 (.Y(n7408), 
	.B(n7407), 
	.AN(mem_write_en));
   NAND2X1 U2181 (.Y(n7407), 
	.B(n6553), 
	.A(n7406));
   OAI22X1 U2182 (.Y(n4133), 
	.B1(n7427), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6311));
   INVX1 U2183 (.Y(n7427), 
	.A(\ram[221][15] ));
   OAI22X1 U2184 (.Y(n4132), 
	.B1(n7428), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6314));
   INVX1 U2185 (.Y(n7428), 
	.A(\ram[221][14] ));
   OAI22X1 U2186 (.Y(n4131), 
	.B1(n7429), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6316));
   INVX1 U2187 (.Y(n7429), 
	.A(\ram[221][13] ));
   OAI22X1 U2188 (.Y(n4130), 
	.B1(n7430), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6318));
   INVX1 U2189 (.Y(n7430), 
	.A(\ram[221][12] ));
   OAI22X1 U2190 (.Y(n4129), 
	.B1(n7431), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6320));
   INVX1 U2191 (.Y(n7431), 
	.A(\ram[221][11] ));
   OAI22X1 U2192 (.Y(n4128), 
	.B1(n7432), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6322));
   INVX1 U2193 (.Y(n7432), 
	.A(\ram[221][10] ));
   OAI22X1 U2194 (.Y(n4127), 
	.B1(n7433), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6324));
   INVX1 U2195 (.Y(n7433), 
	.A(\ram[221][9] ));
   OAI22X1 U2196 (.Y(n4126), 
	.B1(n7434), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6326));
   INVX1 U2197 (.Y(n7434), 
	.A(\ram[221][8] ));
   OAI22X1 U2198 (.Y(n4125), 
	.B1(n7435), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6328));
   INVX1 U2199 (.Y(n7435), 
	.A(\ram[221][7] ));
   OAI22X1 U2200 (.Y(n4124), 
	.B1(n7436), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6330));
   INVX1 U2201 (.Y(n7436), 
	.A(\ram[221][6] ));
   OAI22X1 U2202 (.Y(n4123), 
	.B1(n7437), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6332));
   INVX1 U2203 (.Y(n7437), 
	.A(\ram[221][5] ));
   OAI22X1 U2204 (.Y(n4122), 
	.B1(n7438), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6334));
   INVX1 U2205 (.Y(n7438), 
	.A(\ram[221][4] ));
   OAI22X1 U2206 (.Y(n4121), 
	.B1(n7439), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6336));
   INVX1 U2207 (.Y(n7439), 
	.A(\ram[221][3] ));
   OAI22X1 U2208 (.Y(n4120), 
	.B1(n7440), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6338));
   INVX1 U2209 (.Y(n7440), 
	.A(\ram[221][2] ));
   OAI22X1 U2210 (.Y(n4119), 
	.B1(n7441), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6306));
   INVX1 U2211 (.Y(n7441), 
	.A(\ram[221][1] ));
   OAI22X1 U2212 (.Y(n4118), 
	.B1(n7442), 
	.B0(n7426), 
	.A1(n7425), 
	.A0(n6309));
   INVX1 U2213 (.Y(n7442), 
	.A(\ram[221][0] ));
   NOR2BX1 U2214 (.Y(n7426), 
	.B(n7425), 
	.AN(mem_write_en));
   NAND2X1 U2215 (.Y(n7425), 
	.B(n6572), 
	.A(n7406));
   OAI22X1 U2216 (.Y(n4117), 
	.B1(n7445), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6311));
   INVX1 U2217 (.Y(n7445), 
	.A(\ram[220][15] ));
   OAI22X1 U2218 (.Y(n4116), 
	.B1(n7446), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6314));
   INVX1 U2219 (.Y(n7446), 
	.A(\ram[220][14] ));
   OAI22X1 U2220 (.Y(n4115), 
	.B1(n7447), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6316));
   INVX1 U2221 (.Y(n7447), 
	.A(\ram[220][13] ));
   OAI22X1 U2222 (.Y(n4114), 
	.B1(n7448), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6318));
   INVX1 U2223 (.Y(n7448), 
	.A(\ram[220][12] ));
   OAI22X1 U2224 (.Y(n4113), 
	.B1(n7449), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6320));
   INVX1 U2225 (.Y(n7449), 
	.A(\ram[220][11] ));
   OAI22X1 U2226 (.Y(n4112), 
	.B1(n7450), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6322));
   INVX1 U2227 (.Y(n7450), 
	.A(\ram[220][10] ));
   OAI22X1 U2228 (.Y(n4111), 
	.B1(n7451), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6324));
   INVX1 U2229 (.Y(n7451), 
	.A(\ram[220][9] ));
   OAI22X1 U2230 (.Y(n4110), 
	.B1(n7452), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6326));
   INVX1 U2231 (.Y(n7452), 
	.A(\ram[220][8] ));
   OAI22X1 U2232 (.Y(n4109), 
	.B1(n7453), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6328));
   INVX1 U2233 (.Y(n7453), 
	.A(\ram[220][7] ));
   OAI22X1 U2234 (.Y(n4108), 
	.B1(n7454), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6330));
   INVX1 U2235 (.Y(n7454), 
	.A(\ram[220][6] ));
   OAI22X1 U2236 (.Y(n4107), 
	.B1(n7455), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6332));
   INVX1 U2237 (.Y(n7455), 
	.A(\ram[220][5] ));
   OAI22X1 U2238 (.Y(n4106), 
	.B1(n7456), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6334));
   INVX1 U2239 (.Y(n7456), 
	.A(\ram[220][4] ));
   OAI22X1 U2240 (.Y(n4105), 
	.B1(n7457), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6336));
   INVX1 U2241 (.Y(n7457), 
	.A(\ram[220][3] ));
   OAI22X1 U2242 (.Y(n4104), 
	.B1(n7458), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6338));
   INVX1 U2243 (.Y(n7458), 
	.A(\ram[220][2] ));
   OAI22X1 U2244 (.Y(n4103), 
	.B1(n7459), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6306));
   INVX1 U2245 (.Y(n7459), 
	.A(\ram[220][1] ));
   OAI22X1 U2246 (.Y(n4102), 
	.B1(n7460), 
	.B0(n7444), 
	.A1(n7443), 
	.A0(n6309));
   INVX1 U2247 (.Y(n7460), 
	.A(\ram[220][0] ));
   NOR2BX1 U2248 (.Y(n7444), 
	.B(n7443), 
	.AN(mem_write_en));
   NAND2X1 U2249 (.Y(n7443), 
	.B(n6591), 
	.A(n7406));
   OAI22X1 U2250 (.Y(n4101), 
	.B1(n7463), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6311));
   INVX1 U2251 (.Y(n7463), 
	.A(\ram[219][15] ));
   OAI22X1 U2252 (.Y(n4100), 
	.B1(n7464), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6314));
   INVX1 U2253 (.Y(n7464), 
	.A(\ram[219][14] ));
   OAI22X1 U2254 (.Y(n4099), 
	.B1(n7465), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6316));
   INVX1 U2255 (.Y(n7465), 
	.A(\ram[219][13] ));
   OAI22X1 U2256 (.Y(n4098), 
	.B1(n7466), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6318));
   INVX1 U2257 (.Y(n7466), 
	.A(\ram[219][12] ));
   OAI22X1 U2258 (.Y(n4097), 
	.B1(n7467), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6320));
   INVX1 U2259 (.Y(n7467), 
	.A(\ram[219][11] ));
   OAI22X1 U2260 (.Y(n4096), 
	.B1(n7468), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6322));
   INVX1 U2261 (.Y(n7468), 
	.A(\ram[219][10] ));
   OAI22X1 U2262 (.Y(n4095), 
	.B1(n7469), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6324));
   INVX1 U2263 (.Y(n7469), 
	.A(\ram[219][9] ));
   OAI22X1 U2264 (.Y(n4094), 
	.B1(n7470), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6326));
   INVX1 U2265 (.Y(n7470), 
	.A(\ram[219][8] ));
   OAI22X1 U2266 (.Y(n4093), 
	.B1(n7471), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6328));
   INVX1 U2267 (.Y(n7471), 
	.A(\ram[219][7] ));
   OAI22X1 U2268 (.Y(n4092), 
	.B1(n7472), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6330));
   INVX1 U2269 (.Y(n7472), 
	.A(\ram[219][6] ));
   OAI22X1 U2270 (.Y(n4091), 
	.B1(n7473), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6332));
   INVX1 U2271 (.Y(n7473), 
	.A(\ram[219][5] ));
   OAI22X1 U2272 (.Y(n4090), 
	.B1(n7474), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6334));
   INVX1 U2273 (.Y(n7474), 
	.A(\ram[219][4] ));
   OAI22X1 U2274 (.Y(n4089), 
	.B1(n7475), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6336));
   INVX1 U2275 (.Y(n7475), 
	.A(\ram[219][3] ));
   OAI22X1 U2276 (.Y(n4088), 
	.B1(n7476), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6338));
   INVX1 U2277 (.Y(n7476), 
	.A(\ram[219][2] ));
   OAI22X1 U2278 (.Y(n4087), 
	.B1(n7477), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6306));
   INVX1 U2279 (.Y(n7477), 
	.A(\ram[219][1] ));
   OAI22X1 U2280 (.Y(n4086), 
	.B1(n7478), 
	.B0(n7462), 
	.A1(n7461), 
	.A0(n6309));
   INVX1 U2281 (.Y(n7478), 
	.A(\ram[219][0] ));
   NOR2BX1 U2282 (.Y(n7462), 
	.B(n7461), 
	.AN(mem_write_en));
   NAND2X1 U2283 (.Y(n7461), 
	.B(n6610), 
	.A(n7406));
   OAI22X1 U2284 (.Y(n4085), 
	.B1(n7481), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6311));
   INVX1 U2285 (.Y(n7481), 
	.A(\ram[218][15] ));
   OAI22X1 U2286 (.Y(n4084), 
	.B1(n7482), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6314));
   INVX1 U2287 (.Y(n7482), 
	.A(\ram[218][14] ));
   OAI22X1 U2288 (.Y(n4083), 
	.B1(n7483), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6316));
   INVX1 U2289 (.Y(n7483), 
	.A(\ram[218][13] ));
   OAI22X1 U2290 (.Y(n4082), 
	.B1(n7484), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6318));
   INVX1 U2291 (.Y(n7484), 
	.A(\ram[218][12] ));
   OAI22X1 U2292 (.Y(n4081), 
	.B1(n7485), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6320));
   INVX1 U2293 (.Y(n7485), 
	.A(\ram[218][11] ));
   OAI22X1 U2294 (.Y(n4080), 
	.B1(n7486), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6322));
   INVX1 U2295 (.Y(n7486), 
	.A(\ram[218][10] ));
   OAI22X1 U2296 (.Y(n4079), 
	.B1(n7487), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6324));
   INVX1 U2297 (.Y(n7487), 
	.A(\ram[218][9] ));
   OAI22X1 U2298 (.Y(n4078), 
	.B1(n7488), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6326));
   INVX1 U2299 (.Y(n7488), 
	.A(\ram[218][8] ));
   OAI22X1 U2300 (.Y(n4077), 
	.B1(n7489), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6328));
   INVX1 U2301 (.Y(n7489), 
	.A(\ram[218][7] ));
   OAI22X1 U2302 (.Y(n4076), 
	.B1(n7490), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6330));
   INVX1 U2303 (.Y(n7490), 
	.A(\ram[218][6] ));
   OAI22X1 U2304 (.Y(n4075), 
	.B1(n7491), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6332));
   INVX1 U2305 (.Y(n7491), 
	.A(\ram[218][5] ));
   OAI22X1 U2306 (.Y(n4074), 
	.B1(n7492), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6334));
   INVX1 U2307 (.Y(n7492), 
	.A(\ram[218][4] ));
   OAI22X1 U2308 (.Y(n4073), 
	.B1(n7493), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6336));
   INVX1 U2309 (.Y(n7493), 
	.A(\ram[218][3] ));
   OAI22X1 U2310 (.Y(n4072), 
	.B1(n7494), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6338));
   INVX1 U2311 (.Y(n7494), 
	.A(\ram[218][2] ));
   OAI22X1 U2312 (.Y(n4071), 
	.B1(n7495), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6306));
   INVX1 U2313 (.Y(n7495), 
	.A(\ram[218][1] ));
   OAI22X1 U2314 (.Y(n4070), 
	.B1(n7496), 
	.B0(n7480), 
	.A1(n7479), 
	.A0(n6309));
   INVX1 U2315 (.Y(n7496), 
	.A(\ram[218][0] ));
   NOR2BX1 U2316 (.Y(n7480), 
	.B(n7479), 
	.AN(mem_write_en));
   NAND2X1 U2317 (.Y(n7479), 
	.B(n6629), 
	.A(n7406));
   OAI22X1 U2318 (.Y(n4069), 
	.B1(n7499), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6311));
   INVX1 U2319 (.Y(n7499), 
	.A(\ram[217][15] ));
   OAI22X1 U2320 (.Y(n4068), 
	.B1(n7500), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6314));
   INVX1 U2321 (.Y(n7500), 
	.A(\ram[217][14] ));
   OAI22X1 U2322 (.Y(n4067), 
	.B1(n7501), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6316));
   INVX1 U2323 (.Y(n7501), 
	.A(\ram[217][13] ));
   OAI22X1 U2324 (.Y(n4066), 
	.B1(n7502), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6318));
   INVX1 U2325 (.Y(n7502), 
	.A(\ram[217][12] ));
   OAI22X1 U2326 (.Y(n4065), 
	.B1(n7503), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6320));
   INVX1 U2327 (.Y(n7503), 
	.A(\ram[217][11] ));
   OAI22X1 U2328 (.Y(n4064), 
	.B1(n7504), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6322));
   INVX1 U2329 (.Y(n7504), 
	.A(\ram[217][10] ));
   OAI22X1 U2330 (.Y(n4063), 
	.B1(n7505), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6324));
   INVX1 U2331 (.Y(n7505), 
	.A(\ram[217][9] ));
   OAI22X1 U2332 (.Y(n4062), 
	.B1(n7506), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6326));
   INVX1 U2333 (.Y(n7506), 
	.A(\ram[217][8] ));
   OAI22X1 U2334 (.Y(n4061), 
	.B1(n7507), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6328));
   INVX1 U2335 (.Y(n7507), 
	.A(\ram[217][7] ));
   OAI22X1 U2336 (.Y(n4060), 
	.B1(n7508), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6330));
   INVX1 U2337 (.Y(n7508), 
	.A(\ram[217][6] ));
   OAI22X1 U2338 (.Y(n4059), 
	.B1(n7509), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6332));
   INVX1 U2339 (.Y(n7509), 
	.A(\ram[217][5] ));
   OAI22X1 U2340 (.Y(n4058), 
	.B1(n7510), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6334));
   INVX1 U2341 (.Y(n7510), 
	.A(\ram[217][4] ));
   OAI22X1 U2342 (.Y(n4057), 
	.B1(n7511), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6336));
   INVX1 U2343 (.Y(n7511), 
	.A(\ram[217][3] ));
   OAI22X1 U2344 (.Y(n4056), 
	.B1(n7512), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6338));
   INVX1 U2345 (.Y(n7512), 
	.A(\ram[217][2] ));
   OAI22X1 U2346 (.Y(n4055), 
	.B1(n7513), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6306));
   INVX1 U2347 (.Y(n7513), 
	.A(\ram[217][1] ));
   OAI22X1 U2348 (.Y(n4054), 
	.B1(n7514), 
	.B0(n7498), 
	.A1(n7497), 
	.A0(n6309));
   INVX1 U2349 (.Y(n7514), 
	.A(\ram[217][0] ));
   NOR2BX1 U2350 (.Y(n7498), 
	.B(n7497), 
	.AN(mem_write_en));
   NAND2X1 U2351 (.Y(n7497), 
	.B(n6342), 
	.A(n7406));
   OAI22X1 U2352 (.Y(n4053), 
	.B1(n7517), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6311));
   INVX1 U2353 (.Y(n7517), 
	.A(\ram[216][15] ));
   OAI22X1 U2354 (.Y(n4052), 
	.B1(n7518), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6314));
   INVX1 U2355 (.Y(n7518), 
	.A(\ram[216][14] ));
   OAI22X1 U2356 (.Y(n4051), 
	.B1(n7519), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6316));
   INVX1 U2357 (.Y(n7519), 
	.A(\ram[216][13] ));
   OAI22X1 U2358 (.Y(n4050), 
	.B1(n7520), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6318));
   INVX1 U2359 (.Y(n7520), 
	.A(\ram[216][12] ));
   OAI22X1 U2360 (.Y(n4049), 
	.B1(n7521), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6320));
   INVX1 U2361 (.Y(n7521), 
	.A(\ram[216][11] ));
   OAI22X1 U2362 (.Y(n4048), 
	.B1(n7522), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6322));
   INVX1 U2363 (.Y(n7522), 
	.A(\ram[216][10] ));
   OAI22X1 U2364 (.Y(n4047), 
	.B1(n7523), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6324));
   INVX1 U2365 (.Y(n7523), 
	.A(\ram[216][9] ));
   OAI22X1 U2366 (.Y(n4046), 
	.B1(n7524), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6326));
   INVX1 U2367 (.Y(n7524), 
	.A(\ram[216][8] ));
   OAI22X1 U2368 (.Y(n4045), 
	.B1(n7525), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6328));
   INVX1 U2369 (.Y(n7525), 
	.A(\ram[216][7] ));
   OAI22X1 U2370 (.Y(n4044), 
	.B1(n7526), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6330));
   INVX1 U2371 (.Y(n7526), 
	.A(\ram[216][6] ));
   OAI22X1 U2372 (.Y(n4043), 
	.B1(n7527), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6332));
   INVX1 U2373 (.Y(n7527), 
	.A(\ram[216][5] ));
   OAI22X1 U2374 (.Y(n4042), 
	.B1(n7528), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6334));
   INVX1 U2375 (.Y(n7528), 
	.A(\ram[216][4] ));
   OAI22X1 U2376 (.Y(n4041), 
	.B1(n7529), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6336));
   INVX1 U2377 (.Y(n7529), 
	.A(\ram[216][3] ));
   OAI22X1 U2378 (.Y(n4040), 
	.B1(n7530), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6338));
   INVX1 U2379 (.Y(n7530), 
	.A(\ram[216][2] ));
   OAI22X1 U2380 (.Y(n4039), 
	.B1(n7531), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6306));
   INVX1 U2381 (.Y(n7531), 
	.A(\ram[216][1] ));
   OAI22X1 U2382 (.Y(n4038), 
	.B1(n7532), 
	.B0(n7516), 
	.A1(n7515), 
	.A0(n6309));
   INVX1 U2383 (.Y(n7532), 
	.A(\ram[216][0] ));
   NOR2BX1 U2384 (.Y(n7516), 
	.B(n7515), 
	.AN(mem_write_en));
   NAND2X1 U2385 (.Y(n7515), 
	.B(n6362), 
	.A(n7406));
   OAI22X1 U2386 (.Y(n4037), 
	.B1(n7535), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6311));
   INVX1 U2387 (.Y(n7535), 
	.A(\ram[215][15] ));
   OAI22X1 U2388 (.Y(n4036), 
	.B1(n7536), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6314));
   INVX1 U2389 (.Y(n7536), 
	.A(\ram[215][14] ));
   OAI22X1 U2390 (.Y(n4035), 
	.B1(n7537), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6316));
   INVX1 U2391 (.Y(n7537), 
	.A(\ram[215][13] ));
   OAI22X1 U2392 (.Y(n4034), 
	.B1(n7538), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6318));
   INVX1 U2393 (.Y(n7538), 
	.A(\ram[215][12] ));
   OAI22X1 U2394 (.Y(n4033), 
	.B1(n7539), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6320));
   INVX1 U2395 (.Y(n7539), 
	.A(\ram[215][11] ));
   OAI22X1 U2396 (.Y(n4032), 
	.B1(n7540), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6322));
   INVX1 U2397 (.Y(n7540), 
	.A(\ram[215][10] ));
   OAI22X1 U2398 (.Y(n4031), 
	.B1(n7541), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6324));
   INVX1 U2399 (.Y(n7541), 
	.A(\ram[215][9] ));
   OAI22X1 U2400 (.Y(n4030), 
	.B1(n7542), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6326));
   INVX1 U2401 (.Y(n7542), 
	.A(\ram[215][8] ));
   OAI22X1 U2402 (.Y(n4029), 
	.B1(n7543), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6328));
   INVX1 U2403 (.Y(n7543), 
	.A(\ram[215][7] ));
   OAI22X1 U2404 (.Y(n4028), 
	.B1(n7544), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6330));
   INVX1 U2405 (.Y(n7544), 
	.A(\ram[215][6] ));
   OAI22X1 U2406 (.Y(n4027), 
	.B1(n7545), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6332));
   INVX1 U2407 (.Y(n7545), 
	.A(\ram[215][5] ));
   OAI22X1 U2408 (.Y(n4026), 
	.B1(n7546), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6334));
   INVX1 U2409 (.Y(n7546), 
	.A(\ram[215][4] ));
   OAI22X1 U2410 (.Y(n4025), 
	.B1(n7547), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6336));
   INVX1 U2411 (.Y(n7547), 
	.A(\ram[215][3] ));
   OAI22X1 U2412 (.Y(n4024), 
	.B1(n7548), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6338));
   INVX1 U2413 (.Y(n7548), 
	.A(\ram[215][2] ));
   OAI22X1 U2414 (.Y(n4023), 
	.B1(n7549), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6306));
   INVX1 U2415 (.Y(n7549), 
	.A(\ram[215][1] ));
   OAI22X1 U2416 (.Y(n4022), 
	.B1(n7550), 
	.B0(n7534), 
	.A1(n7533), 
	.A0(n6309));
   INVX1 U2417 (.Y(n7550), 
	.A(\ram[215][0] ));
   NOR2BX1 U2418 (.Y(n7534), 
	.B(n7533), 
	.AN(mem_write_en));
   NAND2X1 U2419 (.Y(n7533), 
	.B(n6381), 
	.A(n7406));
   OAI22X1 U2420 (.Y(n4021), 
	.B1(n7553), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6311));
   INVX1 U2421 (.Y(n7553), 
	.A(\ram[214][15] ));
   OAI22X1 U2422 (.Y(n4020), 
	.B1(n7554), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6314));
   INVX1 U2423 (.Y(n7554), 
	.A(\ram[214][14] ));
   OAI22X1 U2424 (.Y(n4019), 
	.B1(n7555), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6316));
   INVX1 U2425 (.Y(n7555), 
	.A(\ram[214][13] ));
   OAI22X1 U2426 (.Y(n4018), 
	.B1(n7556), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6318));
   INVX1 U2427 (.Y(n7556), 
	.A(\ram[214][12] ));
   OAI22X1 U2428 (.Y(n4017), 
	.B1(n7557), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6320));
   INVX1 U2429 (.Y(n7557), 
	.A(\ram[214][11] ));
   OAI22X1 U2430 (.Y(n4016), 
	.B1(n7558), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6322));
   INVX1 U2431 (.Y(n7558), 
	.A(\ram[214][10] ));
   OAI22X1 U2432 (.Y(n4015), 
	.B1(n7559), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6324));
   INVX1 U2433 (.Y(n7559), 
	.A(\ram[214][9] ));
   OAI22X1 U2434 (.Y(n4014), 
	.B1(n7560), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6326));
   INVX1 U2435 (.Y(n7560), 
	.A(\ram[214][8] ));
   OAI22X1 U2436 (.Y(n4013), 
	.B1(n7561), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6328));
   INVX1 U2437 (.Y(n7561), 
	.A(\ram[214][7] ));
   OAI22X1 U2438 (.Y(n4012), 
	.B1(n7562), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6330));
   INVX1 U2439 (.Y(n7562), 
	.A(\ram[214][6] ));
   OAI22X1 U2440 (.Y(n4011), 
	.B1(n7563), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6332));
   INVX1 U2441 (.Y(n7563), 
	.A(\ram[214][5] ));
   OAI22X1 U2442 (.Y(n4010), 
	.B1(n7564), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6334));
   INVX1 U2443 (.Y(n7564), 
	.A(\ram[214][4] ));
   OAI22X1 U2444 (.Y(n4009), 
	.B1(n7565), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6336));
   INVX1 U2445 (.Y(n7565), 
	.A(\ram[214][3] ));
   OAI22X1 U2446 (.Y(n4008), 
	.B1(n7566), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6338));
   INVX1 U2447 (.Y(n7566), 
	.A(\ram[214][2] ));
   OAI22X1 U2448 (.Y(n4007), 
	.B1(n7567), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6306));
   INVX1 U2449 (.Y(n7567), 
	.A(\ram[214][1] ));
   OAI22X1 U2450 (.Y(n4006), 
	.B1(n7568), 
	.B0(n7552), 
	.A1(n7551), 
	.A0(n6309));
   INVX1 U2451 (.Y(n7568), 
	.A(\ram[214][0] ));
   NOR2BX1 U2452 (.Y(n7552), 
	.B(n7551), 
	.AN(mem_write_en));
   NAND2X1 U2453 (.Y(n7551), 
	.B(n6400), 
	.A(n7406));
   OAI22X1 U2454 (.Y(n4005), 
	.B1(n7571), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6311));
   INVX1 U2455 (.Y(n7571), 
	.A(\ram[213][15] ));
   OAI22X1 U2456 (.Y(n4004), 
	.B1(n7572), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6314));
   INVX1 U2457 (.Y(n7572), 
	.A(\ram[213][14] ));
   OAI22X1 U2458 (.Y(n4003), 
	.B1(n7573), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6316));
   INVX1 U2459 (.Y(n7573), 
	.A(\ram[213][13] ));
   OAI22X1 U2460 (.Y(n4002), 
	.B1(n7574), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6318));
   INVX1 U2461 (.Y(n7574), 
	.A(\ram[213][12] ));
   OAI22X1 U2462 (.Y(n4001), 
	.B1(n7575), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6320));
   INVX1 U2463 (.Y(n7575), 
	.A(\ram[213][11] ));
   OAI22X1 U2464 (.Y(n4000), 
	.B1(n7576), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6322));
   INVX1 U2465 (.Y(n7576), 
	.A(\ram[213][10] ));
   OAI22X1 U2466 (.Y(n3999), 
	.B1(n7577), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6324));
   INVX1 U2467 (.Y(n7577), 
	.A(\ram[213][9] ));
   OAI22X1 U2468 (.Y(n3998), 
	.B1(n7578), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6326));
   INVX1 U2469 (.Y(n7578), 
	.A(\ram[213][8] ));
   OAI22X1 U2470 (.Y(n3997), 
	.B1(n7579), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6328));
   INVX1 U2471 (.Y(n7579), 
	.A(\ram[213][7] ));
   OAI22X1 U2472 (.Y(n3996), 
	.B1(n7580), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6330));
   INVX1 U2473 (.Y(n7580), 
	.A(\ram[213][6] ));
   OAI22X1 U2474 (.Y(n3995), 
	.B1(n7581), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6332));
   INVX1 U2475 (.Y(n7581), 
	.A(\ram[213][5] ));
   OAI22X1 U2476 (.Y(n3994), 
	.B1(n7582), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6334));
   INVX1 U2477 (.Y(n7582), 
	.A(\ram[213][4] ));
   OAI22X1 U2478 (.Y(n3993), 
	.B1(n7583), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6336));
   INVX1 U2479 (.Y(n7583), 
	.A(\ram[213][3] ));
   OAI22X1 U2480 (.Y(n3992), 
	.B1(n7584), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6338));
   INVX1 U2481 (.Y(n7584), 
	.A(\ram[213][2] ));
   OAI22X1 U2482 (.Y(n3991), 
	.B1(n7585), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6306));
   INVX1 U2483 (.Y(n7585), 
	.A(\ram[213][1] ));
   OAI22X1 U2484 (.Y(n3990), 
	.B1(n7586), 
	.B0(n7570), 
	.A1(n7569), 
	.A0(n6309));
   INVX1 U2485 (.Y(n7586), 
	.A(\ram[213][0] ));
   NOR2BX1 U2486 (.Y(n7570), 
	.B(n7569), 
	.AN(mem_write_en));
   NAND2X1 U2487 (.Y(n7569), 
	.B(n6419), 
	.A(n7406));
   OAI22X1 U2488 (.Y(n3989), 
	.B1(n7589), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6311));
   INVX1 U2489 (.Y(n7589), 
	.A(\ram[212][15] ));
   OAI22X1 U2490 (.Y(n3988), 
	.B1(n7590), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6314));
   INVX1 U2491 (.Y(n7590), 
	.A(\ram[212][14] ));
   OAI22X1 U2492 (.Y(n3987), 
	.B1(n7591), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6316));
   INVX1 U2493 (.Y(n7591), 
	.A(\ram[212][13] ));
   OAI22X1 U2494 (.Y(n3986), 
	.B1(n7592), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6318));
   INVX1 U2495 (.Y(n7592), 
	.A(\ram[212][12] ));
   OAI22X1 U2496 (.Y(n3985), 
	.B1(n7593), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6320));
   INVX1 U2497 (.Y(n7593), 
	.A(\ram[212][11] ));
   OAI22X1 U2498 (.Y(n3984), 
	.B1(n7594), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6322));
   INVX1 U2499 (.Y(n7594), 
	.A(\ram[212][10] ));
   OAI22X1 U2500 (.Y(n3983), 
	.B1(n7595), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6324));
   INVX1 U2501 (.Y(n7595), 
	.A(\ram[212][9] ));
   OAI22X1 U2502 (.Y(n3982), 
	.B1(n7596), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6326));
   INVX1 U2503 (.Y(n7596), 
	.A(\ram[212][8] ));
   OAI22X1 U2504 (.Y(n3981), 
	.B1(n7597), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6328));
   INVX1 U2505 (.Y(n7597), 
	.A(\ram[212][7] ));
   OAI22X1 U2506 (.Y(n3980), 
	.B1(n7598), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6330));
   INVX1 U2507 (.Y(n7598), 
	.A(\ram[212][6] ));
   OAI22X1 U2508 (.Y(n3979), 
	.B1(n7599), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6332));
   INVX1 U2509 (.Y(n7599), 
	.A(\ram[212][5] ));
   OAI22X1 U2510 (.Y(n3978), 
	.B1(n7600), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6334));
   INVX1 U2511 (.Y(n7600), 
	.A(\ram[212][4] ));
   OAI22X1 U2512 (.Y(n3977), 
	.B1(n7601), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6336));
   INVX1 U2513 (.Y(n7601), 
	.A(\ram[212][3] ));
   OAI22X1 U2514 (.Y(n3976), 
	.B1(n7602), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6338));
   INVX1 U2515 (.Y(n7602), 
	.A(\ram[212][2] ));
   OAI22X1 U2516 (.Y(n3975), 
	.B1(n7603), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6306));
   INVX1 U2517 (.Y(n7603), 
	.A(\ram[212][1] ));
   OAI22X1 U2518 (.Y(n3974), 
	.B1(n7604), 
	.B0(n7588), 
	.A1(n7587), 
	.A0(n6309));
   INVX1 U2519 (.Y(n7604), 
	.A(\ram[212][0] ));
   NOR2BX1 U2520 (.Y(n7588), 
	.B(n7587), 
	.AN(mem_write_en));
   NAND2X1 U2521 (.Y(n7587), 
	.B(n6438), 
	.A(n7406));
   OAI22X1 U2522 (.Y(n3973), 
	.B1(n7607), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6311));
   INVX1 U2523 (.Y(n7607), 
	.A(\ram[211][15] ));
   OAI22X1 U2524 (.Y(n3972), 
	.B1(n7608), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6314));
   INVX1 U2525 (.Y(n7608), 
	.A(\ram[211][14] ));
   OAI22X1 U2526 (.Y(n3971), 
	.B1(n7609), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6316));
   INVX1 U2527 (.Y(n7609), 
	.A(\ram[211][13] ));
   OAI22X1 U2528 (.Y(n3970), 
	.B1(n7610), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6318));
   INVX1 U2529 (.Y(n7610), 
	.A(\ram[211][12] ));
   OAI22X1 U2530 (.Y(n3969), 
	.B1(n7611), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6320));
   INVX1 U2531 (.Y(n7611), 
	.A(\ram[211][11] ));
   OAI22X1 U2532 (.Y(n3968), 
	.B1(n7612), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6322));
   INVX1 U2533 (.Y(n7612), 
	.A(\ram[211][10] ));
   OAI22X1 U2534 (.Y(n3967), 
	.B1(n7613), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6324));
   INVX1 U2535 (.Y(n7613), 
	.A(\ram[211][9] ));
   OAI22X1 U2536 (.Y(n3966), 
	.B1(n7614), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6326));
   INVX1 U2537 (.Y(n7614), 
	.A(\ram[211][8] ));
   OAI22X1 U2538 (.Y(n3965), 
	.B1(n7615), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6328));
   INVX1 U2539 (.Y(n7615), 
	.A(\ram[211][7] ));
   OAI22X1 U2540 (.Y(n3964), 
	.B1(n7616), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6330));
   INVX1 U2541 (.Y(n7616), 
	.A(\ram[211][6] ));
   OAI22X1 U2542 (.Y(n3963), 
	.B1(n7617), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6332));
   INVX1 U2543 (.Y(n7617), 
	.A(\ram[211][5] ));
   OAI22X1 U2544 (.Y(n3962), 
	.B1(n7618), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6334));
   INVX1 U2545 (.Y(n7618), 
	.A(\ram[211][4] ));
   OAI22X1 U2546 (.Y(n3961), 
	.B1(n7619), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6336));
   INVX1 U2547 (.Y(n7619), 
	.A(\ram[211][3] ));
   OAI22X1 U2548 (.Y(n3960), 
	.B1(n7620), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6338));
   INVX1 U2549 (.Y(n7620), 
	.A(\ram[211][2] ));
   OAI22X1 U2550 (.Y(n3959), 
	.B1(n7621), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6306));
   INVX1 U2551 (.Y(n7621), 
	.A(\ram[211][1] ));
   OAI22X1 U2552 (.Y(n3958), 
	.B1(n7622), 
	.B0(n7606), 
	.A1(n7605), 
	.A0(n6309));
   INVX1 U2553 (.Y(n7622), 
	.A(\ram[211][0] ));
   NOR2BX1 U2554 (.Y(n7606), 
	.B(n7605), 
	.AN(mem_write_en));
   NAND2X1 U2555 (.Y(n7605), 
	.B(n6457), 
	.A(n7406));
   OAI22X1 U2556 (.Y(n3957), 
	.B1(n7625), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6311));
   INVX1 U2557 (.Y(n7625), 
	.A(\ram[210][15] ));
   OAI22X1 U2558 (.Y(n3956), 
	.B1(n7626), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6314));
   INVX1 U2559 (.Y(n7626), 
	.A(\ram[210][14] ));
   OAI22X1 U2560 (.Y(n3955), 
	.B1(n7627), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6316));
   INVX1 U2561 (.Y(n7627), 
	.A(\ram[210][13] ));
   OAI22X1 U2562 (.Y(n3954), 
	.B1(n7628), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6318));
   INVX1 U2563 (.Y(n7628), 
	.A(\ram[210][12] ));
   OAI22X1 U2564 (.Y(n3953), 
	.B1(n7629), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6320));
   INVX1 U2565 (.Y(n7629), 
	.A(\ram[210][11] ));
   OAI22X1 U2566 (.Y(n3952), 
	.B1(n7630), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6322));
   INVX1 U2567 (.Y(n7630), 
	.A(\ram[210][10] ));
   OAI22X1 U2568 (.Y(n3951), 
	.B1(n7631), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6324));
   INVX1 U2569 (.Y(n7631), 
	.A(\ram[210][9] ));
   OAI22X1 U2570 (.Y(n3950), 
	.B1(n7632), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6326));
   INVX1 U2571 (.Y(n7632), 
	.A(\ram[210][8] ));
   OAI22X1 U2572 (.Y(n3949), 
	.B1(n7633), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6328));
   INVX1 U2573 (.Y(n7633), 
	.A(\ram[210][7] ));
   OAI22X1 U2574 (.Y(n3948), 
	.B1(n7634), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6330));
   INVX1 U2575 (.Y(n7634), 
	.A(\ram[210][6] ));
   OAI22X1 U2576 (.Y(n3947), 
	.B1(n7635), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6332));
   INVX1 U2577 (.Y(n7635), 
	.A(\ram[210][5] ));
   OAI22X1 U2578 (.Y(n3946), 
	.B1(n7636), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6334));
   INVX1 U2579 (.Y(n7636), 
	.A(\ram[210][4] ));
   OAI22X1 U2580 (.Y(n3945), 
	.B1(n7637), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6336));
   INVX1 U2581 (.Y(n7637), 
	.A(\ram[210][3] ));
   OAI22X1 U2582 (.Y(n3944), 
	.B1(n7638), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6338));
   INVX1 U2583 (.Y(n7638), 
	.A(\ram[210][2] ));
   OAI22X1 U2584 (.Y(n3943), 
	.B1(n7639), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6306));
   INVX1 U2585 (.Y(n7639), 
	.A(\ram[210][1] ));
   OAI22X1 U2586 (.Y(n3942), 
	.B1(n7640), 
	.B0(n7624), 
	.A1(n7623), 
	.A0(n6309));
   INVX1 U2587 (.Y(n7640), 
	.A(\ram[210][0] ));
   NOR2BX1 U2588 (.Y(n7624), 
	.B(n7623), 
	.AN(mem_write_en));
   NAND2X1 U2589 (.Y(n7623), 
	.B(n6476), 
	.A(n7406));
   OAI22X1 U2590 (.Y(n3941), 
	.B1(n7643), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6311));
   INVX1 U2591 (.Y(n7643), 
	.A(\ram[209][15] ));
   OAI22X1 U2592 (.Y(n3940), 
	.B1(n7644), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6314));
   INVX1 U2593 (.Y(n7644), 
	.A(\ram[209][14] ));
   OAI22X1 U2594 (.Y(n3939), 
	.B1(n7645), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6316));
   INVX1 U2595 (.Y(n7645), 
	.A(\ram[209][13] ));
   OAI22X1 U2596 (.Y(n3938), 
	.B1(n7646), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6318));
   INVX1 U2597 (.Y(n7646), 
	.A(\ram[209][12] ));
   OAI22X1 U2598 (.Y(n3937), 
	.B1(n7647), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6320));
   INVX1 U2599 (.Y(n7647), 
	.A(\ram[209][11] ));
   OAI22X1 U2600 (.Y(n3936), 
	.B1(n7648), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6322));
   INVX1 U2601 (.Y(n7648), 
	.A(\ram[209][10] ));
   OAI22X1 U2602 (.Y(n3935), 
	.B1(n7649), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6324));
   INVX1 U2603 (.Y(n7649), 
	.A(\ram[209][9] ));
   OAI22X1 U2604 (.Y(n3934), 
	.B1(n7650), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6326));
   INVX1 U2605 (.Y(n7650), 
	.A(\ram[209][8] ));
   OAI22X1 U2606 (.Y(n3933), 
	.B1(n7651), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6328));
   INVX1 U2607 (.Y(n7651), 
	.A(\ram[209][7] ));
   OAI22X1 U2608 (.Y(n3932), 
	.B1(n7652), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6330));
   INVX1 U2609 (.Y(n7652), 
	.A(\ram[209][6] ));
   OAI22X1 U2610 (.Y(n3931), 
	.B1(n7653), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6332));
   INVX1 U2611 (.Y(n7653), 
	.A(\ram[209][5] ));
   OAI22X1 U2612 (.Y(n3930), 
	.B1(n7654), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6334));
   INVX1 U2613 (.Y(n7654), 
	.A(\ram[209][4] ));
   OAI22X1 U2614 (.Y(n3929), 
	.B1(n7655), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6336));
   INVX1 U2615 (.Y(n7655), 
	.A(\ram[209][3] ));
   OAI22X1 U2616 (.Y(n3928), 
	.B1(n7656), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6338));
   INVX1 U2617 (.Y(n7656), 
	.A(\ram[209][2] ));
   OAI22X1 U2618 (.Y(n3927), 
	.B1(n7657), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6306));
   INVX1 U2619 (.Y(n7657), 
	.A(\ram[209][1] ));
   OAI22X1 U2620 (.Y(n3926), 
	.B1(n7658), 
	.B0(n7642), 
	.A1(n7641), 
	.A0(n6309));
   INVX1 U2621 (.Y(n7658), 
	.A(\ram[209][0] ));
   NOR2BX1 U2622 (.Y(n7642), 
	.B(n7641), 
	.AN(mem_write_en));
   NAND2X1 U2623 (.Y(n7641), 
	.B(n6495), 
	.A(n7406));
   OAI22X1 U2624 (.Y(n3925), 
	.B1(n7661), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6311));
   INVX1 U2625 (.Y(n7661), 
	.A(\ram[208][15] ));
   OAI22X1 U2626 (.Y(n3924), 
	.B1(n7662), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6314));
   INVX1 U2627 (.Y(n7662), 
	.A(\ram[208][14] ));
   OAI22X1 U2628 (.Y(n3923), 
	.B1(n7663), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6316));
   INVX1 U2629 (.Y(n7663), 
	.A(\ram[208][13] ));
   OAI22X1 U2630 (.Y(n3922), 
	.B1(n7664), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6318));
   INVX1 U2631 (.Y(n7664), 
	.A(\ram[208][12] ));
   OAI22X1 U2632 (.Y(n3921), 
	.B1(n7665), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6320));
   INVX1 U2633 (.Y(n7665), 
	.A(\ram[208][11] ));
   OAI22X1 U2634 (.Y(n3920), 
	.B1(n7666), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6322));
   INVX1 U2635 (.Y(n7666), 
	.A(\ram[208][10] ));
   OAI22X1 U2636 (.Y(n3919), 
	.B1(n7667), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6324));
   INVX1 U2637 (.Y(n7667), 
	.A(\ram[208][9] ));
   OAI22X1 U2638 (.Y(n3918), 
	.B1(n7668), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6326));
   INVX1 U2639 (.Y(n7668), 
	.A(\ram[208][8] ));
   OAI22X1 U2640 (.Y(n3917), 
	.B1(n7669), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6328));
   INVX1 U2641 (.Y(n7669), 
	.A(\ram[208][7] ));
   OAI22X1 U2642 (.Y(n3916), 
	.B1(n7670), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6330));
   INVX1 U2643 (.Y(n7670), 
	.A(\ram[208][6] ));
   OAI22X1 U2644 (.Y(n3915), 
	.B1(n7671), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6332));
   INVX1 U2645 (.Y(n7671), 
	.A(\ram[208][5] ));
   OAI22X1 U2646 (.Y(n3914), 
	.B1(n7672), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6334));
   INVX1 U2647 (.Y(n7672), 
	.A(\ram[208][4] ));
   OAI22X1 U2648 (.Y(n3913), 
	.B1(n7673), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6336));
   INVX1 U2649 (.Y(n7673), 
	.A(\ram[208][3] ));
   OAI22X1 U2650 (.Y(n3912), 
	.B1(n7674), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6338));
   INVX1 U2651 (.Y(n7674), 
	.A(\ram[208][2] ));
   OAI22X1 U2652 (.Y(n3911), 
	.B1(n7675), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6306));
   INVX1 U2653 (.Y(n7675), 
	.A(\ram[208][1] ));
   OAI22X1 U2654 (.Y(n3910), 
	.B1(n7676), 
	.B0(n7660), 
	.A1(n7659), 
	.A0(n6309));
   INVX1 U2655 (.Y(n7676), 
	.A(\ram[208][0] ));
   NOR2BX1 U2656 (.Y(n7660), 
	.B(n7659), 
	.AN(mem_write_en));
   NAND2X1 U2657 (.Y(n7659), 
	.B(n6514), 
	.A(n7406));
   OAI22X1 U2658 (.Y(n3909), 
	.B1(n7679), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6311));
   INVX1 U2659 (.Y(n7679), 
	.A(\ram[207][15] ));
   OAI22X1 U2660 (.Y(n3908), 
	.B1(n7680), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6314));
   INVX1 U2661 (.Y(n7680), 
	.A(\ram[207][14] ));
   OAI22X1 U2662 (.Y(n3907), 
	.B1(n7681), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6316));
   INVX1 U2663 (.Y(n7681), 
	.A(\ram[207][13] ));
   OAI22X1 U2664 (.Y(n3906), 
	.B1(n7682), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6318));
   INVX1 U2665 (.Y(n7682), 
	.A(\ram[207][12] ));
   OAI22X1 U2666 (.Y(n3905), 
	.B1(n7683), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6320));
   INVX1 U2667 (.Y(n7683), 
	.A(\ram[207][11] ));
   OAI22X1 U2668 (.Y(n3904), 
	.B1(n7684), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6322));
   INVX1 U2669 (.Y(n7684), 
	.A(\ram[207][10] ));
   OAI22X1 U2670 (.Y(n3903), 
	.B1(n7685), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6324));
   INVX1 U2671 (.Y(n7685), 
	.A(\ram[207][9] ));
   OAI22X1 U2672 (.Y(n3902), 
	.B1(n7686), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6326));
   INVX1 U2673 (.Y(n7686), 
	.A(\ram[207][8] ));
   OAI22X1 U2674 (.Y(n3901), 
	.B1(n7687), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6328));
   INVX1 U2675 (.Y(n7687), 
	.A(\ram[207][7] ));
   OAI22X1 U2676 (.Y(n3900), 
	.B1(n7688), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6330));
   INVX1 U2677 (.Y(n7688), 
	.A(\ram[207][6] ));
   OAI22X1 U2678 (.Y(n3899), 
	.B1(n7689), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6332));
   INVX1 U2679 (.Y(n7689), 
	.A(\ram[207][5] ));
   OAI22X1 U2680 (.Y(n3898), 
	.B1(n7690), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6334));
   INVX1 U2681 (.Y(n7690), 
	.A(\ram[207][4] ));
   OAI22X1 U2682 (.Y(n3897), 
	.B1(n7691), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6336));
   INVX1 U2683 (.Y(n7691), 
	.A(\ram[207][3] ));
   OAI22X1 U2684 (.Y(n3896), 
	.B1(n7692), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6338));
   INVX1 U2685 (.Y(n7692), 
	.A(\ram[207][2] ));
   OAI22X1 U2686 (.Y(n3895), 
	.B1(n7693), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6306));
   INVX1 U2687 (.Y(n7693), 
	.A(\ram[207][1] ));
   OAI22X1 U2688 (.Y(n3894), 
	.B1(n7694), 
	.B0(n7678), 
	.A1(n7677), 
	.A0(n6309));
   INVX1 U2689 (.Y(n7694), 
	.A(\ram[207][0] ));
   NOR2BX1 U2690 (.Y(n7678), 
	.B(n7677), 
	.AN(mem_write_en));
   NAND2X1 U2691 (.Y(n7677), 
	.B(n6533), 
	.A(n7695));
   OAI22X1 U2692 (.Y(n3893), 
	.B1(n7698), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6311));
   INVX1 U2693 (.Y(n7698), 
	.A(\ram[206][15] ));
   OAI22X1 U2694 (.Y(n3892), 
	.B1(n7699), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6314));
   INVX1 U2695 (.Y(n7699), 
	.A(\ram[206][14] ));
   OAI22X1 U2696 (.Y(n3891), 
	.B1(n7700), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6316));
   INVX1 U2697 (.Y(n7700), 
	.A(\ram[206][13] ));
   OAI22X1 U2698 (.Y(n3890), 
	.B1(n7701), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6318));
   INVX1 U2699 (.Y(n7701), 
	.A(\ram[206][12] ));
   OAI22X1 U2700 (.Y(n3889), 
	.B1(n7702), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6320));
   INVX1 U2701 (.Y(n7702), 
	.A(\ram[206][11] ));
   OAI22X1 U2702 (.Y(n3888), 
	.B1(n7703), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6322));
   INVX1 U2703 (.Y(n7703), 
	.A(\ram[206][10] ));
   OAI22X1 U2704 (.Y(n3887), 
	.B1(n7704), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6324));
   INVX1 U2705 (.Y(n7704), 
	.A(\ram[206][9] ));
   OAI22X1 U2706 (.Y(n3886), 
	.B1(n7705), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6326));
   INVX1 U2707 (.Y(n7705), 
	.A(\ram[206][8] ));
   OAI22X1 U2708 (.Y(n3885), 
	.B1(n7706), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6328));
   INVX1 U2709 (.Y(n7706), 
	.A(\ram[206][7] ));
   OAI22X1 U2710 (.Y(n3884), 
	.B1(n7707), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6330));
   INVX1 U2711 (.Y(n7707), 
	.A(\ram[206][6] ));
   OAI22X1 U2712 (.Y(n3883), 
	.B1(n7708), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6332));
   INVX1 U2713 (.Y(n7708), 
	.A(\ram[206][5] ));
   OAI22X1 U2714 (.Y(n3882), 
	.B1(n7709), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6334));
   INVX1 U2715 (.Y(n7709), 
	.A(\ram[206][4] ));
   OAI22X1 U2716 (.Y(n3881), 
	.B1(n7710), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6336));
   INVX1 U2717 (.Y(n7710), 
	.A(\ram[206][3] ));
   OAI22X1 U2718 (.Y(n3880), 
	.B1(n7711), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6338));
   INVX1 U2719 (.Y(n7711), 
	.A(\ram[206][2] ));
   OAI22X1 U2720 (.Y(n3879), 
	.B1(n7712), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6306));
   INVX1 U2721 (.Y(n7712), 
	.A(\ram[206][1] ));
   OAI22X1 U2722 (.Y(n3878), 
	.B1(n7713), 
	.B0(n7697), 
	.A1(n7696), 
	.A0(n6309));
   INVX1 U2723 (.Y(n7713), 
	.A(\ram[206][0] ));
   NOR2BX1 U2724 (.Y(n7697), 
	.B(n7696), 
	.AN(mem_write_en));
   NAND2X1 U2725 (.Y(n7696), 
	.B(n6553), 
	.A(n7695));
   OAI22X1 U2726 (.Y(n3877), 
	.B1(n7716), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6311));
   INVX1 U2727 (.Y(n7716), 
	.A(\ram[205][15] ));
   OAI22X1 U2728 (.Y(n3876), 
	.B1(n7717), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6314));
   INVX1 U2729 (.Y(n7717), 
	.A(\ram[205][14] ));
   OAI22X1 U2730 (.Y(n3875), 
	.B1(n7718), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6316));
   INVX1 U2731 (.Y(n7718), 
	.A(\ram[205][13] ));
   OAI22X1 U2732 (.Y(n3874), 
	.B1(n7719), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6318));
   INVX1 U2733 (.Y(n7719), 
	.A(\ram[205][12] ));
   OAI22X1 U2734 (.Y(n3873), 
	.B1(n7720), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6320));
   INVX1 U2735 (.Y(n7720), 
	.A(\ram[205][11] ));
   OAI22X1 U2736 (.Y(n3872), 
	.B1(n7721), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6322));
   INVX1 U2737 (.Y(n7721), 
	.A(\ram[205][10] ));
   OAI22X1 U2738 (.Y(n3871), 
	.B1(n7722), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6324));
   INVX1 U2739 (.Y(n7722), 
	.A(\ram[205][9] ));
   OAI22X1 U2740 (.Y(n3870), 
	.B1(n7723), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6326));
   INVX1 U2741 (.Y(n7723), 
	.A(\ram[205][8] ));
   OAI22X1 U2742 (.Y(n3869), 
	.B1(n7724), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6328));
   INVX1 U2743 (.Y(n7724), 
	.A(\ram[205][7] ));
   OAI22X1 U2744 (.Y(n3868), 
	.B1(n7725), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6330));
   INVX1 U2745 (.Y(n7725), 
	.A(\ram[205][6] ));
   OAI22X1 U2746 (.Y(n3867), 
	.B1(n7726), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6332));
   INVX1 U2747 (.Y(n7726), 
	.A(\ram[205][5] ));
   OAI22X1 U2748 (.Y(n3866), 
	.B1(n7727), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6334));
   INVX1 U2749 (.Y(n7727), 
	.A(\ram[205][4] ));
   OAI22X1 U2750 (.Y(n3865), 
	.B1(n7728), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6336));
   INVX1 U2751 (.Y(n7728), 
	.A(\ram[205][3] ));
   OAI22X1 U2752 (.Y(n3864), 
	.B1(n7729), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6338));
   INVX1 U2753 (.Y(n7729), 
	.A(\ram[205][2] ));
   OAI22X1 U2754 (.Y(n3863), 
	.B1(n7730), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6306));
   INVX1 U2755 (.Y(n7730), 
	.A(\ram[205][1] ));
   OAI22X1 U2756 (.Y(n3862), 
	.B1(n7731), 
	.B0(n7715), 
	.A1(n7714), 
	.A0(n6309));
   INVX1 U2757 (.Y(n7731), 
	.A(\ram[205][0] ));
   NOR2BX1 U2758 (.Y(n7715), 
	.B(n7714), 
	.AN(mem_write_en));
   NAND2X1 U2759 (.Y(n7714), 
	.B(n6572), 
	.A(n7695));
   OAI22X1 U2760 (.Y(n3861), 
	.B1(n7734), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6311));
   INVX1 U2761 (.Y(n7734), 
	.A(\ram[204][15] ));
   OAI22X1 U2762 (.Y(n3860), 
	.B1(n7735), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6314));
   INVX1 U2763 (.Y(n7735), 
	.A(\ram[204][14] ));
   OAI22X1 U2764 (.Y(n3859), 
	.B1(n7736), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6316));
   INVX1 U2765 (.Y(n7736), 
	.A(\ram[204][13] ));
   OAI22X1 U2766 (.Y(n3858), 
	.B1(n7737), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6318));
   INVX1 U2767 (.Y(n7737), 
	.A(\ram[204][12] ));
   OAI22X1 U2768 (.Y(n3857), 
	.B1(n7738), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6320));
   INVX1 U2769 (.Y(n7738), 
	.A(\ram[204][11] ));
   OAI22X1 U2770 (.Y(n3856), 
	.B1(n7739), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6322));
   INVX1 U2771 (.Y(n7739), 
	.A(\ram[204][10] ));
   OAI22X1 U2772 (.Y(n3855), 
	.B1(n7740), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6324));
   INVX1 U2773 (.Y(n7740), 
	.A(\ram[204][9] ));
   OAI22X1 U2774 (.Y(n3854), 
	.B1(n7741), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6326));
   INVX1 U2775 (.Y(n7741), 
	.A(\ram[204][8] ));
   OAI22X1 U2776 (.Y(n3853), 
	.B1(n7742), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6328));
   INVX1 U2777 (.Y(n7742), 
	.A(\ram[204][7] ));
   OAI22X1 U2778 (.Y(n3852), 
	.B1(n7743), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6330));
   INVX1 U2779 (.Y(n7743), 
	.A(\ram[204][6] ));
   OAI22X1 U2780 (.Y(n3851), 
	.B1(n7744), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6332));
   INVX1 U2781 (.Y(n7744), 
	.A(\ram[204][5] ));
   OAI22X1 U2782 (.Y(n3850), 
	.B1(n7745), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6334));
   INVX1 U2783 (.Y(n7745), 
	.A(\ram[204][4] ));
   OAI22X1 U2784 (.Y(n3849), 
	.B1(n7746), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6336));
   INVX1 U2785 (.Y(n7746), 
	.A(\ram[204][3] ));
   OAI22X1 U2786 (.Y(n3848), 
	.B1(n7747), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6338));
   INVX1 U2787 (.Y(n7747), 
	.A(\ram[204][2] ));
   OAI22X1 U2788 (.Y(n3847), 
	.B1(n7748), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6306));
   INVX1 U2789 (.Y(n7748), 
	.A(\ram[204][1] ));
   OAI22X1 U2790 (.Y(n3846), 
	.B1(n7749), 
	.B0(n7733), 
	.A1(n7732), 
	.A0(n6309));
   INVX1 U2791 (.Y(n7749), 
	.A(\ram[204][0] ));
   NOR2BX1 U2792 (.Y(n7733), 
	.B(n7732), 
	.AN(mem_write_en));
   NAND2X1 U2793 (.Y(n7732), 
	.B(n6591), 
	.A(n7695));
   OAI22X1 U2794 (.Y(n3845), 
	.B1(n7752), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6311));
   INVX1 U2795 (.Y(n7752), 
	.A(\ram[203][15] ));
   OAI22X1 U2796 (.Y(n3844), 
	.B1(n7753), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6314));
   INVX1 U2797 (.Y(n7753), 
	.A(\ram[203][14] ));
   OAI22X1 U2798 (.Y(n3843), 
	.B1(n7754), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6316));
   INVX1 U2799 (.Y(n7754), 
	.A(\ram[203][13] ));
   OAI22X1 U2800 (.Y(n3842), 
	.B1(n7755), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6318));
   INVX1 U2801 (.Y(n7755), 
	.A(\ram[203][12] ));
   OAI22X1 U2802 (.Y(n3841), 
	.B1(n7756), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6320));
   INVX1 U2803 (.Y(n7756), 
	.A(\ram[203][11] ));
   OAI22X1 U2804 (.Y(n3840), 
	.B1(n7757), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6322));
   INVX1 U2805 (.Y(n7757), 
	.A(\ram[203][10] ));
   OAI22X1 U2806 (.Y(n3839), 
	.B1(n7758), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6324));
   INVX1 U2807 (.Y(n7758), 
	.A(\ram[203][9] ));
   OAI22X1 U2808 (.Y(n3838), 
	.B1(n7759), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6326));
   INVX1 U2809 (.Y(n7759), 
	.A(\ram[203][8] ));
   OAI22X1 U2810 (.Y(n3837), 
	.B1(n7760), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6328));
   INVX1 U2811 (.Y(n7760), 
	.A(\ram[203][7] ));
   OAI22X1 U2812 (.Y(n3836), 
	.B1(n7761), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6330));
   INVX1 U2813 (.Y(n7761), 
	.A(\ram[203][6] ));
   OAI22X1 U2814 (.Y(n3835), 
	.B1(n7762), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6332));
   INVX1 U2815 (.Y(n7762), 
	.A(\ram[203][5] ));
   OAI22X1 U2816 (.Y(n3834), 
	.B1(n7763), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6334));
   INVX1 U2817 (.Y(n7763), 
	.A(\ram[203][4] ));
   OAI22X1 U2818 (.Y(n3833), 
	.B1(n7764), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6336));
   INVX1 U2819 (.Y(n7764), 
	.A(\ram[203][3] ));
   OAI22X1 U2820 (.Y(n3832), 
	.B1(n7765), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6338));
   INVX1 U2821 (.Y(n7765), 
	.A(\ram[203][2] ));
   OAI22X1 U2822 (.Y(n3831), 
	.B1(n7766), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6306));
   INVX1 U2823 (.Y(n7766), 
	.A(\ram[203][1] ));
   OAI22X1 U2824 (.Y(n3830), 
	.B1(n7767), 
	.B0(n7751), 
	.A1(n7750), 
	.A0(n6309));
   INVX1 U2825 (.Y(n7767), 
	.A(\ram[203][0] ));
   NOR2BX1 U2826 (.Y(n7751), 
	.B(n7750), 
	.AN(mem_write_en));
   NAND2X1 U2827 (.Y(n7750), 
	.B(n6610), 
	.A(n7695));
   OAI22X1 U2828 (.Y(n3829), 
	.B1(n7770), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6311));
   INVX1 U2829 (.Y(n7770), 
	.A(\ram[202][15] ));
   OAI22X1 U2830 (.Y(n3828), 
	.B1(n7771), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6314));
   INVX1 U2831 (.Y(n7771), 
	.A(\ram[202][14] ));
   OAI22X1 U2832 (.Y(n3827), 
	.B1(n7772), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6316));
   INVX1 U2833 (.Y(n7772), 
	.A(\ram[202][13] ));
   OAI22X1 U2834 (.Y(n3826), 
	.B1(n7773), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6318));
   INVX1 U2835 (.Y(n7773), 
	.A(\ram[202][12] ));
   OAI22X1 U2836 (.Y(n3825), 
	.B1(n7774), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6320));
   INVX1 U2837 (.Y(n7774), 
	.A(\ram[202][11] ));
   OAI22X1 U2838 (.Y(n3824), 
	.B1(n7775), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6322));
   INVX1 U2839 (.Y(n7775), 
	.A(\ram[202][10] ));
   OAI22X1 U2840 (.Y(n3823), 
	.B1(n7776), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6324));
   INVX1 U2841 (.Y(n7776), 
	.A(\ram[202][9] ));
   OAI22X1 U2842 (.Y(n3822), 
	.B1(n7777), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6326));
   INVX1 U2843 (.Y(n7777), 
	.A(\ram[202][8] ));
   OAI22X1 U2844 (.Y(n3821), 
	.B1(n7778), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6328));
   INVX1 U2845 (.Y(n7778), 
	.A(\ram[202][7] ));
   OAI22X1 U2846 (.Y(n3820), 
	.B1(n7779), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6330));
   INVX1 U2847 (.Y(n7779), 
	.A(\ram[202][6] ));
   OAI22X1 U2848 (.Y(n3819), 
	.B1(n7780), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6332));
   INVX1 U2849 (.Y(n7780), 
	.A(\ram[202][5] ));
   OAI22X1 U2850 (.Y(n3818), 
	.B1(n7781), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6334));
   INVX1 U2851 (.Y(n7781), 
	.A(\ram[202][4] ));
   OAI22X1 U2852 (.Y(n3817), 
	.B1(n7782), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6336));
   INVX1 U2853 (.Y(n7782), 
	.A(\ram[202][3] ));
   OAI22X1 U2854 (.Y(n3816), 
	.B1(n7783), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6338));
   INVX1 U2855 (.Y(n7783), 
	.A(\ram[202][2] ));
   OAI22X1 U2856 (.Y(n3815), 
	.B1(n7784), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6306));
   INVX1 U2857 (.Y(n7784), 
	.A(\ram[202][1] ));
   OAI22X1 U2858 (.Y(n3814), 
	.B1(n7785), 
	.B0(n7769), 
	.A1(n7768), 
	.A0(n6309));
   INVX1 U2859 (.Y(n7785), 
	.A(\ram[202][0] ));
   NOR2BX1 U2860 (.Y(n7769), 
	.B(n7768), 
	.AN(mem_write_en));
   NAND2X1 U2861 (.Y(n7768), 
	.B(n6629), 
	.A(n7695));
   OAI22X1 U2862 (.Y(n3813), 
	.B1(n7788), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6311));
   INVX1 U2863 (.Y(n7788), 
	.A(\ram[201][15] ));
   OAI22X1 U2864 (.Y(n3812), 
	.B1(n7789), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6314));
   INVX1 U2865 (.Y(n7789), 
	.A(\ram[201][14] ));
   OAI22X1 U2866 (.Y(n3811), 
	.B1(n7790), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6316));
   INVX1 U2867 (.Y(n7790), 
	.A(\ram[201][13] ));
   OAI22X1 U2868 (.Y(n3810), 
	.B1(n7791), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6318));
   INVX1 U2869 (.Y(n7791), 
	.A(\ram[201][12] ));
   OAI22X1 U2870 (.Y(n3809), 
	.B1(n7792), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6320));
   INVX1 U2871 (.Y(n7792), 
	.A(\ram[201][11] ));
   OAI22X1 U2872 (.Y(n3808), 
	.B1(n7793), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6322));
   INVX1 U2873 (.Y(n7793), 
	.A(\ram[201][10] ));
   OAI22X1 U2874 (.Y(n3807), 
	.B1(n7794), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6324));
   INVX1 U2875 (.Y(n7794), 
	.A(\ram[201][9] ));
   OAI22X1 U2876 (.Y(n3806), 
	.B1(n7795), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6326));
   INVX1 U2877 (.Y(n7795), 
	.A(\ram[201][8] ));
   OAI22X1 U2878 (.Y(n3805), 
	.B1(n7796), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6328));
   INVX1 U2879 (.Y(n7796), 
	.A(\ram[201][7] ));
   OAI22X1 U2880 (.Y(n3804), 
	.B1(n7797), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6330));
   INVX1 U2881 (.Y(n7797), 
	.A(\ram[201][6] ));
   OAI22X1 U2882 (.Y(n3803), 
	.B1(n7798), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6332));
   INVX1 U2883 (.Y(n7798), 
	.A(\ram[201][5] ));
   OAI22X1 U2884 (.Y(n3802), 
	.B1(n7799), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6334));
   INVX1 U2885 (.Y(n7799), 
	.A(\ram[201][4] ));
   OAI22X1 U2886 (.Y(n3801), 
	.B1(n7800), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6336));
   INVX1 U2887 (.Y(n7800), 
	.A(\ram[201][3] ));
   OAI22X1 U2888 (.Y(n3800), 
	.B1(n7801), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6338));
   INVX1 U2889 (.Y(n7801), 
	.A(\ram[201][2] ));
   OAI22X1 U2890 (.Y(n3799), 
	.B1(n7802), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6306));
   INVX1 U2891 (.Y(n7802), 
	.A(\ram[201][1] ));
   OAI22X1 U2892 (.Y(n3798), 
	.B1(n7803), 
	.B0(n7787), 
	.A1(n7786), 
	.A0(n6309));
   INVX1 U2893 (.Y(n7803), 
	.A(\ram[201][0] ));
   NOR2BX1 U2894 (.Y(n7787), 
	.B(n7786), 
	.AN(mem_write_en));
   NAND2X1 U2895 (.Y(n7786), 
	.B(n6342), 
	.A(n7695));
   OAI22X1 U2896 (.Y(n3797), 
	.B1(n7806), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6311));
   INVX1 U2897 (.Y(n7806), 
	.A(\ram[200][15] ));
   OAI22X1 U2898 (.Y(n3796), 
	.B1(n7807), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6314));
   INVX1 U2899 (.Y(n7807), 
	.A(\ram[200][14] ));
   OAI22X1 U2900 (.Y(n3795), 
	.B1(n7808), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6316));
   INVX1 U2901 (.Y(n7808), 
	.A(\ram[200][13] ));
   OAI22X1 U2902 (.Y(n3794), 
	.B1(n7809), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6318));
   INVX1 U2903 (.Y(n7809), 
	.A(\ram[200][12] ));
   OAI22X1 U2904 (.Y(n3793), 
	.B1(n7810), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6320));
   INVX1 U2905 (.Y(n7810), 
	.A(\ram[200][11] ));
   OAI22X1 U2906 (.Y(n3792), 
	.B1(n7811), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6322));
   INVX1 U2907 (.Y(n7811), 
	.A(\ram[200][10] ));
   OAI22X1 U2908 (.Y(n3791), 
	.B1(n7812), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6324));
   INVX1 U2909 (.Y(n7812), 
	.A(\ram[200][9] ));
   OAI22X1 U2910 (.Y(n3790), 
	.B1(n7813), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6326));
   INVX1 U2911 (.Y(n7813), 
	.A(\ram[200][8] ));
   OAI22X1 U2912 (.Y(n3789), 
	.B1(n7814), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6328));
   INVX1 U2913 (.Y(n7814), 
	.A(\ram[200][7] ));
   OAI22X1 U2914 (.Y(n3788), 
	.B1(n7815), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6330));
   INVX1 U2915 (.Y(n7815), 
	.A(\ram[200][6] ));
   OAI22X1 U2916 (.Y(n3787), 
	.B1(n7816), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6332));
   INVX1 U2917 (.Y(n7816), 
	.A(\ram[200][5] ));
   OAI22X1 U2918 (.Y(n3786), 
	.B1(n7817), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6334));
   INVX1 U2919 (.Y(n7817), 
	.A(\ram[200][4] ));
   OAI22X1 U2920 (.Y(n3785), 
	.B1(n7818), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6336));
   INVX1 U2921 (.Y(n7818), 
	.A(\ram[200][3] ));
   OAI22X1 U2922 (.Y(n3784), 
	.B1(n7819), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6338));
   INVX1 U2923 (.Y(n7819), 
	.A(\ram[200][2] ));
   OAI22X1 U2924 (.Y(n3783), 
	.B1(n7820), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6306));
   INVX1 U2925 (.Y(n7820), 
	.A(\ram[200][1] ));
   OAI22X1 U2926 (.Y(n3782), 
	.B1(n7821), 
	.B0(n7805), 
	.A1(n7804), 
	.A0(n6309));
   INVX1 U2927 (.Y(n7821), 
	.A(\ram[200][0] ));
   NOR2BX1 U2928 (.Y(n7805), 
	.B(n7804), 
	.AN(mem_write_en));
   NAND2X1 U2929 (.Y(n7804), 
	.B(n6362), 
	.A(n7695));
   OAI22X1 U2930 (.Y(n3781), 
	.B1(n7824), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6311));
   INVX1 U2931 (.Y(n7824), 
	.A(\ram[199][15] ));
   OAI22X1 U2932 (.Y(n3780), 
	.B1(n7825), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6314));
   INVX1 U2933 (.Y(n7825), 
	.A(\ram[199][14] ));
   OAI22X1 U2934 (.Y(n3779), 
	.B1(n7826), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6316));
   INVX1 U2935 (.Y(n7826), 
	.A(\ram[199][13] ));
   OAI22X1 U2936 (.Y(n3778), 
	.B1(n7827), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6318));
   INVX1 U2937 (.Y(n7827), 
	.A(\ram[199][12] ));
   OAI22X1 U2938 (.Y(n3777), 
	.B1(n7828), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6320));
   INVX1 U2939 (.Y(n7828), 
	.A(\ram[199][11] ));
   OAI22X1 U2940 (.Y(n3776), 
	.B1(n7829), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6322));
   INVX1 U2941 (.Y(n7829), 
	.A(\ram[199][10] ));
   OAI22X1 U2942 (.Y(n3775), 
	.B1(n7830), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6324));
   INVX1 U2943 (.Y(n7830), 
	.A(\ram[199][9] ));
   OAI22X1 U2944 (.Y(n3774), 
	.B1(n7831), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6326));
   INVX1 U2945 (.Y(n7831), 
	.A(\ram[199][8] ));
   OAI22X1 U2946 (.Y(n3773), 
	.B1(n7832), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6328));
   INVX1 U2947 (.Y(n7832), 
	.A(\ram[199][7] ));
   OAI22X1 U2948 (.Y(n3772), 
	.B1(n7833), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6330));
   INVX1 U2949 (.Y(n7833), 
	.A(\ram[199][6] ));
   OAI22X1 U2950 (.Y(n3771), 
	.B1(n7834), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6332));
   INVX1 U2951 (.Y(n7834), 
	.A(\ram[199][5] ));
   OAI22X1 U2952 (.Y(n3770), 
	.B1(n7835), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6334));
   INVX1 U2953 (.Y(n7835), 
	.A(\ram[199][4] ));
   OAI22X1 U2954 (.Y(n3769), 
	.B1(n7836), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6336));
   INVX1 U2955 (.Y(n7836), 
	.A(\ram[199][3] ));
   OAI22X1 U2956 (.Y(n3768), 
	.B1(n7837), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6338));
   INVX1 U2957 (.Y(n7837), 
	.A(\ram[199][2] ));
   OAI22X1 U2958 (.Y(n3767), 
	.B1(n7838), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6306));
   INVX1 U2959 (.Y(n7838), 
	.A(\ram[199][1] ));
   OAI22X1 U2960 (.Y(n3766), 
	.B1(n7839), 
	.B0(n7823), 
	.A1(n7822), 
	.A0(n6309));
   INVX1 U2961 (.Y(n7839), 
	.A(\ram[199][0] ));
   NOR2BX1 U2962 (.Y(n7823), 
	.B(n7822), 
	.AN(mem_write_en));
   NAND2X1 U2963 (.Y(n7822), 
	.B(n6381), 
	.A(n7695));
   OAI22X1 U2964 (.Y(n3765), 
	.B1(n7842), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6311));
   INVX1 U2965 (.Y(n7842), 
	.A(\ram[198][15] ));
   OAI22X1 U2966 (.Y(n3764), 
	.B1(n7843), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6314));
   INVX1 U2967 (.Y(n7843), 
	.A(\ram[198][14] ));
   OAI22X1 U2968 (.Y(n3763), 
	.B1(n7844), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6316));
   INVX1 U2969 (.Y(n7844), 
	.A(\ram[198][13] ));
   OAI22X1 U2970 (.Y(n3762), 
	.B1(n7845), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6318));
   INVX1 U2971 (.Y(n7845), 
	.A(\ram[198][12] ));
   OAI22X1 U2972 (.Y(n3761), 
	.B1(n7846), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6320));
   INVX1 U2973 (.Y(n7846), 
	.A(\ram[198][11] ));
   OAI22X1 U2974 (.Y(n3760), 
	.B1(n7847), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6322));
   INVX1 U2975 (.Y(n7847), 
	.A(\ram[198][10] ));
   OAI22X1 U2976 (.Y(n3759), 
	.B1(n7848), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6324));
   INVX1 U2977 (.Y(n7848), 
	.A(\ram[198][9] ));
   OAI22X1 U2978 (.Y(n3758), 
	.B1(n7849), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6326));
   INVX1 U2979 (.Y(n7849), 
	.A(\ram[198][8] ));
   OAI22X1 U2980 (.Y(n3757), 
	.B1(n7850), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6328));
   INVX1 U2981 (.Y(n7850), 
	.A(\ram[198][7] ));
   OAI22X1 U2982 (.Y(n3756), 
	.B1(n7851), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6330));
   INVX1 U2983 (.Y(n7851), 
	.A(\ram[198][6] ));
   OAI22X1 U2984 (.Y(n3755), 
	.B1(n7852), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6332));
   INVX1 U2985 (.Y(n7852), 
	.A(\ram[198][5] ));
   OAI22X1 U2986 (.Y(n3754), 
	.B1(n7853), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6334));
   INVX1 U2987 (.Y(n7853), 
	.A(\ram[198][4] ));
   OAI22X1 U2988 (.Y(n3753), 
	.B1(n7854), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6336));
   INVX1 U2989 (.Y(n7854), 
	.A(\ram[198][3] ));
   OAI22X1 U2990 (.Y(n3752), 
	.B1(n7855), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6338));
   INVX1 U2991 (.Y(n7855), 
	.A(\ram[198][2] ));
   OAI22X1 U2992 (.Y(n3751), 
	.B1(n7856), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6306));
   INVX1 U2993 (.Y(n7856), 
	.A(\ram[198][1] ));
   OAI22X1 U2994 (.Y(n3750), 
	.B1(n7857), 
	.B0(n7841), 
	.A1(n7840), 
	.A0(n6309));
   INVX1 U2995 (.Y(n7857), 
	.A(\ram[198][0] ));
   NOR2BX1 U2996 (.Y(n7841), 
	.B(n7840), 
	.AN(mem_write_en));
   NAND2X1 U2997 (.Y(n7840), 
	.B(n6400), 
	.A(n7695));
   OAI22X1 U2998 (.Y(n3749), 
	.B1(n7860), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6311));
   INVX1 U2999 (.Y(n7860), 
	.A(\ram[197][15] ));
   OAI22X1 U3000 (.Y(n3748), 
	.B1(n7861), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6314));
   INVX1 U3001 (.Y(n7861), 
	.A(\ram[197][14] ));
   OAI22X1 U3002 (.Y(n3747), 
	.B1(n7862), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6316));
   INVX1 U3003 (.Y(n7862), 
	.A(\ram[197][13] ));
   OAI22X1 U3004 (.Y(n3746), 
	.B1(n7863), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6318));
   INVX1 U3005 (.Y(n7863), 
	.A(\ram[197][12] ));
   OAI22X1 U3006 (.Y(n3745), 
	.B1(n7864), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6320));
   INVX1 U3007 (.Y(n7864), 
	.A(\ram[197][11] ));
   OAI22X1 U3008 (.Y(n3744), 
	.B1(n7865), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6322));
   INVX1 U3009 (.Y(n7865), 
	.A(\ram[197][10] ));
   OAI22X1 U3010 (.Y(n3743), 
	.B1(n7866), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6324));
   INVX1 U3011 (.Y(n7866), 
	.A(\ram[197][9] ));
   OAI22X1 U3012 (.Y(n3742), 
	.B1(n7867), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6326));
   INVX1 U3013 (.Y(n7867), 
	.A(\ram[197][8] ));
   OAI22X1 U3014 (.Y(n3741), 
	.B1(n7868), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6328));
   INVX1 U3015 (.Y(n7868), 
	.A(\ram[197][7] ));
   OAI22X1 U3016 (.Y(n3740), 
	.B1(n7869), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6330));
   INVX1 U3017 (.Y(n7869), 
	.A(\ram[197][6] ));
   OAI22X1 U3018 (.Y(n3739), 
	.B1(n7870), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6332));
   INVX1 U3019 (.Y(n7870), 
	.A(\ram[197][5] ));
   OAI22X1 U3020 (.Y(n3738), 
	.B1(n7871), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6334));
   INVX1 U3021 (.Y(n7871), 
	.A(\ram[197][4] ));
   OAI22X1 U3022 (.Y(n3737), 
	.B1(n7872), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6336));
   INVX1 U3023 (.Y(n7872), 
	.A(\ram[197][3] ));
   OAI22X1 U3024 (.Y(n3736), 
	.B1(n7873), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6338));
   INVX1 U3025 (.Y(n7873), 
	.A(\ram[197][2] ));
   OAI22X1 U3026 (.Y(n3735), 
	.B1(n7874), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6306));
   INVX1 U3027 (.Y(n7874), 
	.A(\ram[197][1] ));
   OAI22X1 U3028 (.Y(n3734), 
	.B1(n7875), 
	.B0(n7859), 
	.A1(n7858), 
	.A0(n6309));
   INVX1 U3029 (.Y(n7875), 
	.A(\ram[197][0] ));
   NOR2BX1 U3030 (.Y(n7859), 
	.B(n7858), 
	.AN(mem_write_en));
   NAND2X1 U3031 (.Y(n7858), 
	.B(n6419), 
	.A(n7695));
   OAI22X1 U3032 (.Y(n3733), 
	.B1(n7878), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6311));
   INVX1 U3033 (.Y(n7878), 
	.A(\ram[196][15] ));
   OAI22X1 U3034 (.Y(n3732), 
	.B1(n7879), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6314));
   INVX1 U3035 (.Y(n7879), 
	.A(\ram[196][14] ));
   OAI22X1 U3036 (.Y(n3731), 
	.B1(n7880), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6316));
   INVX1 U3037 (.Y(n7880), 
	.A(\ram[196][13] ));
   OAI22X1 U3038 (.Y(n3730), 
	.B1(n7881), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6318));
   INVX1 U3039 (.Y(n7881), 
	.A(\ram[196][12] ));
   OAI22X1 U3040 (.Y(n3729), 
	.B1(n7882), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6320));
   INVX1 U3041 (.Y(n7882), 
	.A(\ram[196][11] ));
   OAI22X1 U3042 (.Y(n3728), 
	.B1(n7883), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6322));
   INVX1 U3043 (.Y(n7883), 
	.A(\ram[196][10] ));
   OAI22X1 U3044 (.Y(n3727), 
	.B1(n7884), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6324));
   INVX1 U3045 (.Y(n7884), 
	.A(\ram[196][9] ));
   OAI22X1 U3046 (.Y(n3726), 
	.B1(n7885), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6326));
   INVX1 U3047 (.Y(n7885), 
	.A(\ram[196][8] ));
   OAI22X1 U3048 (.Y(n3725), 
	.B1(n7886), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6328));
   INVX1 U3049 (.Y(n7886), 
	.A(\ram[196][7] ));
   OAI22X1 U3050 (.Y(n3724), 
	.B1(n7887), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6330));
   INVX1 U3051 (.Y(n7887), 
	.A(\ram[196][6] ));
   OAI22X1 U3052 (.Y(n3723), 
	.B1(n7888), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6332));
   INVX1 U3053 (.Y(n7888), 
	.A(\ram[196][5] ));
   OAI22X1 U3054 (.Y(n3722), 
	.B1(n7889), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6334));
   INVX1 U3055 (.Y(n7889), 
	.A(\ram[196][4] ));
   OAI22X1 U3056 (.Y(n3721), 
	.B1(n7890), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6336));
   INVX1 U3057 (.Y(n7890), 
	.A(\ram[196][3] ));
   OAI22X1 U3058 (.Y(n3720), 
	.B1(n7891), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6338));
   INVX1 U3059 (.Y(n7891), 
	.A(\ram[196][2] ));
   OAI22X1 U3060 (.Y(n3719), 
	.B1(n7892), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6306));
   INVX1 U3061 (.Y(n7892), 
	.A(\ram[196][1] ));
   OAI22X1 U3062 (.Y(n3718), 
	.B1(n7893), 
	.B0(n7877), 
	.A1(n7876), 
	.A0(n6309));
   INVX1 U3063 (.Y(n7893), 
	.A(\ram[196][0] ));
   NOR2BX1 U3064 (.Y(n7877), 
	.B(n7876), 
	.AN(mem_write_en));
   NAND2X1 U3065 (.Y(n7876), 
	.B(n6438), 
	.A(n7695));
   OAI22X1 U3066 (.Y(n3717), 
	.B1(n7896), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6311));
   INVX1 U3067 (.Y(n7896), 
	.A(\ram[195][15] ));
   OAI22X1 U3068 (.Y(n3716), 
	.B1(n7897), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6314));
   INVX1 U3069 (.Y(n7897), 
	.A(\ram[195][14] ));
   OAI22X1 U3070 (.Y(n3715), 
	.B1(n7898), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6316));
   INVX1 U3071 (.Y(n7898), 
	.A(\ram[195][13] ));
   OAI22X1 U3072 (.Y(n3714), 
	.B1(n7899), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6318));
   INVX1 U3073 (.Y(n7899), 
	.A(\ram[195][12] ));
   OAI22X1 U3074 (.Y(n3713), 
	.B1(n7900), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6320));
   INVX1 U3075 (.Y(n7900), 
	.A(\ram[195][11] ));
   OAI22X1 U3076 (.Y(n3712), 
	.B1(n7901), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6322));
   INVX1 U3077 (.Y(n7901), 
	.A(\ram[195][10] ));
   OAI22X1 U3078 (.Y(n3711), 
	.B1(n7902), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6324));
   INVX1 U3079 (.Y(n7902), 
	.A(\ram[195][9] ));
   OAI22X1 U3080 (.Y(n3710), 
	.B1(n7903), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6326));
   INVX1 U3081 (.Y(n7903), 
	.A(\ram[195][8] ));
   OAI22X1 U3082 (.Y(n3709), 
	.B1(n7904), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6328));
   INVX1 U3083 (.Y(n7904), 
	.A(\ram[195][7] ));
   OAI22X1 U3084 (.Y(n3708), 
	.B1(n7905), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6330));
   INVX1 U3085 (.Y(n7905), 
	.A(\ram[195][6] ));
   OAI22X1 U3086 (.Y(n3707), 
	.B1(n7906), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6332));
   INVX1 U3087 (.Y(n7906), 
	.A(\ram[195][5] ));
   OAI22X1 U3088 (.Y(n3706), 
	.B1(n7907), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6334));
   INVX1 U3089 (.Y(n7907), 
	.A(\ram[195][4] ));
   OAI22X1 U3090 (.Y(n3705), 
	.B1(n7908), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6336));
   INVX1 U3091 (.Y(n7908), 
	.A(\ram[195][3] ));
   OAI22X1 U3092 (.Y(n3704), 
	.B1(n7909), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6338));
   INVX1 U3093 (.Y(n7909), 
	.A(\ram[195][2] ));
   OAI22X1 U3094 (.Y(n3703), 
	.B1(n7910), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6306));
   INVX1 U3095 (.Y(n7910), 
	.A(\ram[195][1] ));
   OAI22X1 U3096 (.Y(n3702), 
	.B1(n7911), 
	.B0(n7895), 
	.A1(n7894), 
	.A0(n6309));
   INVX1 U3097 (.Y(n7911), 
	.A(\ram[195][0] ));
   NOR2BX1 U3098 (.Y(n7895), 
	.B(n7894), 
	.AN(mem_write_en));
   NAND2X1 U3099 (.Y(n7894), 
	.B(n6457), 
	.A(n7695));
   OAI22X1 U3100 (.Y(n3701), 
	.B1(n7914), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6311));
   INVX1 U3101 (.Y(n7914), 
	.A(\ram[194][15] ));
   OAI22X1 U3102 (.Y(n3700), 
	.B1(n7915), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6314));
   INVX1 U3103 (.Y(n7915), 
	.A(\ram[194][14] ));
   OAI22X1 U3104 (.Y(n3699), 
	.B1(n7916), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6316));
   INVX1 U3105 (.Y(n7916), 
	.A(\ram[194][13] ));
   OAI22X1 U3106 (.Y(n3698), 
	.B1(n7917), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6318));
   INVX1 U3107 (.Y(n7917), 
	.A(\ram[194][12] ));
   OAI22X1 U3108 (.Y(n3697), 
	.B1(n7918), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6320));
   INVX1 U3109 (.Y(n7918), 
	.A(\ram[194][11] ));
   OAI22X1 U3110 (.Y(n3696), 
	.B1(n7919), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6322));
   INVX1 U3111 (.Y(n7919), 
	.A(\ram[194][10] ));
   OAI22X1 U3112 (.Y(n3695), 
	.B1(n7920), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6324));
   INVX1 U3113 (.Y(n7920), 
	.A(\ram[194][9] ));
   OAI22X1 U3114 (.Y(n3694), 
	.B1(n7921), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6326));
   INVX1 U3115 (.Y(n7921), 
	.A(\ram[194][8] ));
   OAI22X1 U3116 (.Y(n3693), 
	.B1(n7922), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6328));
   INVX1 U3117 (.Y(n7922), 
	.A(\ram[194][7] ));
   OAI22X1 U3118 (.Y(n3692), 
	.B1(n7923), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6330));
   INVX1 U3119 (.Y(n7923), 
	.A(\ram[194][6] ));
   OAI22X1 U3120 (.Y(n3691), 
	.B1(n7924), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6332));
   INVX1 U3121 (.Y(n7924), 
	.A(\ram[194][5] ));
   OAI22X1 U3122 (.Y(n3690), 
	.B1(n7925), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6334));
   INVX1 U3123 (.Y(n7925), 
	.A(\ram[194][4] ));
   OAI22X1 U3124 (.Y(n3689), 
	.B1(n7926), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6336));
   INVX1 U3125 (.Y(n7926), 
	.A(\ram[194][3] ));
   OAI22X1 U3126 (.Y(n3688), 
	.B1(n7927), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6338));
   INVX1 U3127 (.Y(n7927), 
	.A(\ram[194][2] ));
   OAI22X1 U3128 (.Y(n3687), 
	.B1(n7928), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6306));
   INVX1 U3129 (.Y(n7928), 
	.A(\ram[194][1] ));
   OAI22X1 U3130 (.Y(n3686), 
	.B1(n7929), 
	.B0(n7913), 
	.A1(n7912), 
	.A0(n6309));
   INVX1 U3131 (.Y(n7929), 
	.A(\ram[194][0] ));
   NOR2BX1 U3132 (.Y(n7913), 
	.B(n7912), 
	.AN(mem_write_en));
   NAND2X1 U3133 (.Y(n7912), 
	.B(n6476), 
	.A(n7695));
   OAI22X1 U3134 (.Y(n3685), 
	.B1(n7932), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6311));
   INVX1 U3135 (.Y(n7932), 
	.A(\ram[193][15] ));
   OAI22X1 U3136 (.Y(n3684), 
	.B1(n7933), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6314));
   INVX1 U3137 (.Y(n7933), 
	.A(\ram[193][14] ));
   OAI22X1 U3138 (.Y(n3683), 
	.B1(n7934), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6316));
   INVX1 U3139 (.Y(n7934), 
	.A(\ram[193][13] ));
   OAI22X1 U3140 (.Y(n3682), 
	.B1(n7935), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6318));
   INVX1 U3141 (.Y(n7935), 
	.A(\ram[193][12] ));
   OAI22X1 U3142 (.Y(n3681), 
	.B1(n7936), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6320));
   INVX1 U3143 (.Y(n7936), 
	.A(\ram[193][11] ));
   OAI22X1 U3144 (.Y(n3680), 
	.B1(n7937), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6322));
   INVX1 U3145 (.Y(n7937), 
	.A(\ram[193][10] ));
   OAI22X1 U3146 (.Y(n3679), 
	.B1(n7938), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6324));
   INVX1 U3147 (.Y(n7938), 
	.A(\ram[193][9] ));
   OAI22X1 U3148 (.Y(n3678), 
	.B1(n7939), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6326));
   INVX1 U3149 (.Y(n7939), 
	.A(\ram[193][8] ));
   OAI22X1 U3150 (.Y(n3677), 
	.B1(n7940), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6328));
   INVX1 U3151 (.Y(n7940), 
	.A(\ram[193][7] ));
   OAI22X1 U3152 (.Y(n3676), 
	.B1(n7941), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6330));
   INVX1 U3153 (.Y(n7941), 
	.A(\ram[193][6] ));
   OAI22X1 U3154 (.Y(n3675), 
	.B1(n7942), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6332));
   INVX1 U3155 (.Y(n7942), 
	.A(\ram[193][5] ));
   OAI22X1 U3156 (.Y(n3674), 
	.B1(n7943), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6334));
   INVX1 U3157 (.Y(n7943), 
	.A(\ram[193][4] ));
   OAI22X1 U3158 (.Y(n3673), 
	.B1(n7944), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6336));
   INVX1 U3159 (.Y(n7944), 
	.A(\ram[193][3] ));
   OAI22X1 U3160 (.Y(n3672), 
	.B1(n7945), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6338));
   INVX1 U3161 (.Y(n7945), 
	.A(\ram[193][2] ));
   OAI22X1 U3162 (.Y(n3671), 
	.B1(n7946), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6306));
   INVX1 U3163 (.Y(n7946), 
	.A(\ram[193][1] ));
   OAI22X1 U3164 (.Y(n3670), 
	.B1(n7947), 
	.B0(n7931), 
	.A1(n7930), 
	.A0(n6309));
   INVX1 U3165 (.Y(n7947), 
	.A(\ram[193][0] ));
   NOR2BX1 U3166 (.Y(n7931), 
	.B(n7930), 
	.AN(mem_write_en));
   NAND2X1 U3167 (.Y(n7930), 
	.B(n6495), 
	.A(n7695));
   OAI22X1 U3168 (.Y(n3669), 
	.B1(n7950), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6311));
   INVX1 U3169 (.Y(n7950), 
	.A(\ram[192][15] ));
   OAI22X1 U3170 (.Y(n3668), 
	.B1(n7951), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6314));
   INVX1 U3171 (.Y(n7951), 
	.A(\ram[192][14] ));
   OAI22X1 U3172 (.Y(n3667), 
	.B1(n7952), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6316));
   INVX1 U3173 (.Y(n7952), 
	.A(\ram[192][13] ));
   OAI22X1 U3174 (.Y(n3666), 
	.B1(n7953), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6318));
   INVX1 U3175 (.Y(n7953), 
	.A(\ram[192][12] ));
   OAI22X1 U3176 (.Y(n3665), 
	.B1(n7954), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6320));
   INVX1 U3177 (.Y(n7954), 
	.A(\ram[192][11] ));
   OAI22X1 U3178 (.Y(n3664), 
	.B1(n7955), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6322));
   INVX1 U3179 (.Y(n7955), 
	.A(\ram[192][10] ));
   OAI22X1 U3180 (.Y(n3663), 
	.B1(n7956), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6324));
   INVX1 U3181 (.Y(n7956), 
	.A(\ram[192][9] ));
   OAI22X1 U3182 (.Y(n3662), 
	.B1(n7957), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6326));
   INVX1 U3183 (.Y(n7957), 
	.A(\ram[192][8] ));
   OAI22X1 U3184 (.Y(n3661), 
	.B1(n7958), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6328));
   INVX1 U3185 (.Y(n7958), 
	.A(\ram[192][7] ));
   OAI22X1 U3186 (.Y(n3660), 
	.B1(n7959), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6330));
   INVX1 U3187 (.Y(n7959), 
	.A(\ram[192][6] ));
   OAI22X1 U3188 (.Y(n3659), 
	.B1(n7960), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6332));
   INVX1 U3189 (.Y(n7960), 
	.A(\ram[192][5] ));
   OAI22X1 U3190 (.Y(n3658), 
	.B1(n7961), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6334));
   INVX1 U3191 (.Y(n7961), 
	.A(\ram[192][4] ));
   OAI22X1 U3192 (.Y(n3657), 
	.B1(n7962), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6336));
   INVX1 U3193 (.Y(n7962), 
	.A(\ram[192][3] ));
   OAI22X1 U3194 (.Y(n3656), 
	.B1(n7963), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6338));
   INVX1 U3195 (.Y(n7963), 
	.A(\ram[192][2] ));
   OAI22X1 U3196 (.Y(n3655), 
	.B1(n7964), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6306));
   INVX1 U3197 (.Y(n7964), 
	.A(\ram[192][1] ));
   OAI22X1 U3198 (.Y(n3654), 
	.B1(n7965), 
	.B0(n7949), 
	.A1(n7948), 
	.A0(n6309));
   INVX1 U3199 (.Y(n7965), 
	.A(\ram[192][0] ));
   NOR2BX1 U3200 (.Y(n7949), 
	.B(n7948), 
	.AN(mem_write_en));
   NAND2X1 U3201 (.Y(n7948), 
	.B(n6514), 
	.A(n7695));
   OAI22X1 U3202 (.Y(n3653), 
	.B1(n7968), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6311));
   INVX1 U3203 (.Y(n7968), 
	.A(\ram[191][15] ));
   OAI22X1 U3204 (.Y(n3652), 
	.B1(n7969), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6314));
   INVX1 U3205 (.Y(n7969), 
	.A(\ram[191][14] ));
   OAI22X1 U3206 (.Y(n3651), 
	.B1(n7970), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6316));
   INVX1 U3207 (.Y(n7970), 
	.A(\ram[191][13] ));
   OAI22X1 U3208 (.Y(n3650), 
	.B1(n7971), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6318));
   INVX1 U3209 (.Y(n7971), 
	.A(\ram[191][12] ));
   OAI22X1 U3210 (.Y(n3649), 
	.B1(n7972), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6320));
   INVX1 U3211 (.Y(n7972), 
	.A(\ram[191][11] ));
   OAI22X1 U3212 (.Y(n3648), 
	.B1(n7973), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6322));
   INVX1 U3213 (.Y(n7973), 
	.A(\ram[191][10] ));
   OAI22X1 U3214 (.Y(n3647), 
	.B1(n7974), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6324));
   INVX1 U3215 (.Y(n7974), 
	.A(\ram[191][9] ));
   OAI22X1 U3216 (.Y(n3646), 
	.B1(n7975), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6326));
   INVX1 U3217 (.Y(n7975), 
	.A(\ram[191][8] ));
   OAI22X1 U3218 (.Y(n3645), 
	.B1(n7976), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6328));
   INVX1 U3219 (.Y(n7976), 
	.A(\ram[191][7] ));
   OAI22X1 U3220 (.Y(n3644), 
	.B1(n7977), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6330));
   INVX1 U3221 (.Y(n7977), 
	.A(\ram[191][6] ));
   OAI22X1 U3222 (.Y(n3643), 
	.B1(n7978), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6332));
   INVX1 U3223 (.Y(n7978), 
	.A(\ram[191][5] ));
   OAI22X1 U3224 (.Y(n3642), 
	.B1(n7979), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6334));
   INVX1 U3225 (.Y(n7979), 
	.A(\ram[191][4] ));
   OAI22X1 U3226 (.Y(n3641), 
	.B1(n7980), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6336));
   INVX1 U3227 (.Y(n7980), 
	.A(\ram[191][3] ));
   OAI22X1 U3228 (.Y(n3640), 
	.B1(n7981), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6338));
   INVX1 U3229 (.Y(n7981), 
	.A(\ram[191][2] ));
   OAI22X1 U3230 (.Y(n3639), 
	.B1(n7982), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6306));
   INVX1 U3231 (.Y(n7982), 
	.A(\ram[191][1] ));
   OAI22X1 U3232 (.Y(n3638), 
	.B1(n7983), 
	.B0(n7967), 
	.A1(n7966), 
	.A0(n6309));
   INVX1 U3233 (.Y(n7983), 
	.A(\ram[191][0] ));
   NOR2BX1 U3234 (.Y(n7967), 
	.B(n7966), 
	.AN(mem_write_en));
   NAND2X1 U3235 (.Y(n7966), 
	.B(n6533), 
	.A(n7984));
   OAI22X1 U3236 (.Y(n3637), 
	.B1(n7987), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6311));
   INVX1 U3237 (.Y(n7987), 
	.A(\ram[190][15] ));
   OAI22X1 U3238 (.Y(n3636), 
	.B1(n7988), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6314));
   INVX1 U3239 (.Y(n7988), 
	.A(\ram[190][14] ));
   OAI22X1 U3240 (.Y(n3635), 
	.B1(n7989), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6316));
   INVX1 U3241 (.Y(n7989), 
	.A(\ram[190][13] ));
   OAI22X1 U3242 (.Y(n3634), 
	.B1(n7990), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6318));
   INVX1 U3243 (.Y(n7990), 
	.A(\ram[190][12] ));
   OAI22X1 U3244 (.Y(n3633), 
	.B1(n7991), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6320));
   INVX1 U3245 (.Y(n7991), 
	.A(\ram[190][11] ));
   OAI22X1 U3246 (.Y(n3632), 
	.B1(n7992), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6322));
   INVX1 U3247 (.Y(n7992), 
	.A(\ram[190][10] ));
   OAI22X1 U3248 (.Y(n3631), 
	.B1(n7993), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6324));
   INVX1 U3249 (.Y(n7993), 
	.A(\ram[190][9] ));
   OAI22X1 U3250 (.Y(n3630), 
	.B1(n7994), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6326));
   INVX1 U3251 (.Y(n7994), 
	.A(\ram[190][8] ));
   OAI22X1 U3252 (.Y(n3629), 
	.B1(n7995), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6328));
   INVX1 U3253 (.Y(n7995), 
	.A(\ram[190][7] ));
   OAI22X1 U3254 (.Y(n3628), 
	.B1(n7996), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6330));
   INVX1 U3255 (.Y(n7996), 
	.A(\ram[190][6] ));
   OAI22X1 U3256 (.Y(n3627), 
	.B1(n7997), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6332));
   INVX1 U3257 (.Y(n7997), 
	.A(\ram[190][5] ));
   OAI22X1 U3258 (.Y(n3626), 
	.B1(n7998), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6334));
   INVX1 U3259 (.Y(n7998), 
	.A(\ram[190][4] ));
   OAI22X1 U3260 (.Y(n3625), 
	.B1(n7999), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6336));
   INVX1 U3261 (.Y(n7999), 
	.A(\ram[190][3] ));
   OAI22X1 U3262 (.Y(n3624), 
	.B1(n8000), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6338));
   INVX1 U3263 (.Y(n8000), 
	.A(\ram[190][2] ));
   OAI22X1 U3264 (.Y(n3623), 
	.B1(n8001), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6306));
   INVX1 U3265 (.Y(n8001), 
	.A(\ram[190][1] ));
   OAI22X1 U3266 (.Y(n3622), 
	.B1(n8002), 
	.B0(n7986), 
	.A1(n7985), 
	.A0(n6309));
   INVX1 U3267 (.Y(n8002), 
	.A(\ram[190][0] ));
   NOR2BX1 U3268 (.Y(n7986), 
	.B(n7985), 
	.AN(mem_write_en));
   NAND2X1 U3269 (.Y(n7985), 
	.B(n6553), 
	.A(n7984));
   OAI22X1 U3270 (.Y(n3621), 
	.B1(n8005), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6311));
   INVX1 U3271 (.Y(n8005), 
	.A(\ram[189][15] ));
   OAI22X1 U3272 (.Y(n3620), 
	.B1(n8006), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6314));
   INVX1 U3273 (.Y(n8006), 
	.A(\ram[189][14] ));
   OAI22X1 U3274 (.Y(n3619), 
	.B1(n8007), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6316));
   INVX1 U3275 (.Y(n8007), 
	.A(\ram[189][13] ));
   OAI22X1 U3276 (.Y(n3618), 
	.B1(n8008), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6318));
   INVX1 U3277 (.Y(n8008), 
	.A(\ram[189][12] ));
   OAI22X1 U3278 (.Y(n3617), 
	.B1(n8009), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6320));
   INVX1 U3279 (.Y(n8009), 
	.A(\ram[189][11] ));
   OAI22X1 U3280 (.Y(n3616), 
	.B1(n8010), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6322));
   INVX1 U3281 (.Y(n8010), 
	.A(\ram[189][10] ));
   OAI22X1 U3282 (.Y(n3615), 
	.B1(n8011), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6324));
   INVX1 U3283 (.Y(n8011), 
	.A(\ram[189][9] ));
   OAI22X1 U3284 (.Y(n3614), 
	.B1(n8012), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6326));
   INVX1 U3285 (.Y(n8012), 
	.A(\ram[189][8] ));
   OAI22X1 U3286 (.Y(n3613), 
	.B1(n8013), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6328));
   INVX1 U3287 (.Y(n8013), 
	.A(\ram[189][7] ));
   OAI22X1 U3288 (.Y(n3612), 
	.B1(n8014), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6330));
   INVX1 U3289 (.Y(n8014), 
	.A(\ram[189][6] ));
   OAI22X1 U3290 (.Y(n3611), 
	.B1(n8015), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6332));
   INVX1 U3291 (.Y(n8015), 
	.A(\ram[189][5] ));
   OAI22X1 U3292 (.Y(n3610), 
	.B1(n8016), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6334));
   INVX1 U3293 (.Y(n8016), 
	.A(\ram[189][4] ));
   OAI22X1 U3294 (.Y(n3609), 
	.B1(n8017), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6336));
   INVX1 U3295 (.Y(n8017), 
	.A(\ram[189][3] ));
   OAI22X1 U3296 (.Y(n3608), 
	.B1(n8018), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6338));
   INVX1 U3297 (.Y(n8018), 
	.A(\ram[189][2] ));
   OAI22X1 U3298 (.Y(n3607), 
	.B1(n8019), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6306));
   INVX1 U3299 (.Y(n8019), 
	.A(\ram[189][1] ));
   OAI22X1 U3300 (.Y(n3606), 
	.B1(n8020), 
	.B0(n8004), 
	.A1(n8003), 
	.A0(n6309));
   INVX1 U3301 (.Y(n8020), 
	.A(\ram[189][0] ));
   NOR2BX1 U3302 (.Y(n8004), 
	.B(n8003), 
	.AN(mem_write_en));
   NAND2X1 U3303 (.Y(n8003), 
	.B(n6572), 
	.A(n7984));
   OAI22X1 U3304 (.Y(n3605), 
	.B1(n8023), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6311));
   INVX1 U3305 (.Y(n8023), 
	.A(\ram[188][15] ));
   OAI22X1 U3306 (.Y(n3604), 
	.B1(n8024), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6314));
   INVX1 U3307 (.Y(n8024), 
	.A(\ram[188][14] ));
   OAI22X1 U3308 (.Y(n3603), 
	.B1(n8025), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6316));
   INVX1 U3309 (.Y(n8025), 
	.A(\ram[188][13] ));
   OAI22X1 U3310 (.Y(n3602), 
	.B1(n8026), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6318));
   INVX1 U3311 (.Y(n8026), 
	.A(\ram[188][12] ));
   OAI22X1 U3312 (.Y(n3601), 
	.B1(n8027), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6320));
   INVX1 U3313 (.Y(n8027), 
	.A(\ram[188][11] ));
   OAI22X1 U3314 (.Y(n3600), 
	.B1(n8028), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6322));
   INVX1 U3315 (.Y(n8028), 
	.A(\ram[188][10] ));
   OAI22X1 U3316 (.Y(n3599), 
	.B1(n8029), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6324));
   INVX1 U3317 (.Y(n8029), 
	.A(\ram[188][9] ));
   OAI22X1 U3318 (.Y(n3598), 
	.B1(n8030), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6326));
   INVX1 U3319 (.Y(n8030), 
	.A(\ram[188][8] ));
   OAI22X1 U3320 (.Y(n3597), 
	.B1(n8031), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6328));
   INVX1 U3321 (.Y(n8031), 
	.A(\ram[188][7] ));
   OAI22X1 U3322 (.Y(n3596), 
	.B1(n8032), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6330));
   INVX1 U3323 (.Y(n8032), 
	.A(\ram[188][6] ));
   OAI22X1 U3324 (.Y(n3595), 
	.B1(n8033), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6332));
   INVX1 U3325 (.Y(n8033), 
	.A(\ram[188][5] ));
   OAI22X1 U3326 (.Y(n3594), 
	.B1(n8034), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6334));
   INVX1 U3327 (.Y(n8034), 
	.A(\ram[188][4] ));
   OAI22X1 U3328 (.Y(n3593), 
	.B1(n8035), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6336));
   INVX1 U3329 (.Y(n8035), 
	.A(\ram[188][3] ));
   OAI22X1 U3330 (.Y(n3592), 
	.B1(n8036), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6338));
   INVX1 U3331 (.Y(n8036), 
	.A(\ram[188][2] ));
   OAI22X1 U3332 (.Y(n3591), 
	.B1(n8037), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6306));
   INVX1 U3333 (.Y(n8037), 
	.A(\ram[188][1] ));
   OAI22X1 U3334 (.Y(n3590), 
	.B1(n8038), 
	.B0(n8022), 
	.A1(n8021), 
	.A0(n6309));
   INVX1 U3335 (.Y(n8038), 
	.A(\ram[188][0] ));
   NOR2BX1 U3336 (.Y(n8022), 
	.B(n8021), 
	.AN(mem_write_en));
   NAND2X1 U3337 (.Y(n8021), 
	.B(n6591), 
	.A(n7984));
   OAI22X1 U3338 (.Y(n3589), 
	.B1(n8041), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6311));
   INVX1 U3339 (.Y(n8041), 
	.A(\ram[187][15] ));
   OAI22X1 U3340 (.Y(n3588), 
	.B1(n8042), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6314));
   INVX1 U3341 (.Y(n8042), 
	.A(\ram[187][14] ));
   OAI22X1 U3342 (.Y(n3587), 
	.B1(n8043), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6316));
   INVX1 U3343 (.Y(n8043), 
	.A(\ram[187][13] ));
   OAI22X1 U3344 (.Y(n3586), 
	.B1(n8044), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6318));
   INVX1 U3345 (.Y(n8044), 
	.A(\ram[187][12] ));
   OAI22X1 U3346 (.Y(n3585), 
	.B1(n8045), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6320));
   INVX1 U3347 (.Y(n8045), 
	.A(\ram[187][11] ));
   OAI22X1 U3348 (.Y(n3584), 
	.B1(n8046), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6322));
   INVX1 U3349 (.Y(n8046), 
	.A(\ram[187][10] ));
   OAI22X1 U3350 (.Y(n3583), 
	.B1(n8047), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6324));
   INVX1 U3351 (.Y(n8047), 
	.A(\ram[187][9] ));
   OAI22X1 U3352 (.Y(n3582), 
	.B1(n8048), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6326));
   INVX1 U3353 (.Y(n8048), 
	.A(\ram[187][8] ));
   OAI22X1 U3354 (.Y(n3581), 
	.B1(n8049), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6328));
   INVX1 U3355 (.Y(n8049), 
	.A(\ram[187][7] ));
   OAI22X1 U3356 (.Y(n3580), 
	.B1(n8050), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6330));
   INVX1 U3357 (.Y(n8050), 
	.A(\ram[187][6] ));
   OAI22X1 U3358 (.Y(n3579), 
	.B1(n8051), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6332));
   INVX1 U3359 (.Y(n8051), 
	.A(\ram[187][5] ));
   OAI22X1 U3360 (.Y(n3578), 
	.B1(n8052), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6334));
   INVX1 U3361 (.Y(n8052), 
	.A(\ram[187][4] ));
   OAI22X1 U3362 (.Y(n3577), 
	.B1(n8053), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6336));
   INVX1 U3363 (.Y(n8053), 
	.A(\ram[187][3] ));
   OAI22X1 U3364 (.Y(n3576), 
	.B1(n8054), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6338));
   INVX1 U3365 (.Y(n8054), 
	.A(\ram[187][2] ));
   OAI22X1 U3366 (.Y(n3575), 
	.B1(n8055), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6306));
   INVX1 U3367 (.Y(n8055), 
	.A(\ram[187][1] ));
   OAI22X1 U3368 (.Y(n3574), 
	.B1(n8056), 
	.B0(n8040), 
	.A1(n8039), 
	.A0(n6309));
   INVX1 U3369 (.Y(n8056), 
	.A(\ram[187][0] ));
   NOR2BX1 U3370 (.Y(n8040), 
	.B(n8039), 
	.AN(mem_write_en));
   NAND2X1 U3371 (.Y(n8039), 
	.B(n6610), 
	.A(n7984));
   OAI22X1 U3372 (.Y(n3573), 
	.B1(n8059), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6311));
   INVX1 U3373 (.Y(n8059), 
	.A(\ram[186][15] ));
   OAI22X1 U3374 (.Y(n3572), 
	.B1(n8060), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6314));
   INVX1 U3375 (.Y(n8060), 
	.A(\ram[186][14] ));
   OAI22X1 U3376 (.Y(n3571), 
	.B1(n8061), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6316));
   INVX1 U3377 (.Y(n8061), 
	.A(\ram[186][13] ));
   OAI22X1 U3378 (.Y(n3570), 
	.B1(n8062), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6318));
   INVX1 U3379 (.Y(n8062), 
	.A(\ram[186][12] ));
   OAI22X1 U3380 (.Y(n3569), 
	.B1(n8063), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6320));
   INVX1 U3381 (.Y(n8063), 
	.A(\ram[186][11] ));
   OAI22X1 U3382 (.Y(n3568), 
	.B1(n8064), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6322));
   INVX1 U3383 (.Y(n8064), 
	.A(\ram[186][10] ));
   OAI22X1 U3384 (.Y(n3567), 
	.B1(n8065), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6324));
   INVX1 U3385 (.Y(n8065), 
	.A(\ram[186][9] ));
   OAI22X1 U3386 (.Y(n3566), 
	.B1(n8066), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6326));
   INVX1 U3387 (.Y(n8066), 
	.A(\ram[186][8] ));
   OAI22X1 U3388 (.Y(n3565), 
	.B1(n8067), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6328));
   INVX1 U3389 (.Y(n8067), 
	.A(\ram[186][7] ));
   OAI22X1 U3390 (.Y(n3564), 
	.B1(n8068), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6330));
   INVX1 U3391 (.Y(n8068), 
	.A(\ram[186][6] ));
   OAI22X1 U3392 (.Y(n3563), 
	.B1(n8069), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6332));
   INVX1 U3393 (.Y(n8069), 
	.A(\ram[186][5] ));
   OAI22X1 U3394 (.Y(n3562), 
	.B1(n8070), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6334));
   INVX1 U3395 (.Y(n8070), 
	.A(\ram[186][4] ));
   OAI22X1 U3396 (.Y(n3561), 
	.B1(n8071), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6336));
   INVX1 U3397 (.Y(n8071), 
	.A(\ram[186][3] ));
   OAI22X1 U3398 (.Y(n3560), 
	.B1(n8072), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6338));
   INVX1 U3399 (.Y(n8072), 
	.A(\ram[186][2] ));
   OAI22X1 U3400 (.Y(n3559), 
	.B1(n8073), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6306));
   INVX1 U3401 (.Y(n8073), 
	.A(\ram[186][1] ));
   OAI22X1 U3402 (.Y(n3558), 
	.B1(n8074), 
	.B0(n8058), 
	.A1(n8057), 
	.A0(n6309));
   INVX1 U3403 (.Y(n8074), 
	.A(\ram[186][0] ));
   NOR2BX1 U3404 (.Y(n8058), 
	.B(n8057), 
	.AN(mem_write_en));
   NAND2X1 U3405 (.Y(n8057), 
	.B(n6629), 
	.A(n7984));
   OAI22X1 U3406 (.Y(n3557), 
	.B1(n8077), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6311));
   INVX1 U3407 (.Y(n8077), 
	.A(\ram[185][15] ));
   OAI22X1 U3408 (.Y(n3556), 
	.B1(n8078), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6314));
   INVX1 U3409 (.Y(n8078), 
	.A(\ram[185][14] ));
   OAI22X1 U3410 (.Y(n3555), 
	.B1(n8079), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6316));
   INVX1 U3411 (.Y(n8079), 
	.A(\ram[185][13] ));
   OAI22X1 U3412 (.Y(n3554), 
	.B1(n8080), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6318));
   INVX1 U3413 (.Y(n8080), 
	.A(\ram[185][12] ));
   OAI22X1 U3414 (.Y(n3553), 
	.B1(n8081), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6320));
   INVX1 U3415 (.Y(n8081), 
	.A(\ram[185][11] ));
   OAI22X1 U3416 (.Y(n3552), 
	.B1(n8082), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6322));
   INVX1 U3417 (.Y(n8082), 
	.A(\ram[185][10] ));
   OAI22X1 U3418 (.Y(n3551), 
	.B1(n8083), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6324));
   INVX1 U3419 (.Y(n8083), 
	.A(\ram[185][9] ));
   OAI22X1 U3420 (.Y(n3550), 
	.B1(n8084), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6326));
   INVX1 U3421 (.Y(n8084), 
	.A(\ram[185][8] ));
   OAI22X1 U3422 (.Y(n3549), 
	.B1(n8085), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6328));
   INVX1 U3423 (.Y(n8085), 
	.A(\ram[185][7] ));
   OAI22X1 U3424 (.Y(n3548), 
	.B1(n8086), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6330));
   INVX1 U3425 (.Y(n8086), 
	.A(\ram[185][6] ));
   OAI22X1 U3426 (.Y(n3547), 
	.B1(n8087), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6332));
   INVX1 U3427 (.Y(n8087), 
	.A(\ram[185][5] ));
   OAI22X1 U3428 (.Y(n3546), 
	.B1(n8088), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6334));
   INVX1 U3429 (.Y(n8088), 
	.A(\ram[185][4] ));
   OAI22X1 U3430 (.Y(n3545), 
	.B1(n8089), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6336));
   INVX1 U3431 (.Y(n8089), 
	.A(\ram[185][3] ));
   OAI22X1 U3432 (.Y(n3544), 
	.B1(n8090), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6338));
   INVX1 U3433 (.Y(n8090), 
	.A(\ram[185][2] ));
   OAI22X1 U3434 (.Y(n3543), 
	.B1(n8091), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6306));
   INVX1 U3435 (.Y(n8091), 
	.A(\ram[185][1] ));
   OAI22X1 U3436 (.Y(n3542), 
	.B1(n8092), 
	.B0(n8076), 
	.A1(n8075), 
	.A0(n6309));
   INVX1 U3437 (.Y(n8092), 
	.A(\ram[185][0] ));
   NOR2BX1 U3438 (.Y(n8076), 
	.B(n8075), 
	.AN(mem_write_en));
   NAND2X1 U3439 (.Y(n8075), 
	.B(n6342), 
	.A(n7984));
   OAI22X1 U3440 (.Y(n3541), 
	.B1(n8095), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6311));
   INVX1 U3441 (.Y(n8095), 
	.A(\ram[184][15] ));
   OAI22X1 U3442 (.Y(n3540), 
	.B1(n8096), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6314));
   INVX1 U3443 (.Y(n8096), 
	.A(\ram[184][14] ));
   OAI22X1 U3444 (.Y(n3539), 
	.B1(n8097), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6316));
   INVX1 U3445 (.Y(n8097), 
	.A(\ram[184][13] ));
   OAI22X1 U3446 (.Y(n3538), 
	.B1(n8098), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6318));
   INVX1 U3447 (.Y(n8098), 
	.A(\ram[184][12] ));
   OAI22X1 U3448 (.Y(n3537), 
	.B1(n8099), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6320));
   INVX1 U3449 (.Y(n8099), 
	.A(\ram[184][11] ));
   OAI22X1 U3450 (.Y(n3536), 
	.B1(n8100), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6322));
   INVX1 U3451 (.Y(n8100), 
	.A(\ram[184][10] ));
   OAI22X1 U3452 (.Y(n3535), 
	.B1(n8101), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6324));
   INVX1 U3453 (.Y(n8101), 
	.A(\ram[184][9] ));
   OAI22X1 U3454 (.Y(n3534), 
	.B1(n8102), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6326));
   INVX1 U3455 (.Y(n8102), 
	.A(\ram[184][8] ));
   OAI22X1 U3456 (.Y(n3533), 
	.B1(n8103), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6328));
   INVX1 U3457 (.Y(n8103), 
	.A(\ram[184][7] ));
   OAI22X1 U3458 (.Y(n3532), 
	.B1(n8104), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6330));
   INVX1 U3459 (.Y(n8104), 
	.A(\ram[184][6] ));
   OAI22X1 U3460 (.Y(n3531), 
	.B1(n8105), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6332));
   INVX1 U3461 (.Y(n8105), 
	.A(\ram[184][5] ));
   OAI22X1 U3462 (.Y(n3530), 
	.B1(n8106), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6334));
   INVX1 U3463 (.Y(n8106), 
	.A(\ram[184][4] ));
   OAI22X1 U3464 (.Y(n3529), 
	.B1(n8107), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6336));
   INVX1 U3465 (.Y(n8107), 
	.A(\ram[184][3] ));
   OAI22X1 U3466 (.Y(n3528), 
	.B1(n8108), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6338));
   INVX1 U3467 (.Y(n8108), 
	.A(\ram[184][2] ));
   OAI22X1 U3468 (.Y(n3527), 
	.B1(n8109), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6306));
   INVX1 U3469 (.Y(n8109), 
	.A(\ram[184][1] ));
   OAI22X1 U3470 (.Y(n3526), 
	.B1(n8110), 
	.B0(n8094), 
	.A1(n8093), 
	.A0(n6309));
   INVX1 U3471 (.Y(n8110), 
	.A(\ram[184][0] ));
   NOR2BX1 U3472 (.Y(n8094), 
	.B(n8093), 
	.AN(mem_write_en));
   NAND2X1 U3473 (.Y(n8093), 
	.B(n6362), 
	.A(n7984));
   OAI22X1 U3474 (.Y(n3525), 
	.B1(n8113), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6311));
   INVX1 U3475 (.Y(n8113), 
	.A(\ram[183][15] ));
   OAI22X1 U3476 (.Y(n3524), 
	.B1(n8114), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6314));
   INVX1 U3477 (.Y(n8114), 
	.A(\ram[183][14] ));
   OAI22X1 U3478 (.Y(n3523), 
	.B1(n8115), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6316));
   INVX1 U3479 (.Y(n8115), 
	.A(\ram[183][13] ));
   OAI22X1 U3480 (.Y(n3522), 
	.B1(n8116), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6318));
   INVX1 U3481 (.Y(n8116), 
	.A(\ram[183][12] ));
   OAI22X1 U3482 (.Y(n3521), 
	.B1(n8117), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6320));
   INVX1 U3483 (.Y(n8117), 
	.A(\ram[183][11] ));
   OAI22X1 U3484 (.Y(n3520), 
	.B1(n8118), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6322));
   INVX1 U3485 (.Y(n8118), 
	.A(\ram[183][10] ));
   OAI22X1 U3486 (.Y(n3519), 
	.B1(n8119), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6324));
   INVX1 U3487 (.Y(n8119), 
	.A(\ram[183][9] ));
   OAI22X1 U3488 (.Y(n3518), 
	.B1(n8120), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6326));
   INVX1 U3489 (.Y(n8120), 
	.A(\ram[183][8] ));
   OAI22X1 U3490 (.Y(n3517), 
	.B1(n8121), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6328));
   INVX1 U3491 (.Y(n8121), 
	.A(\ram[183][7] ));
   OAI22X1 U3492 (.Y(n3516), 
	.B1(n8122), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6330));
   INVX1 U3493 (.Y(n8122), 
	.A(\ram[183][6] ));
   OAI22X1 U3494 (.Y(n3515), 
	.B1(n8123), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6332));
   INVX1 U3495 (.Y(n8123), 
	.A(\ram[183][5] ));
   OAI22X1 U3496 (.Y(n3514), 
	.B1(n8124), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6334));
   INVX1 U3497 (.Y(n8124), 
	.A(\ram[183][4] ));
   OAI22X1 U3498 (.Y(n3513), 
	.B1(n8125), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6336));
   INVX1 U3499 (.Y(n8125), 
	.A(\ram[183][3] ));
   OAI22X1 U3500 (.Y(n3512), 
	.B1(n8126), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6338));
   INVX1 U3501 (.Y(n8126), 
	.A(\ram[183][2] ));
   OAI22X1 U3502 (.Y(n3511), 
	.B1(n8127), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6306));
   INVX1 U3503 (.Y(n8127), 
	.A(\ram[183][1] ));
   OAI22X1 U3504 (.Y(n3510), 
	.B1(n8128), 
	.B0(n8112), 
	.A1(n8111), 
	.A0(n6309));
   INVX1 U3505 (.Y(n8128), 
	.A(\ram[183][0] ));
   NOR2BX1 U3506 (.Y(n8112), 
	.B(n8111), 
	.AN(mem_write_en));
   NAND2X1 U3507 (.Y(n8111), 
	.B(n6381), 
	.A(n7984));
   OAI22X1 U3508 (.Y(n3509), 
	.B1(n8131), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6311));
   INVX1 U3509 (.Y(n8131), 
	.A(\ram[182][15] ));
   OAI22X1 U3510 (.Y(n3508), 
	.B1(n8132), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6314));
   INVX1 U3511 (.Y(n8132), 
	.A(\ram[182][14] ));
   OAI22X1 U3512 (.Y(n3507), 
	.B1(n8133), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6316));
   INVX1 U3513 (.Y(n8133), 
	.A(\ram[182][13] ));
   OAI22X1 U3514 (.Y(n3506), 
	.B1(n8134), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6318));
   INVX1 U3515 (.Y(n8134), 
	.A(\ram[182][12] ));
   OAI22X1 U3516 (.Y(n3505), 
	.B1(n8135), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6320));
   INVX1 U3517 (.Y(n8135), 
	.A(\ram[182][11] ));
   OAI22X1 U3518 (.Y(n3504), 
	.B1(n8136), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6322));
   INVX1 U3519 (.Y(n8136), 
	.A(\ram[182][10] ));
   OAI22X1 U3520 (.Y(n3503), 
	.B1(n8137), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6324));
   INVX1 U3521 (.Y(n8137), 
	.A(\ram[182][9] ));
   OAI22X1 U3522 (.Y(n3502), 
	.B1(n8138), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6326));
   INVX1 U3523 (.Y(n8138), 
	.A(\ram[182][8] ));
   OAI22X1 U3524 (.Y(n3501), 
	.B1(n8139), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6328));
   INVX1 U3525 (.Y(n8139), 
	.A(\ram[182][7] ));
   OAI22X1 U3526 (.Y(n3500), 
	.B1(n8140), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6330));
   INVX1 U3527 (.Y(n8140), 
	.A(\ram[182][6] ));
   OAI22X1 U3528 (.Y(n3499), 
	.B1(n8141), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6332));
   INVX1 U3529 (.Y(n8141), 
	.A(\ram[182][5] ));
   OAI22X1 U3530 (.Y(n3498), 
	.B1(n8142), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6334));
   INVX1 U3531 (.Y(n8142), 
	.A(\ram[182][4] ));
   OAI22X1 U3532 (.Y(n3497), 
	.B1(n8143), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6336));
   INVX1 U3533 (.Y(n8143), 
	.A(\ram[182][3] ));
   OAI22X1 U3534 (.Y(n3496), 
	.B1(n8144), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6338));
   INVX1 U3535 (.Y(n8144), 
	.A(\ram[182][2] ));
   OAI22X1 U3536 (.Y(n3495), 
	.B1(n8145), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6306));
   INVX1 U3537 (.Y(n8145), 
	.A(\ram[182][1] ));
   OAI22X1 U3538 (.Y(n3494), 
	.B1(n8146), 
	.B0(n8130), 
	.A1(n8129), 
	.A0(n6309));
   INVX1 U3539 (.Y(n8146), 
	.A(\ram[182][0] ));
   NOR2BX1 U3540 (.Y(n8130), 
	.B(n8129), 
	.AN(mem_write_en));
   NAND2X1 U3541 (.Y(n8129), 
	.B(n6400), 
	.A(n7984));
   OAI22X1 U3542 (.Y(n3493), 
	.B1(n8149), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6311));
   INVX1 U3543 (.Y(n8149), 
	.A(\ram[181][15] ));
   OAI22X1 U3544 (.Y(n3492), 
	.B1(n8150), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6314));
   INVX1 U3545 (.Y(n8150), 
	.A(\ram[181][14] ));
   OAI22X1 U3546 (.Y(n3491), 
	.B1(n8151), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6316));
   INVX1 U3547 (.Y(n8151), 
	.A(\ram[181][13] ));
   OAI22X1 U3548 (.Y(n3490), 
	.B1(n8152), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6318));
   INVX1 U3549 (.Y(n8152), 
	.A(\ram[181][12] ));
   OAI22X1 U3550 (.Y(n3489), 
	.B1(n8153), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6320));
   INVX1 U3551 (.Y(n8153), 
	.A(\ram[181][11] ));
   OAI22X1 U3552 (.Y(n3488), 
	.B1(n8154), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6322));
   INVX1 U3553 (.Y(n8154), 
	.A(\ram[181][10] ));
   OAI22X1 U3554 (.Y(n3487), 
	.B1(n8155), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6324));
   INVX1 U3555 (.Y(n8155), 
	.A(\ram[181][9] ));
   OAI22X1 U3556 (.Y(n3486), 
	.B1(n8156), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6326));
   INVX1 U3557 (.Y(n8156), 
	.A(\ram[181][8] ));
   OAI22X1 U3558 (.Y(n3485), 
	.B1(n8157), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6328));
   INVX1 U3559 (.Y(n8157), 
	.A(\ram[181][7] ));
   OAI22X1 U3560 (.Y(n3484), 
	.B1(n8158), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6330));
   INVX1 U3561 (.Y(n8158), 
	.A(\ram[181][6] ));
   OAI22X1 U3562 (.Y(n3483), 
	.B1(n8159), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6332));
   INVX1 U3563 (.Y(n8159), 
	.A(\ram[181][5] ));
   OAI22X1 U3564 (.Y(n3482), 
	.B1(n8160), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6334));
   INVX1 U3565 (.Y(n8160), 
	.A(\ram[181][4] ));
   OAI22X1 U3566 (.Y(n3481), 
	.B1(n8161), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6336));
   INVX1 U3567 (.Y(n8161), 
	.A(\ram[181][3] ));
   OAI22X1 U3568 (.Y(n3480), 
	.B1(n8162), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6338));
   INVX1 U3569 (.Y(n8162), 
	.A(\ram[181][2] ));
   OAI22X1 U3570 (.Y(n3479), 
	.B1(n8163), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6306));
   INVX1 U3571 (.Y(n8163), 
	.A(\ram[181][1] ));
   OAI22X1 U3572 (.Y(n3478), 
	.B1(n8164), 
	.B0(n8148), 
	.A1(n8147), 
	.A0(n6309));
   INVX1 U3573 (.Y(n8164), 
	.A(\ram[181][0] ));
   NOR2BX1 U3574 (.Y(n8148), 
	.B(n8147), 
	.AN(mem_write_en));
   NAND2X1 U3575 (.Y(n8147), 
	.B(n6419), 
	.A(n7984));
   OAI22X1 U3576 (.Y(n3477), 
	.B1(n8167), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6311));
   INVX1 U3577 (.Y(n8167), 
	.A(\ram[180][15] ));
   OAI22X1 U3578 (.Y(n3476), 
	.B1(n8168), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6314));
   INVX1 U3579 (.Y(n8168), 
	.A(\ram[180][14] ));
   OAI22X1 U3580 (.Y(n3475), 
	.B1(n8169), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6316));
   INVX1 U3581 (.Y(n8169), 
	.A(\ram[180][13] ));
   OAI22X1 U3582 (.Y(n3474), 
	.B1(n8170), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6318));
   INVX1 U3583 (.Y(n8170), 
	.A(\ram[180][12] ));
   OAI22X1 U3584 (.Y(n3473), 
	.B1(n8171), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6320));
   INVX1 U3585 (.Y(n8171), 
	.A(\ram[180][11] ));
   OAI22X1 U3586 (.Y(n3472), 
	.B1(n8172), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6322));
   INVX1 U3587 (.Y(n8172), 
	.A(\ram[180][10] ));
   OAI22X1 U3588 (.Y(n3471), 
	.B1(n8173), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6324));
   INVX1 U3589 (.Y(n8173), 
	.A(\ram[180][9] ));
   OAI22X1 U3590 (.Y(n3470), 
	.B1(n8174), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6326));
   INVX1 U3591 (.Y(n8174), 
	.A(\ram[180][8] ));
   OAI22X1 U3592 (.Y(n3469), 
	.B1(n8175), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6328));
   INVX1 U3593 (.Y(n8175), 
	.A(\ram[180][7] ));
   OAI22X1 U3594 (.Y(n3468), 
	.B1(n8176), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6330));
   INVX1 U3595 (.Y(n8176), 
	.A(\ram[180][6] ));
   OAI22X1 U3596 (.Y(n3467), 
	.B1(n8177), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6332));
   INVX1 U3597 (.Y(n8177), 
	.A(\ram[180][5] ));
   OAI22X1 U3598 (.Y(n3466), 
	.B1(n8178), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6334));
   INVX1 U3599 (.Y(n8178), 
	.A(\ram[180][4] ));
   OAI22X1 U3600 (.Y(n3465), 
	.B1(n8179), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6336));
   INVX1 U3601 (.Y(n8179), 
	.A(\ram[180][3] ));
   OAI22X1 U3602 (.Y(n3464), 
	.B1(n8180), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6338));
   INVX1 U3603 (.Y(n8180), 
	.A(\ram[180][2] ));
   OAI22X1 U3604 (.Y(n3463), 
	.B1(n8181), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6306));
   INVX1 U3605 (.Y(n8181), 
	.A(\ram[180][1] ));
   OAI22X1 U3606 (.Y(n3462), 
	.B1(n8182), 
	.B0(n8166), 
	.A1(n8165), 
	.A0(n6309));
   INVX1 U3607 (.Y(n8182), 
	.A(\ram[180][0] ));
   NOR2BX1 U3608 (.Y(n8166), 
	.B(n8165), 
	.AN(mem_write_en));
   NAND2X1 U3609 (.Y(n8165), 
	.B(n6438), 
	.A(n7984));
   OAI22X1 U3610 (.Y(n3461), 
	.B1(n8185), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6311));
   INVX1 U3611 (.Y(n8185), 
	.A(\ram[179][15] ));
   OAI22X1 U3612 (.Y(n3460), 
	.B1(n8186), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6314));
   INVX1 U3613 (.Y(n8186), 
	.A(\ram[179][14] ));
   OAI22X1 U3614 (.Y(n3459), 
	.B1(n8187), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6316));
   INVX1 U3615 (.Y(n8187), 
	.A(\ram[179][13] ));
   OAI22X1 U3616 (.Y(n3458), 
	.B1(n8188), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6318));
   INVX1 U3617 (.Y(n8188), 
	.A(\ram[179][12] ));
   OAI22X1 U3618 (.Y(n3457), 
	.B1(n8189), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6320));
   INVX1 U3619 (.Y(n8189), 
	.A(\ram[179][11] ));
   OAI22X1 U3620 (.Y(n3456), 
	.B1(n8190), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6322));
   INVX1 U3621 (.Y(n8190), 
	.A(\ram[179][10] ));
   OAI22X1 U3622 (.Y(n3455), 
	.B1(n8191), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6324));
   INVX1 U3623 (.Y(n8191), 
	.A(\ram[179][9] ));
   OAI22X1 U3624 (.Y(n3454), 
	.B1(n8192), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6326));
   INVX1 U3625 (.Y(n8192), 
	.A(\ram[179][8] ));
   OAI22X1 U3626 (.Y(n3453), 
	.B1(n8193), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6328));
   INVX1 U3627 (.Y(n8193), 
	.A(\ram[179][7] ));
   OAI22X1 U3628 (.Y(n3452), 
	.B1(n8194), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6330));
   INVX1 U3629 (.Y(n8194), 
	.A(\ram[179][6] ));
   OAI22X1 U3630 (.Y(n3451), 
	.B1(n8195), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6332));
   INVX1 U3631 (.Y(n8195), 
	.A(\ram[179][5] ));
   OAI22X1 U3632 (.Y(n3450), 
	.B1(n8196), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6334));
   INVX1 U3633 (.Y(n8196), 
	.A(\ram[179][4] ));
   OAI22X1 U3634 (.Y(n3449), 
	.B1(n8197), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6336));
   INVX1 U3635 (.Y(n8197), 
	.A(\ram[179][3] ));
   OAI22X1 U3636 (.Y(n3448), 
	.B1(n8198), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6338));
   INVX1 U3637 (.Y(n8198), 
	.A(\ram[179][2] ));
   OAI22X1 U3638 (.Y(n3447), 
	.B1(n8199), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6306));
   INVX1 U3639 (.Y(n8199), 
	.A(\ram[179][1] ));
   OAI22X1 U3640 (.Y(n3446), 
	.B1(n8200), 
	.B0(n8184), 
	.A1(n8183), 
	.A0(n6309));
   INVX1 U3641 (.Y(n8200), 
	.A(\ram[179][0] ));
   NOR2BX1 U3642 (.Y(n8184), 
	.B(n8183), 
	.AN(mem_write_en));
   NAND2X1 U3643 (.Y(n8183), 
	.B(n6457), 
	.A(n7984));
   OAI22X1 U3644 (.Y(n3445), 
	.B1(n8203), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6311));
   INVX1 U3645 (.Y(n8203), 
	.A(\ram[178][15] ));
   OAI22X1 U3646 (.Y(n3444), 
	.B1(n8204), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6314));
   INVX1 U3647 (.Y(n8204), 
	.A(\ram[178][14] ));
   OAI22X1 U3648 (.Y(n3443), 
	.B1(n8205), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6316));
   INVX1 U3649 (.Y(n8205), 
	.A(\ram[178][13] ));
   OAI22X1 U3650 (.Y(n3442), 
	.B1(n8206), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6318));
   INVX1 U3651 (.Y(n8206), 
	.A(\ram[178][12] ));
   OAI22X1 U3652 (.Y(n3441), 
	.B1(n8207), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6320));
   INVX1 U3653 (.Y(n8207), 
	.A(\ram[178][11] ));
   OAI22X1 U3654 (.Y(n3440), 
	.B1(n8208), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6322));
   INVX1 U3655 (.Y(n8208), 
	.A(\ram[178][10] ));
   OAI22X1 U3656 (.Y(n3439), 
	.B1(n8209), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6324));
   INVX1 U3657 (.Y(n8209), 
	.A(\ram[178][9] ));
   OAI22X1 U3658 (.Y(n3438), 
	.B1(n8210), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6326));
   INVX1 U3659 (.Y(n8210), 
	.A(\ram[178][8] ));
   OAI22X1 U3660 (.Y(n3437), 
	.B1(n8211), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6328));
   INVX1 U3661 (.Y(n8211), 
	.A(\ram[178][7] ));
   OAI22X1 U3662 (.Y(n3436), 
	.B1(n8212), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6330));
   INVX1 U3663 (.Y(n8212), 
	.A(\ram[178][6] ));
   OAI22X1 U3664 (.Y(n3435), 
	.B1(n8213), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6332));
   INVX1 U3665 (.Y(n8213), 
	.A(\ram[178][5] ));
   OAI22X1 U3666 (.Y(n3434), 
	.B1(n8214), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6334));
   INVX1 U3667 (.Y(n8214), 
	.A(\ram[178][4] ));
   OAI22X1 U3668 (.Y(n3433), 
	.B1(n8215), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6336));
   INVX1 U3669 (.Y(n8215), 
	.A(\ram[178][3] ));
   OAI22X1 U3670 (.Y(n3432), 
	.B1(n8216), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6338));
   INVX1 U3671 (.Y(n8216), 
	.A(\ram[178][2] ));
   OAI22X1 U3672 (.Y(n3431), 
	.B1(n8217), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6306));
   INVX1 U3673 (.Y(n8217), 
	.A(\ram[178][1] ));
   OAI22X1 U3674 (.Y(n3430), 
	.B1(n8218), 
	.B0(n8202), 
	.A1(n8201), 
	.A0(n6309));
   INVX1 U3675 (.Y(n8218), 
	.A(\ram[178][0] ));
   NOR2BX1 U3676 (.Y(n8202), 
	.B(n8201), 
	.AN(mem_write_en));
   NAND2X1 U3677 (.Y(n8201), 
	.B(n6476), 
	.A(n7984));
   OAI22X1 U3678 (.Y(n3429), 
	.B1(n8221), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6311));
   INVX1 U3679 (.Y(n8221), 
	.A(\ram[177][15] ));
   OAI22X1 U3680 (.Y(n3428), 
	.B1(n8222), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6314));
   INVX1 U3681 (.Y(n8222), 
	.A(\ram[177][14] ));
   OAI22X1 U3682 (.Y(n3427), 
	.B1(n8223), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6316));
   INVX1 U3683 (.Y(n8223), 
	.A(\ram[177][13] ));
   OAI22X1 U3684 (.Y(n3426), 
	.B1(n8224), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6318));
   INVX1 U3685 (.Y(n8224), 
	.A(\ram[177][12] ));
   OAI22X1 U3686 (.Y(n3425), 
	.B1(n8225), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6320));
   INVX1 U3687 (.Y(n8225), 
	.A(\ram[177][11] ));
   OAI22X1 U3688 (.Y(n3424), 
	.B1(n8226), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6322));
   INVX1 U3689 (.Y(n8226), 
	.A(\ram[177][10] ));
   OAI22X1 U3690 (.Y(n3423), 
	.B1(n8227), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6324));
   INVX1 U3691 (.Y(n8227), 
	.A(\ram[177][9] ));
   OAI22X1 U3692 (.Y(n3422), 
	.B1(n8228), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6326));
   INVX1 U3693 (.Y(n8228), 
	.A(\ram[177][8] ));
   OAI22X1 U3694 (.Y(n3421), 
	.B1(n8229), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6328));
   INVX1 U3695 (.Y(n8229), 
	.A(\ram[177][7] ));
   OAI22X1 U3696 (.Y(n3420), 
	.B1(n8230), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6330));
   INVX1 U3697 (.Y(n8230), 
	.A(\ram[177][6] ));
   OAI22X1 U3698 (.Y(n3419), 
	.B1(n8231), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6332));
   INVX1 U3699 (.Y(n8231), 
	.A(\ram[177][5] ));
   OAI22X1 U3700 (.Y(n3418), 
	.B1(n8232), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6334));
   INVX1 U3701 (.Y(n8232), 
	.A(\ram[177][4] ));
   OAI22X1 U3702 (.Y(n3417), 
	.B1(n8233), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6336));
   INVX1 U3703 (.Y(n8233), 
	.A(\ram[177][3] ));
   OAI22X1 U3704 (.Y(n3416), 
	.B1(n8234), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6338));
   INVX1 U3705 (.Y(n8234), 
	.A(\ram[177][2] ));
   OAI22X1 U3706 (.Y(n3415), 
	.B1(n8235), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6306));
   INVX1 U3707 (.Y(n8235), 
	.A(\ram[177][1] ));
   OAI22X1 U3708 (.Y(n3414), 
	.B1(n8236), 
	.B0(n8220), 
	.A1(n8219), 
	.A0(n6309));
   INVX1 U3709 (.Y(n8236), 
	.A(\ram[177][0] ));
   NOR2BX1 U3710 (.Y(n8220), 
	.B(n8219), 
	.AN(mem_write_en));
   NAND2X1 U3711 (.Y(n8219), 
	.B(n6495), 
	.A(n7984));
   OAI22X1 U3712 (.Y(n3413), 
	.B1(n8239), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6311));
   INVX1 U3713 (.Y(n8239), 
	.A(\ram[176][15] ));
   OAI22X1 U3714 (.Y(n3412), 
	.B1(n8240), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6314));
   INVX1 U3715 (.Y(n8240), 
	.A(\ram[176][14] ));
   OAI22X1 U3716 (.Y(n3411), 
	.B1(n8241), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6316));
   INVX1 U3717 (.Y(n8241), 
	.A(\ram[176][13] ));
   OAI22X1 U3718 (.Y(n3410), 
	.B1(n8242), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6318));
   INVX1 U3719 (.Y(n8242), 
	.A(\ram[176][12] ));
   OAI22X1 U3720 (.Y(n3409), 
	.B1(n8243), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6320));
   INVX1 U3721 (.Y(n8243), 
	.A(\ram[176][11] ));
   OAI22X1 U3722 (.Y(n3408), 
	.B1(n8244), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6322));
   INVX1 U3723 (.Y(n8244), 
	.A(\ram[176][10] ));
   OAI22X1 U3724 (.Y(n3407), 
	.B1(n8245), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6324));
   INVX1 U3725 (.Y(n8245), 
	.A(\ram[176][9] ));
   OAI22X1 U3726 (.Y(n3406), 
	.B1(n8246), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6326));
   INVX1 U3727 (.Y(n8246), 
	.A(\ram[176][8] ));
   OAI22X1 U3728 (.Y(n3405), 
	.B1(n8247), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6328));
   INVX1 U3729 (.Y(n8247), 
	.A(\ram[176][7] ));
   OAI22X1 U3730 (.Y(n3404), 
	.B1(n8248), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6330));
   INVX1 U3731 (.Y(n8248), 
	.A(\ram[176][6] ));
   OAI22X1 U3732 (.Y(n3403), 
	.B1(n8249), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6332));
   INVX1 U3733 (.Y(n8249), 
	.A(\ram[176][5] ));
   OAI22X1 U3734 (.Y(n3402), 
	.B1(n8250), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6334));
   INVX1 U3735 (.Y(n8250), 
	.A(\ram[176][4] ));
   OAI22X1 U3736 (.Y(n3401), 
	.B1(n8251), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6336));
   INVX1 U3737 (.Y(n8251), 
	.A(\ram[176][3] ));
   OAI22X1 U3738 (.Y(n3400), 
	.B1(n8252), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6338));
   INVX1 U3739 (.Y(n8252), 
	.A(\ram[176][2] ));
   OAI22X1 U3740 (.Y(n3399), 
	.B1(n8253), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6306));
   INVX1 U3741 (.Y(n8253), 
	.A(\ram[176][1] ));
   OAI22X1 U3742 (.Y(n3398), 
	.B1(n8254), 
	.B0(n8238), 
	.A1(n8237), 
	.A0(n6309));
   INVX1 U3743 (.Y(n8254), 
	.A(\ram[176][0] ));
   NOR2BX1 U3744 (.Y(n8238), 
	.B(n8237), 
	.AN(mem_write_en));
   NAND2X1 U3745 (.Y(n8237), 
	.B(n6514), 
	.A(n7984));
   OAI22X1 U3746 (.Y(n3397), 
	.B1(n8257), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6311));
   INVX1 U3747 (.Y(n8257), 
	.A(\ram[175][15] ));
   OAI22X1 U3748 (.Y(n3396), 
	.B1(n8258), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6314));
   INVX1 U3749 (.Y(n8258), 
	.A(\ram[175][14] ));
   OAI22X1 U3750 (.Y(n3395), 
	.B1(n8259), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6316));
   INVX1 U3751 (.Y(n8259), 
	.A(\ram[175][13] ));
   OAI22X1 U3752 (.Y(n3394), 
	.B1(n8260), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6318));
   INVX1 U3753 (.Y(n8260), 
	.A(\ram[175][12] ));
   OAI22X1 U3754 (.Y(n3393), 
	.B1(n8261), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6320));
   INVX1 U3755 (.Y(n8261), 
	.A(\ram[175][11] ));
   OAI22X1 U3756 (.Y(n3392), 
	.B1(n8262), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6322));
   INVX1 U3757 (.Y(n8262), 
	.A(\ram[175][10] ));
   OAI22X1 U3758 (.Y(n3391), 
	.B1(n8263), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6324));
   INVX1 U3759 (.Y(n8263), 
	.A(\ram[175][9] ));
   OAI22X1 U3760 (.Y(n3390), 
	.B1(n8264), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6326));
   INVX1 U3761 (.Y(n8264), 
	.A(\ram[175][8] ));
   OAI22X1 U3762 (.Y(n3389), 
	.B1(n8265), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6328));
   INVX1 U3763 (.Y(n8265), 
	.A(\ram[175][7] ));
   OAI22X1 U3764 (.Y(n3388), 
	.B1(n8266), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6330));
   INVX1 U3765 (.Y(n8266), 
	.A(\ram[175][6] ));
   OAI22X1 U3766 (.Y(n3387), 
	.B1(n8267), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6332));
   INVX1 U3767 (.Y(n8267), 
	.A(\ram[175][5] ));
   OAI22X1 U3768 (.Y(n3386), 
	.B1(n8268), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6334));
   INVX1 U3769 (.Y(n8268), 
	.A(\ram[175][4] ));
   OAI22X1 U3770 (.Y(n3385), 
	.B1(n8269), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6336));
   INVX1 U3771 (.Y(n8269), 
	.A(\ram[175][3] ));
   OAI22X1 U3772 (.Y(n3384), 
	.B1(n8270), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6338));
   INVX1 U3773 (.Y(n8270), 
	.A(\ram[175][2] ));
   OAI22X1 U3774 (.Y(n3383), 
	.B1(n8271), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6306));
   INVX1 U3775 (.Y(n8271), 
	.A(\ram[175][1] ));
   OAI22X1 U3776 (.Y(n3382), 
	.B1(n8272), 
	.B0(n8256), 
	.A1(n8255), 
	.A0(n6309));
   INVX1 U3777 (.Y(n8272), 
	.A(\ram[175][0] ));
   NOR2BX1 U3778 (.Y(n8256), 
	.B(n8255), 
	.AN(mem_write_en));
   NAND2X1 U3779 (.Y(n8255), 
	.B(n6533), 
	.A(n8273));
   OAI22X1 U3780 (.Y(n3381), 
	.B1(n8276), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6311));
   INVX1 U3781 (.Y(n8276), 
	.A(\ram[174][15] ));
   OAI22X1 U3782 (.Y(n3380), 
	.B1(n8277), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6314));
   INVX1 U3783 (.Y(n8277), 
	.A(\ram[174][14] ));
   OAI22X1 U3784 (.Y(n3379), 
	.B1(n8278), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6316));
   INVX1 U3785 (.Y(n8278), 
	.A(\ram[174][13] ));
   OAI22X1 U3786 (.Y(n3378), 
	.B1(n8279), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6318));
   INVX1 U3787 (.Y(n8279), 
	.A(\ram[174][12] ));
   OAI22X1 U3788 (.Y(n3377), 
	.B1(n8280), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6320));
   INVX1 U3789 (.Y(n8280), 
	.A(\ram[174][11] ));
   OAI22X1 U3790 (.Y(n3376), 
	.B1(n8281), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6322));
   INVX1 U3791 (.Y(n8281), 
	.A(\ram[174][10] ));
   OAI22X1 U3792 (.Y(n3375), 
	.B1(n8282), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6324));
   INVX1 U3793 (.Y(n8282), 
	.A(\ram[174][9] ));
   OAI22X1 U3794 (.Y(n3374), 
	.B1(n8283), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6326));
   INVX1 U3795 (.Y(n8283), 
	.A(\ram[174][8] ));
   OAI22X1 U3796 (.Y(n3373), 
	.B1(n8284), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6328));
   INVX1 U3797 (.Y(n8284), 
	.A(\ram[174][7] ));
   OAI22X1 U3798 (.Y(n3372), 
	.B1(n8285), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6330));
   INVX1 U3799 (.Y(n8285), 
	.A(\ram[174][6] ));
   OAI22X1 U3800 (.Y(n3371), 
	.B1(n8286), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6332));
   INVX1 U3801 (.Y(n8286), 
	.A(\ram[174][5] ));
   OAI22X1 U3802 (.Y(n3370), 
	.B1(n8287), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6334));
   INVX1 U3803 (.Y(n8287), 
	.A(\ram[174][4] ));
   OAI22X1 U3804 (.Y(n3369), 
	.B1(n8288), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6336));
   INVX1 U3805 (.Y(n8288), 
	.A(\ram[174][3] ));
   OAI22X1 U3806 (.Y(n3368), 
	.B1(n8289), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6338));
   INVX1 U3807 (.Y(n8289), 
	.A(\ram[174][2] ));
   OAI22X1 U3808 (.Y(n3367), 
	.B1(n8290), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6306));
   INVX1 U3809 (.Y(n8290), 
	.A(\ram[174][1] ));
   OAI22X1 U3810 (.Y(n3366), 
	.B1(n8291), 
	.B0(n8275), 
	.A1(n8274), 
	.A0(n6309));
   INVX1 U3811 (.Y(n8291), 
	.A(\ram[174][0] ));
   NOR2BX1 U3812 (.Y(n8275), 
	.B(n8274), 
	.AN(mem_write_en));
   NAND2X1 U3813 (.Y(n8274), 
	.B(n6553), 
	.A(n8273));
   OAI22X1 U3814 (.Y(n3365), 
	.B1(n8294), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6311));
   INVX1 U3815 (.Y(n8294), 
	.A(\ram[173][15] ));
   OAI22X1 U3816 (.Y(n3364), 
	.B1(n8295), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6314));
   INVX1 U3817 (.Y(n8295), 
	.A(\ram[173][14] ));
   OAI22X1 U3818 (.Y(n3363), 
	.B1(n8296), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6316));
   INVX1 U3819 (.Y(n8296), 
	.A(\ram[173][13] ));
   OAI22X1 U3820 (.Y(n3362), 
	.B1(n8297), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6318));
   INVX1 U3821 (.Y(n8297), 
	.A(\ram[173][12] ));
   OAI22X1 U3822 (.Y(n3361), 
	.B1(n8298), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6320));
   INVX1 U3823 (.Y(n8298), 
	.A(\ram[173][11] ));
   OAI22X1 U3824 (.Y(n3360), 
	.B1(n8299), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6322));
   INVX1 U3825 (.Y(n8299), 
	.A(\ram[173][10] ));
   OAI22X1 U3826 (.Y(n3359), 
	.B1(n8300), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6324));
   INVX1 U3827 (.Y(n8300), 
	.A(\ram[173][9] ));
   OAI22X1 U3828 (.Y(n3358), 
	.B1(n8301), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6326));
   INVX1 U3829 (.Y(n8301), 
	.A(\ram[173][8] ));
   OAI22X1 U3830 (.Y(n3357), 
	.B1(n8302), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6328));
   INVX1 U3831 (.Y(n8302), 
	.A(\ram[173][7] ));
   OAI22X1 U3832 (.Y(n3356), 
	.B1(n8303), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6330));
   INVX1 U3833 (.Y(n8303), 
	.A(\ram[173][6] ));
   OAI22X1 U3834 (.Y(n3355), 
	.B1(n8304), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6332));
   INVX1 U3835 (.Y(n8304), 
	.A(\ram[173][5] ));
   OAI22X1 U3836 (.Y(n3354), 
	.B1(n8305), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6334));
   INVX1 U3837 (.Y(n8305), 
	.A(\ram[173][4] ));
   OAI22X1 U3838 (.Y(n3353), 
	.B1(n8306), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6336));
   INVX1 U3839 (.Y(n8306), 
	.A(\ram[173][3] ));
   OAI22X1 U3840 (.Y(n3352), 
	.B1(n8307), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6338));
   INVX1 U3841 (.Y(n8307), 
	.A(\ram[173][2] ));
   OAI22X1 U3842 (.Y(n3351), 
	.B1(n8308), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6306));
   INVX1 U3843 (.Y(n8308), 
	.A(\ram[173][1] ));
   OAI22X1 U3844 (.Y(n3350), 
	.B1(n8309), 
	.B0(n8293), 
	.A1(n8292), 
	.A0(n6309));
   INVX1 U3845 (.Y(n8309), 
	.A(\ram[173][0] ));
   NOR2BX1 U3846 (.Y(n8293), 
	.B(n8292), 
	.AN(mem_write_en));
   NAND2X1 U3847 (.Y(n8292), 
	.B(n6572), 
	.A(n8273));
   OAI22X1 U3848 (.Y(n3349), 
	.B1(n8312), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6311));
   INVX1 U3849 (.Y(n8312), 
	.A(\ram[172][15] ));
   OAI22X1 U3850 (.Y(n3348), 
	.B1(n8313), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6314));
   INVX1 U3851 (.Y(n8313), 
	.A(\ram[172][14] ));
   OAI22X1 U3852 (.Y(n3347), 
	.B1(n8314), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6316));
   INVX1 U3853 (.Y(n8314), 
	.A(\ram[172][13] ));
   OAI22X1 U3854 (.Y(n3346), 
	.B1(n8315), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6318));
   INVX1 U3855 (.Y(n8315), 
	.A(\ram[172][12] ));
   OAI22X1 U3856 (.Y(n3345), 
	.B1(n8316), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6320));
   INVX1 U3857 (.Y(n8316), 
	.A(\ram[172][11] ));
   OAI22X1 U3858 (.Y(n3344), 
	.B1(n8317), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6322));
   INVX1 U3859 (.Y(n8317), 
	.A(\ram[172][10] ));
   OAI22X1 U3860 (.Y(n3343), 
	.B1(n8318), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6324));
   INVX1 U3861 (.Y(n8318), 
	.A(\ram[172][9] ));
   OAI22X1 U3862 (.Y(n3342), 
	.B1(n8319), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6326));
   INVX1 U3863 (.Y(n8319), 
	.A(\ram[172][8] ));
   OAI22X1 U3864 (.Y(n3341), 
	.B1(n8320), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6328));
   INVX1 U3865 (.Y(n8320), 
	.A(\ram[172][7] ));
   OAI22X1 U3866 (.Y(n3340), 
	.B1(n8321), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6330));
   INVX1 U3867 (.Y(n8321), 
	.A(\ram[172][6] ));
   OAI22X1 U3868 (.Y(n3339), 
	.B1(n8322), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6332));
   INVX1 U3869 (.Y(n8322), 
	.A(\ram[172][5] ));
   OAI22X1 U3870 (.Y(n3338), 
	.B1(n8323), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6334));
   INVX1 U3871 (.Y(n8323), 
	.A(\ram[172][4] ));
   OAI22X1 U3872 (.Y(n3337), 
	.B1(n8324), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6336));
   INVX1 U3873 (.Y(n8324), 
	.A(\ram[172][3] ));
   OAI22X1 U3874 (.Y(n3336), 
	.B1(n8325), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6338));
   INVX1 U3875 (.Y(n8325), 
	.A(\ram[172][2] ));
   OAI22X1 U3876 (.Y(n3335), 
	.B1(n8326), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6306));
   INVX1 U3877 (.Y(n8326), 
	.A(\ram[172][1] ));
   OAI22X1 U3878 (.Y(n3334), 
	.B1(n8327), 
	.B0(n8311), 
	.A1(n8310), 
	.A0(n6309));
   INVX1 U3879 (.Y(n8327), 
	.A(\ram[172][0] ));
   NOR2BX1 U3880 (.Y(n8311), 
	.B(n8310), 
	.AN(mem_write_en));
   NAND2X1 U3881 (.Y(n8310), 
	.B(n6591), 
	.A(n8273));
   OAI22X1 U3882 (.Y(n3333), 
	.B1(n8330), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6311));
   INVX1 U3883 (.Y(n8330), 
	.A(\ram[171][15] ));
   OAI22X1 U3884 (.Y(n3332), 
	.B1(n8331), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6314));
   INVX1 U3885 (.Y(n8331), 
	.A(\ram[171][14] ));
   OAI22X1 U3886 (.Y(n3331), 
	.B1(n8332), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6316));
   INVX1 U3887 (.Y(n8332), 
	.A(\ram[171][13] ));
   OAI22X1 U3888 (.Y(n3330), 
	.B1(n8333), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6318));
   INVX1 U3889 (.Y(n8333), 
	.A(\ram[171][12] ));
   OAI22X1 U3890 (.Y(n3329), 
	.B1(n8334), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6320));
   INVX1 U3891 (.Y(n8334), 
	.A(\ram[171][11] ));
   OAI22X1 U3892 (.Y(n3328), 
	.B1(n8335), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6322));
   INVX1 U3893 (.Y(n8335), 
	.A(\ram[171][10] ));
   OAI22X1 U3894 (.Y(n3327), 
	.B1(n8336), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6324));
   INVX1 U3895 (.Y(n8336), 
	.A(\ram[171][9] ));
   OAI22X1 U3896 (.Y(n3326), 
	.B1(n8337), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6326));
   INVX1 U3897 (.Y(n8337), 
	.A(\ram[171][8] ));
   OAI22X1 U3898 (.Y(n3325), 
	.B1(n8338), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6328));
   INVX1 U3899 (.Y(n8338), 
	.A(\ram[171][7] ));
   OAI22X1 U3900 (.Y(n3324), 
	.B1(n8339), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6330));
   INVX1 U3901 (.Y(n8339), 
	.A(\ram[171][6] ));
   OAI22X1 U3902 (.Y(n3323), 
	.B1(n8340), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6332));
   INVX1 U3903 (.Y(n8340), 
	.A(\ram[171][5] ));
   OAI22X1 U3904 (.Y(n3322), 
	.B1(n8341), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6334));
   INVX1 U3905 (.Y(n8341), 
	.A(\ram[171][4] ));
   OAI22X1 U3906 (.Y(n3321), 
	.B1(n8342), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6336));
   INVX1 U3907 (.Y(n8342), 
	.A(\ram[171][3] ));
   OAI22X1 U3908 (.Y(n3320), 
	.B1(n8343), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6338));
   INVX1 U3909 (.Y(n8343), 
	.A(\ram[171][2] ));
   OAI22X1 U3910 (.Y(n3319), 
	.B1(n8344), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6306));
   INVX1 U3911 (.Y(n8344), 
	.A(\ram[171][1] ));
   OAI22X1 U3912 (.Y(n3318), 
	.B1(n8345), 
	.B0(n8329), 
	.A1(n8328), 
	.A0(n6309));
   INVX1 U3913 (.Y(n8345), 
	.A(\ram[171][0] ));
   NOR2BX1 U3914 (.Y(n8329), 
	.B(n8328), 
	.AN(mem_write_en));
   NAND2X1 U3915 (.Y(n8328), 
	.B(n6610), 
	.A(n8273));
   OAI22X1 U3916 (.Y(n3317), 
	.B1(n8348), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6311));
   INVX1 U3917 (.Y(n8348), 
	.A(\ram[170][15] ));
   OAI22X1 U3918 (.Y(n3316), 
	.B1(n8349), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6314));
   INVX1 U3919 (.Y(n8349), 
	.A(\ram[170][14] ));
   OAI22X1 U3920 (.Y(n3315), 
	.B1(n8350), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6316));
   INVX1 U3921 (.Y(n8350), 
	.A(\ram[170][13] ));
   OAI22X1 U3922 (.Y(n3314), 
	.B1(n8351), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6318));
   INVX1 U3923 (.Y(n8351), 
	.A(\ram[170][12] ));
   OAI22X1 U3924 (.Y(n3313), 
	.B1(n8352), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6320));
   INVX1 U3925 (.Y(n8352), 
	.A(\ram[170][11] ));
   OAI22X1 U3926 (.Y(n3312), 
	.B1(n8353), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6322));
   INVX1 U3927 (.Y(n8353), 
	.A(\ram[170][10] ));
   OAI22X1 U3928 (.Y(n3311), 
	.B1(n8354), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6324));
   INVX1 U3929 (.Y(n8354), 
	.A(\ram[170][9] ));
   OAI22X1 U3930 (.Y(n3310), 
	.B1(n8355), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6326));
   INVX1 U3931 (.Y(n8355), 
	.A(\ram[170][8] ));
   OAI22X1 U3932 (.Y(n3309), 
	.B1(n8356), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6328));
   INVX1 U3933 (.Y(n8356), 
	.A(\ram[170][7] ));
   OAI22X1 U3934 (.Y(n3308), 
	.B1(n8357), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6330));
   INVX1 U3935 (.Y(n8357), 
	.A(\ram[170][6] ));
   OAI22X1 U3936 (.Y(n3307), 
	.B1(n8358), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6332));
   INVX1 U3937 (.Y(n8358), 
	.A(\ram[170][5] ));
   OAI22X1 U3938 (.Y(n3306), 
	.B1(n8359), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6334));
   INVX1 U3939 (.Y(n8359), 
	.A(\ram[170][4] ));
   OAI22X1 U3940 (.Y(n3305), 
	.B1(n8360), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6336));
   INVX1 U3941 (.Y(n8360), 
	.A(\ram[170][3] ));
   OAI22X1 U3942 (.Y(n3304), 
	.B1(n8361), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6338));
   INVX1 U3943 (.Y(n8361), 
	.A(\ram[170][2] ));
   OAI22X1 U3944 (.Y(n3303), 
	.B1(n8362), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6306));
   INVX1 U3945 (.Y(n8362), 
	.A(\ram[170][1] ));
   OAI22X1 U3946 (.Y(n3302), 
	.B1(n8363), 
	.B0(n8347), 
	.A1(n8346), 
	.A0(n6309));
   INVX1 U3947 (.Y(n8363), 
	.A(\ram[170][0] ));
   NOR2BX1 U3948 (.Y(n8347), 
	.B(n8346), 
	.AN(mem_write_en));
   NAND2X1 U3949 (.Y(n8346), 
	.B(n6629), 
	.A(n8273));
   OAI22X1 U3950 (.Y(n3301), 
	.B1(n8366), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6311));
   INVX1 U3951 (.Y(n8366), 
	.A(\ram[169][15] ));
   OAI22X1 U3952 (.Y(n3300), 
	.B1(n8367), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6314));
   INVX1 U3953 (.Y(n8367), 
	.A(\ram[169][14] ));
   OAI22X1 U3954 (.Y(n3299), 
	.B1(n8368), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6316));
   INVX1 U3955 (.Y(n8368), 
	.A(\ram[169][13] ));
   OAI22X1 U3956 (.Y(n3298), 
	.B1(n8369), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6318));
   INVX1 U3957 (.Y(n8369), 
	.A(\ram[169][12] ));
   OAI22X1 U3958 (.Y(n3297), 
	.B1(n8370), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6320));
   INVX1 U3959 (.Y(n8370), 
	.A(\ram[169][11] ));
   OAI22X1 U3960 (.Y(n3296), 
	.B1(n8371), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6322));
   INVX1 U3961 (.Y(n8371), 
	.A(\ram[169][10] ));
   OAI22X1 U3962 (.Y(n3295), 
	.B1(n8372), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6324));
   INVX1 U3963 (.Y(n8372), 
	.A(\ram[169][9] ));
   OAI22X1 U3964 (.Y(n3294), 
	.B1(n8373), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6326));
   INVX1 U3965 (.Y(n8373), 
	.A(\ram[169][8] ));
   OAI22X1 U3966 (.Y(n3293), 
	.B1(n8374), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6328));
   INVX1 U3967 (.Y(n8374), 
	.A(\ram[169][7] ));
   OAI22X1 U3968 (.Y(n3292), 
	.B1(n8375), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6330));
   INVX1 U3969 (.Y(n8375), 
	.A(\ram[169][6] ));
   OAI22X1 U3970 (.Y(n3291), 
	.B1(n8376), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6332));
   INVX1 U3971 (.Y(n8376), 
	.A(\ram[169][5] ));
   OAI22X1 U3972 (.Y(n3290), 
	.B1(n8377), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6334));
   INVX1 U3973 (.Y(n8377), 
	.A(\ram[169][4] ));
   OAI22X1 U3974 (.Y(n3289), 
	.B1(n8378), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6336));
   INVX1 U3975 (.Y(n8378), 
	.A(\ram[169][3] ));
   OAI22X1 U3976 (.Y(n3288), 
	.B1(n8379), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6338));
   INVX1 U3977 (.Y(n8379), 
	.A(\ram[169][2] ));
   OAI22X1 U3978 (.Y(n3287), 
	.B1(n8380), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6306));
   INVX1 U3979 (.Y(n8380), 
	.A(\ram[169][1] ));
   OAI22X1 U3980 (.Y(n3286), 
	.B1(n8381), 
	.B0(n8365), 
	.A1(n8364), 
	.A0(n6309));
   INVX1 U3981 (.Y(n8381), 
	.A(\ram[169][0] ));
   NOR2BX1 U3982 (.Y(n8365), 
	.B(n8364), 
	.AN(mem_write_en));
   NAND2X1 U3983 (.Y(n8364), 
	.B(n6342), 
	.A(n8273));
   OAI22X1 U3984 (.Y(n3285), 
	.B1(n8384), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6311));
   INVX1 U3985 (.Y(n8384), 
	.A(\ram[168][15] ));
   OAI22X1 U3986 (.Y(n3284), 
	.B1(n8385), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6314));
   INVX1 U3987 (.Y(n8385), 
	.A(\ram[168][14] ));
   OAI22X1 U3988 (.Y(n3283), 
	.B1(n8386), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6316));
   INVX1 U3989 (.Y(n8386), 
	.A(\ram[168][13] ));
   OAI22X1 U3990 (.Y(n3282), 
	.B1(n8387), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6318));
   INVX1 U3991 (.Y(n8387), 
	.A(\ram[168][12] ));
   OAI22X1 U3992 (.Y(n3281), 
	.B1(n8388), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6320));
   INVX1 U3993 (.Y(n8388), 
	.A(\ram[168][11] ));
   OAI22X1 U3994 (.Y(n3280), 
	.B1(n8389), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6322));
   INVX1 U3995 (.Y(n8389), 
	.A(\ram[168][10] ));
   OAI22X1 U3996 (.Y(n3279), 
	.B1(n8390), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6324));
   INVX1 U3997 (.Y(n8390), 
	.A(\ram[168][9] ));
   OAI22X1 U3998 (.Y(n3278), 
	.B1(n8391), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6326));
   INVX1 U3999 (.Y(n8391), 
	.A(\ram[168][8] ));
   OAI22X1 U4000 (.Y(n3277), 
	.B1(n8392), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6328));
   INVX1 U4001 (.Y(n8392), 
	.A(\ram[168][7] ));
   OAI22X1 U4002 (.Y(n3276), 
	.B1(n8393), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6330));
   INVX1 U4003 (.Y(n8393), 
	.A(\ram[168][6] ));
   OAI22X1 U4004 (.Y(n3275), 
	.B1(n8394), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6332));
   INVX1 U4005 (.Y(n8394), 
	.A(\ram[168][5] ));
   OAI22X1 U4006 (.Y(n3274), 
	.B1(n8395), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6334));
   INVX1 U4007 (.Y(n8395), 
	.A(\ram[168][4] ));
   OAI22X1 U4008 (.Y(n3273), 
	.B1(n8396), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6336));
   INVX1 U4009 (.Y(n8396), 
	.A(\ram[168][3] ));
   OAI22X1 U4010 (.Y(n3272), 
	.B1(n8397), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6338));
   INVX1 U4011 (.Y(n8397), 
	.A(\ram[168][2] ));
   OAI22X1 U4012 (.Y(n3271), 
	.B1(n8398), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6306));
   INVX1 U4013 (.Y(n8398), 
	.A(\ram[168][1] ));
   OAI22X1 U4014 (.Y(n3270), 
	.B1(n8399), 
	.B0(n8383), 
	.A1(n8382), 
	.A0(n6309));
   INVX1 U4015 (.Y(n8399), 
	.A(\ram[168][0] ));
   NOR2BX1 U4016 (.Y(n8383), 
	.B(n8382), 
	.AN(mem_write_en));
   NAND2X1 U4017 (.Y(n8382), 
	.B(n6362), 
	.A(n8273));
   OAI22X1 U4018 (.Y(n3269), 
	.B1(n8402), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6311));
   INVX1 U4019 (.Y(n8402), 
	.A(\ram[167][15] ));
   OAI22X1 U4020 (.Y(n3268), 
	.B1(n8403), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6314));
   INVX1 U4021 (.Y(n8403), 
	.A(\ram[167][14] ));
   OAI22X1 U4022 (.Y(n3267), 
	.B1(n8404), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6316));
   INVX1 U4023 (.Y(n8404), 
	.A(\ram[167][13] ));
   OAI22X1 U4024 (.Y(n3266), 
	.B1(n8405), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6318));
   INVX1 U4025 (.Y(n8405), 
	.A(\ram[167][12] ));
   OAI22X1 U4026 (.Y(n3265), 
	.B1(n8406), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6320));
   INVX1 U4027 (.Y(n8406), 
	.A(\ram[167][11] ));
   OAI22X1 U4028 (.Y(n3264), 
	.B1(n8407), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6322));
   INVX1 U4029 (.Y(n8407), 
	.A(\ram[167][10] ));
   OAI22X1 U4030 (.Y(n3263), 
	.B1(n8408), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6324));
   INVX1 U4031 (.Y(n8408), 
	.A(\ram[167][9] ));
   OAI22X1 U4032 (.Y(n3262), 
	.B1(n8409), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6326));
   INVX1 U4033 (.Y(n8409), 
	.A(\ram[167][8] ));
   OAI22X1 U4034 (.Y(n3261), 
	.B1(n8410), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6328));
   INVX1 U4035 (.Y(n8410), 
	.A(\ram[167][7] ));
   OAI22X1 U4036 (.Y(n3260), 
	.B1(n8411), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6330));
   INVX1 U4037 (.Y(n8411), 
	.A(\ram[167][6] ));
   OAI22X1 U4038 (.Y(n3259), 
	.B1(n8412), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6332));
   INVX1 U4039 (.Y(n8412), 
	.A(\ram[167][5] ));
   OAI22X1 U4040 (.Y(n3258), 
	.B1(n8413), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6334));
   INVX1 U4041 (.Y(n8413), 
	.A(\ram[167][4] ));
   OAI22X1 U4042 (.Y(n3257), 
	.B1(n8414), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6336));
   INVX1 U4043 (.Y(n8414), 
	.A(\ram[167][3] ));
   OAI22X1 U4044 (.Y(n3256), 
	.B1(n8415), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6338));
   INVX1 U4045 (.Y(n8415), 
	.A(\ram[167][2] ));
   OAI22X1 U4046 (.Y(n3255), 
	.B1(n8416), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6306));
   INVX1 U4047 (.Y(n8416), 
	.A(\ram[167][1] ));
   OAI22X1 U4048 (.Y(n3254), 
	.B1(n8417), 
	.B0(n8401), 
	.A1(n8400), 
	.A0(n6309));
   INVX1 U4049 (.Y(n8417), 
	.A(\ram[167][0] ));
   NOR2BX1 U4050 (.Y(n8401), 
	.B(n8400), 
	.AN(mem_write_en));
   NAND2X1 U4051 (.Y(n8400), 
	.B(n6381), 
	.A(n8273));
   OAI22X1 U4052 (.Y(n3253), 
	.B1(n8420), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6311));
   INVX1 U4053 (.Y(n8420), 
	.A(\ram[166][15] ));
   OAI22X1 U4054 (.Y(n3252), 
	.B1(n8421), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6314));
   INVX1 U4055 (.Y(n8421), 
	.A(\ram[166][14] ));
   OAI22X1 U4056 (.Y(n3251), 
	.B1(n8422), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6316));
   INVX1 U4057 (.Y(n8422), 
	.A(\ram[166][13] ));
   OAI22X1 U4058 (.Y(n3250), 
	.B1(n8423), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6318));
   INVX1 U4059 (.Y(n8423), 
	.A(\ram[166][12] ));
   OAI22X1 U4060 (.Y(n3249), 
	.B1(n8424), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6320));
   INVX1 U4061 (.Y(n8424), 
	.A(\ram[166][11] ));
   OAI22X1 U4062 (.Y(n3248), 
	.B1(n8425), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6322));
   INVX1 U4063 (.Y(n8425), 
	.A(\ram[166][10] ));
   OAI22X1 U4064 (.Y(n3247), 
	.B1(n8426), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6324));
   INVX1 U4065 (.Y(n8426), 
	.A(\ram[166][9] ));
   OAI22X1 U4066 (.Y(n3246), 
	.B1(n8427), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6326));
   INVX1 U4067 (.Y(n8427), 
	.A(\ram[166][8] ));
   OAI22X1 U4068 (.Y(n3245), 
	.B1(n8428), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6328));
   INVX1 U4069 (.Y(n8428), 
	.A(\ram[166][7] ));
   OAI22X1 U4070 (.Y(n3244), 
	.B1(n8429), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6330));
   INVX1 U4071 (.Y(n8429), 
	.A(\ram[166][6] ));
   OAI22X1 U4072 (.Y(n3243), 
	.B1(n8430), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6332));
   INVX1 U4073 (.Y(n8430), 
	.A(\ram[166][5] ));
   OAI22X1 U4074 (.Y(n3242), 
	.B1(n8431), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6334));
   INVX1 U4075 (.Y(n8431), 
	.A(\ram[166][4] ));
   OAI22X1 U4076 (.Y(n3241), 
	.B1(n8432), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6336));
   INVX1 U4077 (.Y(n8432), 
	.A(\ram[166][3] ));
   OAI22X1 U4078 (.Y(n3240), 
	.B1(n8433), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6338));
   INVX1 U4079 (.Y(n8433), 
	.A(\ram[166][2] ));
   OAI22X1 U4080 (.Y(n3239), 
	.B1(n8434), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6306));
   INVX1 U4081 (.Y(n8434), 
	.A(\ram[166][1] ));
   OAI22X1 U4082 (.Y(n3238), 
	.B1(n8435), 
	.B0(n8419), 
	.A1(n8418), 
	.A0(n6309));
   INVX1 U4083 (.Y(n8435), 
	.A(\ram[166][0] ));
   NOR2BX1 U4084 (.Y(n8419), 
	.B(n8418), 
	.AN(mem_write_en));
   NAND2X1 U4085 (.Y(n8418), 
	.B(n6400), 
	.A(n8273));
   OAI22X1 U4086 (.Y(n3237), 
	.B1(n8438), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6311));
   INVX1 U4087 (.Y(n8438), 
	.A(\ram[165][15] ));
   OAI22X1 U4088 (.Y(n3236), 
	.B1(n8439), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6314));
   INVX1 U4089 (.Y(n8439), 
	.A(\ram[165][14] ));
   OAI22X1 U4090 (.Y(n3235), 
	.B1(n8440), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6316));
   INVX1 U4091 (.Y(n8440), 
	.A(\ram[165][13] ));
   OAI22X1 U4092 (.Y(n3234), 
	.B1(n8441), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6318));
   INVX1 U4093 (.Y(n8441), 
	.A(\ram[165][12] ));
   OAI22X1 U4094 (.Y(n3233), 
	.B1(n8442), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6320));
   INVX1 U4095 (.Y(n8442), 
	.A(\ram[165][11] ));
   OAI22X1 U4096 (.Y(n3232), 
	.B1(n8443), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6322));
   INVX1 U4097 (.Y(n8443), 
	.A(\ram[165][10] ));
   OAI22X1 U4098 (.Y(n3231), 
	.B1(n8444), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6324));
   INVX1 U4099 (.Y(n8444), 
	.A(\ram[165][9] ));
   OAI22X1 U4100 (.Y(n3230), 
	.B1(n8445), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6326));
   INVX1 U4101 (.Y(n8445), 
	.A(\ram[165][8] ));
   OAI22X1 U4102 (.Y(n3229), 
	.B1(n8446), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6328));
   INVX1 U4103 (.Y(n8446), 
	.A(\ram[165][7] ));
   OAI22X1 U4104 (.Y(n3228), 
	.B1(n8447), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6330));
   INVX1 U4105 (.Y(n8447), 
	.A(\ram[165][6] ));
   OAI22X1 U4106 (.Y(n3227), 
	.B1(n8448), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6332));
   INVX1 U4107 (.Y(n8448), 
	.A(\ram[165][5] ));
   OAI22X1 U4108 (.Y(n3226), 
	.B1(n8449), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6334));
   INVX1 U4109 (.Y(n8449), 
	.A(\ram[165][4] ));
   OAI22X1 U4110 (.Y(n3225), 
	.B1(n8450), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6336));
   INVX1 U4111 (.Y(n8450), 
	.A(\ram[165][3] ));
   OAI22X1 U4112 (.Y(n3224), 
	.B1(n8451), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6338));
   INVX1 U4113 (.Y(n8451), 
	.A(\ram[165][2] ));
   OAI22X1 U4114 (.Y(n3223), 
	.B1(n8452), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6306));
   INVX1 U4115 (.Y(n8452), 
	.A(\ram[165][1] ));
   OAI22X1 U4116 (.Y(n3222), 
	.B1(n8453), 
	.B0(n8437), 
	.A1(n8436), 
	.A0(n6309));
   INVX1 U4117 (.Y(n8453), 
	.A(\ram[165][0] ));
   NOR2BX1 U4118 (.Y(n8437), 
	.B(n8436), 
	.AN(mem_write_en));
   NAND2X1 U4119 (.Y(n8436), 
	.B(n6419), 
	.A(n8273));
   OAI22X1 U4120 (.Y(n3221), 
	.B1(n8456), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6311));
   INVX1 U4121 (.Y(n8456), 
	.A(\ram[164][15] ));
   OAI22X1 U4122 (.Y(n3220), 
	.B1(n8457), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6314));
   INVX1 U4123 (.Y(n8457), 
	.A(\ram[164][14] ));
   OAI22X1 U4124 (.Y(n3219), 
	.B1(n8458), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6316));
   INVX1 U4125 (.Y(n8458), 
	.A(\ram[164][13] ));
   OAI22X1 U4126 (.Y(n3218), 
	.B1(n8459), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6318));
   INVX1 U4127 (.Y(n8459), 
	.A(\ram[164][12] ));
   OAI22X1 U4128 (.Y(n3217), 
	.B1(n8460), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6320));
   INVX1 U4129 (.Y(n8460), 
	.A(\ram[164][11] ));
   OAI22X1 U4130 (.Y(n3216), 
	.B1(n8461), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6322));
   INVX1 U4131 (.Y(n8461), 
	.A(\ram[164][10] ));
   OAI22X1 U4132 (.Y(n3215), 
	.B1(n8462), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6324));
   INVX1 U4133 (.Y(n8462), 
	.A(\ram[164][9] ));
   OAI22X1 U4134 (.Y(n3214), 
	.B1(n8463), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6326));
   INVX1 U4135 (.Y(n8463), 
	.A(\ram[164][8] ));
   OAI22X1 U4136 (.Y(n3213), 
	.B1(n8464), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6328));
   INVX1 U4137 (.Y(n8464), 
	.A(\ram[164][7] ));
   OAI22X1 U4138 (.Y(n3212), 
	.B1(n8465), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6330));
   INVX1 U4139 (.Y(n8465), 
	.A(\ram[164][6] ));
   OAI22X1 U4140 (.Y(n3211), 
	.B1(n8466), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6332));
   INVX1 U4141 (.Y(n8466), 
	.A(\ram[164][5] ));
   OAI22X1 U4142 (.Y(n3210), 
	.B1(n8467), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6334));
   INVX1 U4143 (.Y(n8467), 
	.A(\ram[164][4] ));
   OAI22X1 U4144 (.Y(n3209), 
	.B1(n8468), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6336));
   INVX1 U4145 (.Y(n8468), 
	.A(\ram[164][3] ));
   OAI22X1 U4146 (.Y(n3208), 
	.B1(n8469), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6338));
   INVX1 U4147 (.Y(n8469), 
	.A(\ram[164][2] ));
   OAI22X1 U4148 (.Y(n3207), 
	.B1(n8470), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6306));
   INVX1 U4149 (.Y(n8470), 
	.A(\ram[164][1] ));
   OAI22X1 U4150 (.Y(n3206), 
	.B1(n8471), 
	.B0(n8455), 
	.A1(n8454), 
	.A0(n6309));
   INVX1 U4151 (.Y(n8471), 
	.A(\ram[164][0] ));
   NOR2BX1 U4152 (.Y(n8455), 
	.B(n8454), 
	.AN(mem_write_en));
   NAND2X1 U4153 (.Y(n8454), 
	.B(n6438), 
	.A(n8273));
   OAI22X1 U4154 (.Y(n3205), 
	.B1(n8474), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6311));
   INVX1 U4155 (.Y(n8474), 
	.A(\ram[163][15] ));
   OAI22X1 U4156 (.Y(n3204), 
	.B1(n8475), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6314));
   INVX1 U4157 (.Y(n8475), 
	.A(\ram[163][14] ));
   OAI22X1 U4158 (.Y(n3203), 
	.B1(n8476), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6316));
   INVX1 U4159 (.Y(n8476), 
	.A(\ram[163][13] ));
   OAI22X1 U4160 (.Y(n3202), 
	.B1(n8477), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6318));
   INVX1 U4161 (.Y(n8477), 
	.A(\ram[163][12] ));
   OAI22X1 U4162 (.Y(n3201), 
	.B1(n8478), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6320));
   INVX1 U4163 (.Y(n8478), 
	.A(\ram[163][11] ));
   OAI22X1 U4164 (.Y(n3200), 
	.B1(n8479), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6322));
   INVX1 U4165 (.Y(n8479), 
	.A(\ram[163][10] ));
   OAI22X1 U4166 (.Y(n3199), 
	.B1(n8480), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6324));
   INVX1 U4167 (.Y(n8480), 
	.A(\ram[163][9] ));
   OAI22X1 U4168 (.Y(n3198), 
	.B1(n8481), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6326));
   INVX1 U4169 (.Y(n8481), 
	.A(\ram[163][8] ));
   OAI22X1 U4170 (.Y(n3197), 
	.B1(n8482), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6328));
   INVX1 U4171 (.Y(n8482), 
	.A(\ram[163][7] ));
   OAI22X1 U4172 (.Y(n3196), 
	.B1(n8483), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6330));
   INVX1 U4173 (.Y(n8483), 
	.A(\ram[163][6] ));
   OAI22X1 U4174 (.Y(n3195), 
	.B1(n8484), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6332));
   INVX1 U4175 (.Y(n8484), 
	.A(\ram[163][5] ));
   OAI22X1 U4176 (.Y(n3194), 
	.B1(n8485), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6334));
   INVX1 U4177 (.Y(n8485), 
	.A(\ram[163][4] ));
   OAI22X1 U4178 (.Y(n3193), 
	.B1(n8486), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6336));
   INVX1 U4179 (.Y(n8486), 
	.A(\ram[163][3] ));
   OAI22X1 U4180 (.Y(n3192), 
	.B1(n8487), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6338));
   INVX1 U4181 (.Y(n8487), 
	.A(\ram[163][2] ));
   OAI22X1 U4182 (.Y(n3191), 
	.B1(n8488), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6306));
   INVX1 U4183 (.Y(n8488), 
	.A(\ram[163][1] ));
   OAI22X1 U4184 (.Y(n3190), 
	.B1(n8489), 
	.B0(n8473), 
	.A1(n8472), 
	.A0(n6309));
   INVX1 U4185 (.Y(n8489), 
	.A(\ram[163][0] ));
   NOR2BX1 U4186 (.Y(n8473), 
	.B(n8472), 
	.AN(mem_write_en));
   NAND2X1 U4187 (.Y(n8472), 
	.B(n6457), 
	.A(n8273));
   OAI22X1 U4188 (.Y(n3189), 
	.B1(n8492), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6311));
   INVX1 U4189 (.Y(n8492), 
	.A(\ram[162][15] ));
   OAI22X1 U4190 (.Y(n3188), 
	.B1(n8493), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6314));
   INVX1 U4191 (.Y(n8493), 
	.A(\ram[162][14] ));
   OAI22X1 U4192 (.Y(n3187), 
	.B1(n8494), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6316));
   INVX1 U4193 (.Y(n8494), 
	.A(\ram[162][13] ));
   OAI22X1 U4194 (.Y(n3186), 
	.B1(n8495), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6318));
   INVX1 U4195 (.Y(n8495), 
	.A(\ram[162][12] ));
   OAI22X1 U4196 (.Y(n3185), 
	.B1(n8496), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6320));
   INVX1 U4197 (.Y(n8496), 
	.A(\ram[162][11] ));
   OAI22X1 U4198 (.Y(n3184), 
	.B1(n8497), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6322));
   INVX1 U4199 (.Y(n8497), 
	.A(\ram[162][10] ));
   OAI22X1 U4200 (.Y(n3183), 
	.B1(n8498), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6324));
   INVX1 U4201 (.Y(n8498), 
	.A(\ram[162][9] ));
   OAI22X1 U4202 (.Y(n3182), 
	.B1(n8499), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6326));
   INVX1 U4203 (.Y(n8499), 
	.A(\ram[162][8] ));
   OAI22X1 U4204 (.Y(n3181), 
	.B1(n8500), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6328));
   INVX1 U4205 (.Y(n8500), 
	.A(\ram[162][7] ));
   OAI22X1 U4206 (.Y(n3180), 
	.B1(n8501), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6330));
   INVX1 U4207 (.Y(n8501), 
	.A(\ram[162][6] ));
   OAI22X1 U4208 (.Y(n3179), 
	.B1(n8502), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6332));
   INVX1 U4209 (.Y(n8502), 
	.A(\ram[162][5] ));
   OAI22X1 U4210 (.Y(n3178), 
	.B1(n8503), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6334));
   INVX1 U4211 (.Y(n8503), 
	.A(\ram[162][4] ));
   OAI22X1 U4212 (.Y(n3177), 
	.B1(n8504), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6336));
   INVX1 U4213 (.Y(n8504), 
	.A(\ram[162][3] ));
   OAI22X1 U4214 (.Y(n3176), 
	.B1(n8505), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6338));
   INVX1 U4215 (.Y(n8505), 
	.A(\ram[162][2] ));
   OAI22X1 U4216 (.Y(n3175), 
	.B1(n8506), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6306));
   INVX1 U4217 (.Y(n8506), 
	.A(\ram[162][1] ));
   OAI22X1 U4218 (.Y(n3174), 
	.B1(n8507), 
	.B0(n8491), 
	.A1(n8490), 
	.A0(n6309));
   INVX1 U4219 (.Y(n8507), 
	.A(\ram[162][0] ));
   NOR2BX1 U4220 (.Y(n8491), 
	.B(n8490), 
	.AN(mem_write_en));
   NAND2X1 U4221 (.Y(n8490), 
	.B(n6476), 
	.A(n8273));
   OAI22X1 U4222 (.Y(n3173), 
	.B1(n8510), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6311));
   INVX1 U4223 (.Y(n8510), 
	.A(\ram[161][15] ));
   OAI22X1 U4224 (.Y(n3172), 
	.B1(n8511), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6314));
   INVX1 U4225 (.Y(n8511), 
	.A(\ram[161][14] ));
   OAI22X1 U4226 (.Y(n3171), 
	.B1(n8512), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6316));
   INVX1 U4227 (.Y(n8512), 
	.A(\ram[161][13] ));
   OAI22X1 U4228 (.Y(n3170), 
	.B1(n8513), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6318));
   INVX1 U4229 (.Y(n8513), 
	.A(\ram[161][12] ));
   OAI22X1 U4230 (.Y(n3169), 
	.B1(n8514), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6320));
   INVX1 U4231 (.Y(n8514), 
	.A(\ram[161][11] ));
   OAI22X1 U4232 (.Y(n3168), 
	.B1(n8515), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6322));
   INVX1 U4233 (.Y(n8515), 
	.A(\ram[161][10] ));
   OAI22X1 U4234 (.Y(n3167), 
	.B1(n8516), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6324));
   INVX1 U4235 (.Y(n8516), 
	.A(\ram[161][9] ));
   OAI22X1 U4236 (.Y(n3166), 
	.B1(n8517), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6326));
   INVX1 U4237 (.Y(n8517), 
	.A(\ram[161][8] ));
   OAI22X1 U4238 (.Y(n3165), 
	.B1(n8518), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6328));
   INVX1 U4239 (.Y(n8518), 
	.A(\ram[161][7] ));
   OAI22X1 U4240 (.Y(n3164), 
	.B1(n8519), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6330));
   INVX1 U4241 (.Y(n8519), 
	.A(\ram[161][6] ));
   OAI22X1 U4242 (.Y(n3163), 
	.B1(n8520), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6332));
   INVX1 U4243 (.Y(n8520), 
	.A(\ram[161][5] ));
   OAI22X1 U4244 (.Y(n3162), 
	.B1(n8521), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6334));
   INVX1 U4245 (.Y(n8521), 
	.A(\ram[161][4] ));
   OAI22X1 U4246 (.Y(n3161), 
	.B1(n8522), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6336));
   INVX1 U4247 (.Y(n8522), 
	.A(\ram[161][3] ));
   OAI22X1 U4248 (.Y(n3160), 
	.B1(n8523), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6338));
   INVX1 U4249 (.Y(n8523), 
	.A(\ram[161][2] ));
   OAI22X1 U4250 (.Y(n3159), 
	.B1(n8524), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6306));
   INVX1 U4251 (.Y(n8524), 
	.A(\ram[161][1] ));
   OAI22X1 U4252 (.Y(n3158), 
	.B1(n8525), 
	.B0(n8509), 
	.A1(n8508), 
	.A0(n6309));
   INVX1 U4253 (.Y(n8525), 
	.A(\ram[161][0] ));
   NOR2BX1 U4254 (.Y(n8509), 
	.B(n8508), 
	.AN(mem_write_en));
   NAND2X1 U4255 (.Y(n8508), 
	.B(n6495), 
	.A(n8273));
   OAI22X1 U4256 (.Y(n3157), 
	.B1(n8528), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6311));
   INVX1 U4257 (.Y(n8528), 
	.A(\ram[160][15] ));
   OAI22X1 U4258 (.Y(n3156), 
	.B1(n8529), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6314));
   INVX1 U4259 (.Y(n8529), 
	.A(\ram[160][14] ));
   OAI22X1 U4260 (.Y(n3155), 
	.B1(n8530), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6316));
   INVX1 U4261 (.Y(n8530), 
	.A(\ram[160][13] ));
   OAI22X1 U4262 (.Y(n3154), 
	.B1(n8531), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6318));
   INVX1 U4263 (.Y(n8531), 
	.A(\ram[160][12] ));
   OAI22X1 U4264 (.Y(n3153), 
	.B1(n8532), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6320));
   INVX1 U4265 (.Y(n8532), 
	.A(\ram[160][11] ));
   OAI22X1 U4266 (.Y(n3152), 
	.B1(n8533), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6322));
   INVX1 U4267 (.Y(n8533), 
	.A(\ram[160][10] ));
   OAI22X1 U4268 (.Y(n3151), 
	.B1(n8534), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6324));
   INVX1 U4269 (.Y(n8534), 
	.A(\ram[160][9] ));
   OAI22X1 U4270 (.Y(n3150), 
	.B1(n8535), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6326));
   INVX1 U4271 (.Y(n8535), 
	.A(\ram[160][8] ));
   OAI22X1 U4272 (.Y(n3149), 
	.B1(n8536), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6328));
   INVX1 U4273 (.Y(n8536), 
	.A(\ram[160][7] ));
   OAI22X1 U4274 (.Y(n3148), 
	.B1(n8537), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6330));
   INVX1 U4275 (.Y(n8537), 
	.A(\ram[160][6] ));
   OAI22X1 U4276 (.Y(n3147), 
	.B1(n8538), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6332));
   INVX1 U4277 (.Y(n8538), 
	.A(\ram[160][5] ));
   OAI22X1 U4278 (.Y(n3146), 
	.B1(n8539), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6334));
   INVX1 U4279 (.Y(n8539), 
	.A(\ram[160][4] ));
   OAI22X1 U4280 (.Y(n3145), 
	.B1(n8540), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6336));
   INVX1 U4281 (.Y(n8540), 
	.A(\ram[160][3] ));
   OAI22X1 U4282 (.Y(n3144), 
	.B1(n8541), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6338));
   INVX1 U4283 (.Y(n8541), 
	.A(\ram[160][2] ));
   OAI22X1 U4284 (.Y(n3143), 
	.B1(n8542), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6306));
   INVX1 U4285 (.Y(n8542), 
	.A(\ram[160][1] ));
   OAI22X1 U4286 (.Y(n3142), 
	.B1(n8543), 
	.B0(n8527), 
	.A1(n8526), 
	.A0(n6309));
   INVX1 U4287 (.Y(n8543), 
	.A(\ram[160][0] ));
   NOR2BX1 U4288 (.Y(n8527), 
	.B(n8526), 
	.AN(mem_write_en));
   NAND2X1 U4289 (.Y(n8526), 
	.B(n6514), 
	.A(n8273));
   OAI22X1 U4290 (.Y(n3141), 
	.B1(n8546), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6311));
   INVX1 U4291 (.Y(n8546), 
	.A(\ram[159][15] ));
   OAI22X1 U4292 (.Y(n3140), 
	.B1(n8547), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6314));
   INVX1 U4293 (.Y(n8547), 
	.A(\ram[159][14] ));
   OAI22X1 U4294 (.Y(n3139), 
	.B1(n8548), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6316));
   INVX1 U4295 (.Y(n8548), 
	.A(\ram[159][13] ));
   OAI22X1 U4296 (.Y(n3138), 
	.B1(n8549), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6318));
   INVX1 U4297 (.Y(n8549), 
	.A(\ram[159][12] ));
   OAI22X1 U4298 (.Y(n3137), 
	.B1(n8550), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6320));
   INVX1 U4299 (.Y(n8550), 
	.A(\ram[159][11] ));
   OAI22X1 U4300 (.Y(n3136), 
	.B1(n8551), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6322));
   INVX1 U4301 (.Y(n8551), 
	.A(\ram[159][10] ));
   OAI22X1 U4302 (.Y(n3135), 
	.B1(n8552), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6324));
   INVX1 U4303 (.Y(n8552), 
	.A(\ram[159][9] ));
   OAI22X1 U4304 (.Y(n3134), 
	.B1(n8553), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6326));
   INVX1 U4305 (.Y(n8553), 
	.A(\ram[159][8] ));
   OAI22X1 U4306 (.Y(n3133), 
	.B1(n8554), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6328));
   INVX1 U4307 (.Y(n8554), 
	.A(\ram[159][7] ));
   OAI22X1 U4308 (.Y(n3132), 
	.B1(n8555), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6330));
   INVX1 U4309 (.Y(n8555), 
	.A(\ram[159][6] ));
   OAI22X1 U4310 (.Y(n3131), 
	.B1(n8556), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6332));
   INVX1 U4311 (.Y(n8556), 
	.A(\ram[159][5] ));
   OAI22X1 U4312 (.Y(n3130), 
	.B1(n8557), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6334));
   INVX1 U4313 (.Y(n8557), 
	.A(\ram[159][4] ));
   OAI22X1 U4314 (.Y(n3129), 
	.B1(n8558), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6336));
   INVX1 U4315 (.Y(n8558), 
	.A(\ram[159][3] ));
   OAI22X1 U4316 (.Y(n3128), 
	.B1(n8559), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6338));
   INVX1 U4317 (.Y(n8559), 
	.A(\ram[159][2] ));
   OAI22X1 U4318 (.Y(n3127), 
	.B1(n8560), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6306));
   INVX1 U4319 (.Y(n8560), 
	.A(\ram[159][1] ));
   OAI22X1 U4320 (.Y(n3126), 
	.B1(n8561), 
	.B0(n8545), 
	.A1(n8544), 
	.A0(n6309));
   INVX1 U4321 (.Y(n8561), 
	.A(\ram[159][0] ));
   NOR2BX1 U4322 (.Y(n8545), 
	.B(n8544), 
	.AN(mem_write_en));
   NAND2X1 U4323 (.Y(n8544), 
	.B(n6533), 
	.A(n8562));
   OAI22X1 U4324 (.Y(n3125), 
	.B1(n8565), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6311));
   INVX1 U4325 (.Y(n8565), 
	.A(\ram[158][15] ));
   OAI22X1 U4326 (.Y(n3124), 
	.B1(n8566), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6314));
   INVX1 U4327 (.Y(n8566), 
	.A(\ram[158][14] ));
   OAI22X1 U4328 (.Y(n3123), 
	.B1(n8567), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6316));
   INVX1 U4329 (.Y(n8567), 
	.A(\ram[158][13] ));
   OAI22X1 U4330 (.Y(n3122), 
	.B1(n8568), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6318));
   INVX1 U4331 (.Y(n8568), 
	.A(\ram[158][12] ));
   OAI22X1 U4332 (.Y(n3121), 
	.B1(n8569), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6320));
   INVX1 U4333 (.Y(n8569), 
	.A(\ram[158][11] ));
   OAI22X1 U4334 (.Y(n3120), 
	.B1(n8570), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6322));
   INVX1 U4335 (.Y(n8570), 
	.A(\ram[158][10] ));
   OAI22X1 U4336 (.Y(n3119), 
	.B1(n8571), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6324));
   INVX1 U4337 (.Y(n8571), 
	.A(\ram[158][9] ));
   OAI22X1 U4338 (.Y(n3118), 
	.B1(n8572), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6326));
   INVX1 U4339 (.Y(n8572), 
	.A(\ram[158][8] ));
   OAI22X1 U4340 (.Y(n3117), 
	.B1(n8573), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6328));
   INVX1 U4341 (.Y(n8573), 
	.A(\ram[158][7] ));
   OAI22X1 U4342 (.Y(n3116), 
	.B1(n8574), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6330));
   INVX1 U4343 (.Y(n8574), 
	.A(\ram[158][6] ));
   OAI22X1 U4344 (.Y(n3115), 
	.B1(n8575), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6332));
   INVX1 U4345 (.Y(n8575), 
	.A(\ram[158][5] ));
   OAI22X1 U4346 (.Y(n3114), 
	.B1(n8576), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6334));
   INVX1 U4347 (.Y(n8576), 
	.A(\ram[158][4] ));
   OAI22X1 U4348 (.Y(n3113), 
	.B1(n8577), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6336));
   INVX1 U4349 (.Y(n8577), 
	.A(\ram[158][3] ));
   OAI22X1 U4350 (.Y(n3112), 
	.B1(n8578), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6338));
   INVX1 U4351 (.Y(n8578), 
	.A(\ram[158][2] ));
   OAI22X1 U4352 (.Y(n3111), 
	.B1(n8579), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6306));
   INVX1 U4353 (.Y(n8579), 
	.A(\ram[158][1] ));
   OAI22X1 U4354 (.Y(n3110), 
	.B1(n8580), 
	.B0(n8564), 
	.A1(n8563), 
	.A0(n6309));
   INVX1 U4355 (.Y(n8580), 
	.A(\ram[158][0] ));
   NOR2BX1 U4356 (.Y(n8564), 
	.B(n8563), 
	.AN(mem_write_en));
   NAND2X1 U4357 (.Y(n8563), 
	.B(n6553), 
	.A(n8562));
   OAI22X1 U4358 (.Y(n3109), 
	.B1(n8583), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6311));
   INVX1 U4359 (.Y(n8583), 
	.A(\ram[157][15] ));
   OAI22X1 U4360 (.Y(n3108), 
	.B1(n8584), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6314));
   INVX1 U4361 (.Y(n8584), 
	.A(\ram[157][14] ));
   OAI22X1 U4362 (.Y(n3107), 
	.B1(n8585), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6316));
   INVX1 U4363 (.Y(n8585), 
	.A(\ram[157][13] ));
   OAI22X1 U4364 (.Y(n3106), 
	.B1(n8586), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6318));
   INVX1 U4365 (.Y(n8586), 
	.A(\ram[157][12] ));
   OAI22X1 U4366 (.Y(n3105), 
	.B1(n8587), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6320));
   INVX1 U4367 (.Y(n8587), 
	.A(\ram[157][11] ));
   OAI22X1 U4368 (.Y(n3104), 
	.B1(n8588), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6322));
   INVX1 U4369 (.Y(n8588), 
	.A(\ram[157][10] ));
   OAI22X1 U4370 (.Y(n3103), 
	.B1(n8589), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6324));
   INVX1 U4371 (.Y(n8589), 
	.A(\ram[157][9] ));
   OAI22X1 U4372 (.Y(n3102), 
	.B1(n8590), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6326));
   INVX1 U4373 (.Y(n8590), 
	.A(\ram[157][8] ));
   OAI22X1 U4374 (.Y(n3101), 
	.B1(n8591), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6328));
   INVX1 U4375 (.Y(n8591), 
	.A(\ram[157][7] ));
   OAI22X1 U4376 (.Y(n3100), 
	.B1(n8592), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6330));
   INVX1 U4377 (.Y(n8592), 
	.A(\ram[157][6] ));
   OAI22X1 U4378 (.Y(n3099), 
	.B1(n8593), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6332));
   INVX1 U4379 (.Y(n8593), 
	.A(\ram[157][5] ));
   OAI22X1 U4380 (.Y(n3098), 
	.B1(n8594), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6334));
   INVX1 U4381 (.Y(n8594), 
	.A(\ram[157][4] ));
   OAI22X1 U4382 (.Y(n3097), 
	.B1(n8595), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6336));
   INVX1 U4383 (.Y(n8595), 
	.A(\ram[157][3] ));
   OAI22X1 U4384 (.Y(n3096), 
	.B1(n8596), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6338));
   INVX1 U4385 (.Y(n8596), 
	.A(\ram[157][2] ));
   OAI22X1 U4386 (.Y(n3095), 
	.B1(n8597), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6306));
   INVX1 U4387 (.Y(n8597), 
	.A(\ram[157][1] ));
   OAI22X1 U4388 (.Y(n3094), 
	.B1(n8598), 
	.B0(n8582), 
	.A1(n8581), 
	.A0(n6309));
   INVX1 U4389 (.Y(n8598), 
	.A(\ram[157][0] ));
   NOR2BX1 U4390 (.Y(n8582), 
	.B(n8581), 
	.AN(mem_write_en));
   NAND2X1 U4391 (.Y(n8581), 
	.B(n6572), 
	.A(n8562));
   OAI22X1 U4392 (.Y(n3093), 
	.B1(n8601), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6311));
   INVX1 U4393 (.Y(n8601), 
	.A(\ram[156][15] ));
   OAI22X1 U4394 (.Y(n3092), 
	.B1(n8602), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6314));
   INVX1 U4395 (.Y(n8602), 
	.A(\ram[156][14] ));
   OAI22X1 U4396 (.Y(n3091), 
	.B1(n8603), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6316));
   INVX1 U4397 (.Y(n8603), 
	.A(\ram[156][13] ));
   OAI22X1 U4398 (.Y(n3090), 
	.B1(n8604), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6318));
   INVX1 U4399 (.Y(n8604), 
	.A(\ram[156][12] ));
   OAI22X1 U4400 (.Y(n3089), 
	.B1(n8605), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6320));
   INVX1 U4401 (.Y(n8605), 
	.A(\ram[156][11] ));
   OAI22X1 U4402 (.Y(n3088), 
	.B1(n8606), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6322));
   INVX1 U4403 (.Y(n8606), 
	.A(\ram[156][10] ));
   OAI22X1 U4404 (.Y(n3087), 
	.B1(n8607), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6324));
   INVX1 U4405 (.Y(n8607), 
	.A(\ram[156][9] ));
   OAI22X1 U4406 (.Y(n3086), 
	.B1(n8608), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6326));
   INVX1 U4407 (.Y(n8608), 
	.A(\ram[156][8] ));
   OAI22X1 U4408 (.Y(n3085), 
	.B1(n8609), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6328));
   INVX1 U4409 (.Y(n8609), 
	.A(\ram[156][7] ));
   OAI22X1 U4410 (.Y(n3084), 
	.B1(n8610), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6330));
   INVX1 U4411 (.Y(n8610), 
	.A(\ram[156][6] ));
   OAI22X1 U4412 (.Y(n3083), 
	.B1(n8611), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6332));
   INVX1 U4413 (.Y(n8611), 
	.A(\ram[156][5] ));
   OAI22X1 U4414 (.Y(n3082), 
	.B1(n8612), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6334));
   INVX1 U4415 (.Y(n8612), 
	.A(\ram[156][4] ));
   OAI22X1 U4416 (.Y(n3081), 
	.B1(n8613), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6336));
   INVX1 U4417 (.Y(n8613), 
	.A(\ram[156][3] ));
   OAI22X1 U4418 (.Y(n3080), 
	.B1(n8614), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6338));
   INVX1 U4419 (.Y(n8614), 
	.A(\ram[156][2] ));
   OAI22X1 U4420 (.Y(n3079), 
	.B1(n8615), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6306));
   INVX1 U4421 (.Y(n8615), 
	.A(\ram[156][1] ));
   OAI22X1 U4422 (.Y(n3078), 
	.B1(n8616), 
	.B0(n8600), 
	.A1(n8599), 
	.A0(n6309));
   INVX1 U4423 (.Y(n8616), 
	.A(\ram[156][0] ));
   NOR2BX1 U4424 (.Y(n8600), 
	.B(n8599), 
	.AN(mem_write_en));
   NAND2X1 U4425 (.Y(n8599), 
	.B(n6591), 
	.A(n8562));
   OAI22X1 U4426 (.Y(n3077), 
	.B1(n8619), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6311));
   INVX1 U4427 (.Y(n8619), 
	.A(\ram[155][15] ));
   OAI22X1 U4428 (.Y(n3076), 
	.B1(n8620), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6314));
   INVX1 U4429 (.Y(n8620), 
	.A(\ram[155][14] ));
   OAI22X1 U4430 (.Y(n3075), 
	.B1(n8621), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6316));
   INVX1 U4431 (.Y(n8621), 
	.A(\ram[155][13] ));
   OAI22X1 U4432 (.Y(n3074), 
	.B1(n8622), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6318));
   INVX1 U4433 (.Y(n8622), 
	.A(\ram[155][12] ));
   OAI22X1 U4434 (.Y(n3073), 
	.B1(n8623), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6320));
   INVX1 U4435 (.Y(n8623), 
	.A(\ram[155][11] ));
   OAI22X1 U4436 (.Y(n3072), 
	.B1(n8624), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6322));
   INVX1 U4437 (.Y(n8624), 
	.A(\ram[155][10] ));
   OAI22X1 U4438 (.Y(n3071), 
	.B1(n8625), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6324));
   INVX1 U4439 (.Y(n8625), 
	.A(\ram[155][9] ));
   OAI22X1 U4440 (.Y(n3070), 
	.B1(n8626), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6326));
   INVX1 U4441 (.Y(n8626), 
	.A(\ram[155][8] ));
   OAI22X1 U4442 (.Y(n3069), 
	.B1(n8627), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6328));
   INVX1 U4443 (.Y(n8627), 
	.A(\ram[155][7] ));
   OAI22X1 U4444 (.Y(n3068), 
	.B1(n8628), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6330));
   INVX1 U4445 (.Y(n8628), 
	.A(\ram[155][6] ));
   OAI22X1 U4446 (.Y(n3067), 
	.B1(n8629), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6332));
   INVX1 U4447 (.Y(n8629), 
	.A(\ram[155][5] ));
   OAI22X1 U4448 (.Y(n3066), 
	.B1(n8630), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6334));
   INVX1 U4449 (.Y(n8630), 
	.A(\ram[155][4] ));
   OAI22X1 U4450 (.Y(n3065), 
	.B1(n8631), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6336));
   INVX1 U4451 (.Y(n8631), 
	.A(\ram[155][3] ));
   OAI22X1 U4452 (.Y(n3064), 
	.B1(n8632), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6338));
   INVX1 U4453 (.Y(n8632), 
	.A(\ram[155][2] ));
   OAI22X1 U4454 (.Y(n3063), 
	.B1(n8633), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6306));
   INVX1 U4455 (.Y(n8633), 
	.A(\ram[155][1] ));
   OAI22X1 U4456 (.Y(n3062), 
	.B1(n8634), 
	.B0(n8618), 
	.A1(n8617), 
	.A0(n6309));
   INVX1 U4457 (.Y(n8634), 
	.A(\ram[155][0] ));
   NOR2BX1 U4458 (.Y(n8618), 
	.B(n8617), 
	.AN(mem_write_en));
   NAND2X1 U4459 (.Y(n8617), 
	.B(n6610), 
	.A(n8562));
   OAI22X1 U4460 (.Y(n3061), 
	.B1(n8637), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6311));
   INVX1 U4461 (.Y(n8637), 
	.A(\ram[154][15] ));
   OAI22X1 U4462 (.Y(n3060), 
	.B1(n8638), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6314));
   INVX1 U4463 (.Y(n8638), 
	.A(\ram[154][14] ));
   OAI22X1 U4464 (.Y(n3059), 
	.B1(n8639), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6316));
   INVX1 U4465 (.Y(n8639), 
	.A(\ram[154][13] ));
   OAI22X1 U4466 (.Y(n3058), 
	.B1(n8640), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6318));
   INVX1 U4467 (.Y(n8640), 
	.A(\ram[154][12] ));
   OAI22X1 U4468 (.Y(n3057), 
	.B1(n8641), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6320));
   INVX1 U4469 (.Y(n8641), 
	.A(\ram[154][11] ));
   OAI22X1 U4470 (.Y(n3056), 
	.B1(n8642), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6322));
   INVX1 U4471 (.Y(n8642), 
	.A(\ram[154][10] ));
   OAI22X1 U4472 (.Y(n3055), 
	.B1(n8643), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6324));
   INVX1 U4473 (.Y(n8643), 
	.A(\ram[154][9] ));
   OAI22X1 U4474 (.Y(n3054), 
	.B1(n8644), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6326));
   INVX1 U4475 (.Y(n8644), 
	.A(\ram[154][8] ));
   OAI22X1 U4476 (.Y(n3053), 
	.B1(n8645), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6328));
   INVX1 U4477 (.Y(n8645), 
	.A(\ram[154][7] ));
   OAI22X1 U4478 (.Y(n3052), 
	.B1(n8646), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6330));
   INVX1 U4479 (.Y(n8646), 
	.A(\ram[154][6] ));
   OAI22X1 U4480 (.Y(n3051), 
	.B1(n8647), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6332));
   INVX1 U4481 (.Y(n8647), 
	.A(\ram[154][5] ));
   OAI22X1 U4482 (.Y(n3050), 
	.B1(n8648), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6334));
   INVX1 U4483 (.Y(n8648), 
	.A(\ram[154][4] ));
   OAI22X1 U4484 (.Y(n3049), 
	.B1(n8649), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6336));
   INVX1 U4485 (.Y(n8649), 
	.A(\ram[154][3] ));
   OAI22X1 U4486 (.Y(n3048), 
	.B1(n8650), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6338));
   INVX1 U4487 (.Y(n8650), 
	.A(\ram[154][2] ));
   OAI22X1 U4488 (.Y(n3047), 
	.B1(n8651), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6306));
   INVX1 U4489 (.Y(n8651), 
	.A(\ram[154][1] ));
   OAI22X1 U4490 (.Y(n3046), 
	.B1(n8652), 
	.B0(n8636), 
	.A1(n8635), 
	.A0(n6309));
   INVX1 U4491 (.Y(n8652), 
	.A(\ram[154][0] ));
   NOR2BX1 U4492 (.Y(n8636), 
	.B(n8635), 
	.AN(mem_write_en));
   NAND2X1 U4493 (.Y(n8635), 
	.B(n6629), 
	.A(n8562));
   OAI22X1 U4494 (.Y(n3045), 
	.B1(n8655), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6311));
   INVX1 U4495 (.Y(n8655), 
	.A(\ram[153][15] ));
   OAI22X1 U4496 (.Y(n3044), 
	.B1(n8656), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6314));
   INVX1 U4497 (.Y(n8656), 
	.A(\ram[153][14] ));
   OAI22X1 U4498 (.Y(n3043), 
	.B1(n8657), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6316));
   INVX1 U4499 (.Y(n8657), 
	.A(\ram[153][13] ));
   OAI22X1 U4500 (.Y(n3042), 
	.B1(n8658), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6318));
   INVX1 U4501 (.Y(n8658), 
	.A(\ram[153][12] ));
   OAI22X1 U4502 (.Y(n3041), 
	.B1(n8659), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6320));
   INVX1 U4503 (.Y(n8659), 
	.A(\ram[153][11] ));
   OAI22X1 U4504 (.Y(n3040), 
	.B1(n8660), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6322));
   INVX1 U4505 (.Y(n8660), 
	.A(\ram[153][10] ));
   OAI22X1 U4506 (.Y(n3039), 
	.B1(n8661), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6324));
   INVX1 U4507 (.Y(n8661), 
	.A(\ram[153][9] ));
   OAI22X1 U4508 (.Y(n3038), 
	.B1(n8662), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6326));
   INVX1 U4509 (.Y(n8662), 
	.A(\ram[153][8] ));
   OAI22X1 U4510 (.Y(n3037), 
	.B1(n8663), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6328));
   INVX1 U4511 (.Y(n8663), 
	.A(\ram[153][7] ));
   OAI22X1 U4512 (.Y(n3036), 
	.B1(n8664), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6330));
   INVX1 U4513 (.Y(n8664), 
	.A(\ram[153][6] ));
   OAI22X1 U4514 (.Y(n3035), 
	.B1(n8665), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6332));
   INVX1 U4515 (.Y(n8665), 
	.A(\ram[153][5] ));
   OAI22X1 U4516 (.Y(n3034), 
	.B1(n8666), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6334));
   INVX1 U4517 (.Y(n8666), 
	.A(\ram[153][4] ));
   OAI22X1 U4518 (.Y(n3033), 
	.B1(n8667), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6336));
   INVX1 U4519 (.Y(n8667), 
	.A(\ram[153][3] ));
   OAI22X1 U4520 (.Y(n3032), 
	.B1(n8668), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6338));
   INVX1 U4521 (.Y(n8668), 
	.A(\ram[153][2] ));
   OAI22X1 U4522 (.Y(n3031), 
	.B1(n8669), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6306));
   INVX1 U4523 (.Y(n8669), 
	.A(\ram[153][1] ));
   OAI22X1 U4524 (.Y(n3030), 
	.B1(n8670), 
	.B0(n8654), 
	.A1(n8653), 
	.A0(n6309));
   INVX1 U4525 (.Y(n8670), 
	.A(\ram[153][0] ));
   NOR2BX1 U4526 (.Y(n8654), 
	.B(n8653), 
	.AN(mem_write_en));
   NAND2X1 U4527 (.Y(n8653), 
	.B(n6342), 
	.A(n8562));
   OAI22X1 U4528 (.Y(n3029), 
	.B1(n8673), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6311));
   INVX1 U4529 (.Y(n8673), 
	.A(\ram[152][15] ));
   OAI22X1 U4530 (.Y(n3028), 
	.B1(n8674), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6314));
   INVX1 U4531 (.Y(n8674), 
	.A(\ram[152][14] ));
   OAI22X1 U4532 (.Y(n3027), 
	.B1(n8675), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6316));
   INVX1 U4533 (.Y(n8675), 
	.A(\ram[152][13] ));
   OAI22X1 U4534 (.Y(n3026), 
	.B1(n8676), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6318));
   INVX1 U4535 (.Y(n8676), 
	.A(\ram[152][12] ));
   OAI22X1 U4536 (.Y(n3025), 
	.B1(n8677), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6320));
   INVX1 U4537 (.Y(n8677), 
	.A(\ram[152][11] ));
   OAI22X1 U4538 (.Y(n3024), 
	.B1(n8678), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6322));
   INVX1 U4539 (.Y(n8678), 
	.A(\ram[152][10] ));
   OAI22X1 U4540 (.Y(n3023), 
	.B1(n8679), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6324));
   INVX1 U4541 (.Y(n8679), 
	.A(\ram[152][9] ));
   OAI22X1 U4542 (.Y(n3022), 
	.B1(n8680), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6326));
   INVX1 U4543 (.Y(n8680), 
	.A(\ram[152][8] ));
   OAI22X1 U4544 (.Y(n3021), 
	.B1(n8681), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6328));
   INVX1 U4545 (.Y(n8681), 
	.A(\ram[152][7] ));
   OAI22X1 U4546 (.Y(n3020), 
	.B1(n8682), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6330));
   INVX1 U4547 (.Y(n8682), 
	.A(\ram[152][6] ));
   OAI22X1 U4548 (.Y(n3019), 
	.B1(n8683), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6332));
   INVX1 U4549 (.Y(n8683), 
	.A(\ram[152][5] ));
   OAI22X1 U4550 (.Y(n3018), 
	.B1(n8684), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6334));
   INVX1 U4551 (.Y(n8684), 
	.A(\ram[152][4] ));
   OAI22X1 U4552 (.Y(n3017), 
	.B1(n8685), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6336));
   INVX1 U4553 (.Y(n8685), 
	.A(\ram[152][3] ));
   OAI22X1 U4554 (.Y(n3016), 
	.B1(n8686), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6338));
   INVX1 U4555 (.Y(n8686), 
	.A(\ram[152][2] ));
   OAI22X1 U4556 (.Y(n3015), 
	.B1(n8687), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6306));
   INVX1 U4557 (.Y(n8687), 
	.A(\ram[152][1] ));
   OAI22X1 U4558 (.Y(n3014), 
	.B1(n8688), 
	.B0(n8672), 
	.A1(n8671), 
	.A0(n6309));
   INVX1 U4559 (.Y(n8688), 
	.A(\ram[152][0] ));
   NOR2BX1 U4560 (.Y(n8672), 
	.B(n8671), 
	.AN(mem_write_en));
   NAND2X1 U4561 (.Y(n8671), 
	.B(n6362), 
	.A(n8562));
   OAI22X1 U4562 (.Y(n3013), 
	.B1(n8691), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6311));
   INVX1 U4563 (.Y(n8691), 
	.A(\ram[151][15] ));
   OAI22X1 U4564 (.Y(n3012), 
	.B1(n8692), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6314));
   INVX1 U4565 (.Y(n8692), 
	.A(\ram[151][14] ));
   OAI22X1 U4566 (.Y(n3011), 
	.B1(n8693), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6316));
   INVX1 U4567 (.Y(n8693), 
	.A(\ram[151][13] ));
   OAI22X1 U4568 (.Y(n3010), 
	.B1(n8694), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6318));
   INVX1 U4569 (.Y(n8694), 
	.A(\ram[151][12] ));
   OAI22X1 U4570 (.Y(n3009), 
	.B1(n8695), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6320));
   INVX1 U4571 (.Y(n8695), 
	.A(\ram[151][11] ));
   OAI22X1 U4572 (.Y(n3008), 
	.B1(n8696), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6322));
   INVX1 U4573 (.Y(n8696), 
	.A(\ram[151][10] ));
   OAI22X1 U4574 (.Y(n3007), 
	.B1(n8697), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6324));
   INVX1 U4575 (.Y(n8697), 
	.A(\ram[151][9] ));
   OAI22X1 U4576 (.Y(n3006), 
	.B1(n8698), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6326));
   INVX1 U4577 (.Y(n8698), 
	.A(\ram[151][8] ));
   OAI22X1 U4578 (.Y(n3005), 
	.B1(n8699), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6328));
   INVX1 U4579 (.Y(n8699), 
	.A(\ram[151][7] ));
   OAI22X1 U4580 (.Y(n3004), 
	.B1(n8700), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6330));
   INVX1 U4581 (.Y(n8700), 
	.A(\ram[151][6] ));
   OAI22X1 U4582 (.Y(n3003), 
	.B1(n8701), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6332));
   INVX1 U4583 (.Y(n8701), 
	.A(\ram[151][5] ));
   OAI22X1 U4584 (.Y(n3002), 
	.B1(n8702), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6334));
   INVX1 U4585 (.Y(n8702), 
	.A(\ram[151][4] ));
   OAI22X1 U4586 (.Y(n3001), 
	.B1(n8703), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6336));
   INVX1 U4587 (.Y(n8703), 
	.A(\ram[151][3] ));
   OAI22X1 U4588 (.Y(n3000), 
	.B1(n8704), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6338));
   INVX1 U4589 (.Y(n8704), 
	.A(\ram[151][2] ));
   OAI22X1 U4590 (.Y(n2999), 
	.B1(n8705), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6306));
   INVX1 U4591 (.Y(n8705), 
	.A(\ram[151][1] ));
   OAI22X1 U4592 (.Y(n2998), 
	.B1(n8706), 
	.B0(n8690), 
	.A1(n8689), 
	.A0(n6309));
   INVX1 U4593 (.Y(n8706), 
	.A(\ram[151][0] ));
   NOR2BX1 U4594 (.Y(n8690), 
	.B(n8689), 
	.AN(mem_write_en));
   NAND2X1 U4595 (.Y(n8689), 
	.B(n6381), 
	.A(n8562));
   OAI22X1 U4596 (.Y(n2997), 
	.B1(n8709), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6311));
   INVX1 U4597 (.Y(n8709), 
	.A(\ram[150][15] ));
   OAI22X1 U4598 (.Y(n2996), 
	.B1(n8710), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6314));
   INVX1 U4599 (.Y(n8710), 
	.A(\ram[150][14] ));
   OAI22X1 U4600 (.Y(n2995), 
	.B1(n8711), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6316));
   INVX1 U4601 (.Y(n8711), 
	.A(\ram[150][13] ));
   OAI22X1 U4602 (.Y(n2994), 
	.B1(n8712), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6318));
   INVX1 U4603 (.Y(n8712), 
	.A(\ram[150][12] ));
   OAI22X1 U4604 (.Y(n2993), 
	.B1(n8713), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6320));
   INVX1 U4605 (.Y(n8713), 
	.A(\ram[150][11] ));
   OAI22X1 U4606 (.Y(n2992), 
	.B1(n8714), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6322));
   INVX1 U4607 (.Y(n8714), 
	.A(\ram[150][10] ));
   OAI22X1 U4608 (.Y(n2991), 
	.B1(n8715), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6324));
   INVX1 U4609 (.Y(n8715), 
	.A(\ram[150][9] ));
   OAI22X1 U4610 (.Y(n2990), 
	.B1(n8716), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6326));
   INVX1 U4611 (.Y(n8716), 
	.A(\ram[150][8] ));
   OAI22X1 U4612 (.Y(n2989), 
	.B1(n8717), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6328));
   INVX1 U4613 (.Y(n8717), 
	.A(\ram[150][7] ));
   OAI22X1 U4614 (.Y(n2988), 
	.B1(n8718), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6330));
   INVX1 U4615 (.Y(n8718), 
	.A(\ram[150][6] ));
   OAI22X1 U4616 (.Y(n2987), 
	.B1(n8719), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6332));
   INVX1 U4617 (.Y(n8719), 
	.A(\ram[150][5] ));
   OAI22X1 U4618 (.Y(n2986), 
	.B1(n8720), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6334));
   INVX1 U4619 (.Y(n8720), 
	.A(\ram[150][4] ));
   OAI22X1 U4620 (.Y(n2985), 
	.B1(n8721), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6336));
   INVX1 U4621 (.Y(n8721), 
	.A(\ram[150][3] ));
   OAI22X1 U4622 (.Y(n2984), 
	.B1(n8722), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6338));
   INVX1 U4623 (.Y(n8722), 
	.A(\ram[150][2] ));
   OAI22X1 U4624 (.Y(n2983), 
	.B1(n8723), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6306));
   INVX1 U4625 (.Y(n8723), 
	.A(\ram[150][1] ));
   OAI22X1 U4626 (.Y(n2982), 
	.B1(n8724), 
	.B0(n8708), 
	.A1(n8707), 
	.A0(n6309));
   INVX1 U4627 (.Y(n8724), 
	.A(\ram[150][0] ));
   NOR2BX1 U4628 (.Y(n8708), 
	.B(n8707), 
	.AN(mem_write_en));
   NAND2X1 U4629 (.Y(n8707), 
	.B(n6400), 
	.A(n8562));
   OAI22X1 U4630 (.Y(n2981), 
	.B1(n8727), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6311));
   INVX1 U4631 (.Y(n8727), 
	.A(\ram[149][15] ));
   OAI22X1 U4632 (.Y(n2980), 
	.B1(n8728), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6314));
   INVX1 U4633 (.Y(n8728), 
	.A(\ram[149][14] ));
   OAI22X1 U4634 (.Y(n2979), 
	.B1(n8729), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6316));
   INVX1 U4635 (.Y(n8729), 
	.A(\ram[149][13] ));
   OAI22X1 U4636 (.Y(n2978), 
	.B1(n8730), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6318));
   INVX1 U4637 (.Y(n8730), 
	.A(\ram[149][12] ));
   OAI22X1 U4638 (.Y(n2977), 
	.B1(n8731), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6320));
   INVX1 U4639 (.Y(n8731), 
	.A(\ram[149][11] ));
   OAI22X1 U4640 (.Y(n2976), 
	.B1(n8732), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6322));
   INVX1 U4641 (.Y(n8732), 
	.A(\ram[149][10] ));
   OAI22X1 U4642 (.Y(n2975), 
	.B1(n8733), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6324));
   INVX1 U4643 (.Y(n8733), 
	.A(\ram[149][9] ));
   OAI22X1 U4644 (.Y(n2974), 
	.B1(n8734), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6326));
   INVX1 U4645 (.Y(n8734), 
	.A(\ram[149][8] ));
   OAI22X1 U4646 (.Y(n2973), 
	.B1(n8735), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6328));
   INVX1 U4647 (.Y(n8735), 
	.A(\ram[149][7] ));
   OAI22X1 U4648 (.Y(n2972), 
	.B1(n8736), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6330));
   INVX1 U4649 (.Y(n8736), 
	.A(\ram[149][6] ));
   OAI22X1 U4650 (.Y(n2971), 
	.B1(n8737), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6332));
   INVX1 U4651 (.Y(n8737), 
	.A(\ram[149][5] ));
   OAI22X1 U4652 (.Y(n2970), 
	.B1(n8738), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6334));
   INVX1 U4653 (.Y(n8738), 
	.A(\ram[149][4] ));
   OAI22X1 U4654 (.Y(n2969), 
	.B1(n8739), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6336));
   INVX1 U4655 (.Y(n8739), 
	.A(\ram[149][3] ));
   OAI22X1 U4656 (.Y(n2968), 
	.B1(n8740), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6338));
   INVX1 U4657 (.Y(n8740), 
	.A(\ram[149][2] ));
   OAI22X1 U4658 (.Y(n2967), 
	.B1(n8741), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6306));
   INVX1 U4659 (.Y(n8741), 
	.A(\ram[149][1] ));
   OAI22X1 U4660 (.Y(n2966), 
	.B1(n8742), 
	.B0(n8726), 
	.A1(n8725), 
	.A0(n6309));
   INVX1 U4661 (.Y(n8742), 
	.A(\ram[149][0] ));
   NOR2BX1 U4662 (.Y(n8726), 
	.B(n8725), 
	.AN(mem_write_en));
   NAND2X1 U4663 (.Y(n8725), 
	.B(n6419), 
	.A(n8562));
   OAI22X1 U4664 (.Y(n2965), 
	.B1(n8745), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6311));
   INVX1 U4665 (.Y(n8745), 
	.A(\ram[148][15] ));
   OAI22X1 U4666 (.Y(n2964), 
	.B1(n8746), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6314));
   INVX1 U4667 (.Y(n8746), 
	.A(\ram[148][14] ));
   OAI22X1 U4668 (.Y(n2963), 
	.B1(n8747), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6316));
   INVX1 U4669 (.Y(n8747), 
	.A(\ram[148][13] ));
   OAI22X1 U4670 (.Y(n2962), 
	.B1(n8748), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6318));
   INVX1 U4671 (.Y(n8748), 
	.A(\ram[148][12] ));
   OAI22X1 U4672 (.Y(n2961), 
	.B1(n8749), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6320));
   INVX1 U4673 (.Y(n8749), 
	.A(\ram[148][11] ));
   OAI22X1 U4674 (.Y(n2960), 
	.B1(n8750), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6322));
   INVX1 U4675 (.Y(n8750), 
	.A(\ram[148][10] ));
   OAI22X1 U4676 (.Y(n2959), 
	.B1(n8751), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6324));
   INVX1 U4677 (.Y(n8751), 
	.A(\ram[148][9] ));
   OAI22X1 U4678 (.Y(n2958), 
	.B1(n8752), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6326));
   INVX1 U4679 (.Y(n8752), 
	.A(\ram[148][8] ));
   OAI22X1 U4680 (.Y(n2957), 
	.B1(n8753), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6328));
   INVX1 U4681 (.Y(n8753), 
	.A(\ram[148][7] ));
   OAI22X1 U4682 (.Y(n2956), 
	.B1(n8754), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6330));
   INVX1 U4683 (.Y(n8754), 
	.A(\ram[148][6] ));
   OAI22X1 U4684 (.Y(n2955), 
	.B1(n8755), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6332));
   INVX1 U4685 (.Y(n8755), 
	.A(\ram[148][5] ));
   OAI22X1 U4686 (.Y(n2954), 
	.B1(n8756), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6334));
   INVX1 U4687 (.Y(n8756), 
	.A(\ram[148][4] ));
   OAI22X1 U4688 (.Y(n2953), 
	.B1(n8757), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6336));
   INVX1 U4689 (.Y(n8757), 
	.A(\ram[148][3] ));
   OAI22X1 U4690 (.Y(n2952), 
	.B1(n8758), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6338));
   INVX1 U4691 (.Y(n8758), 
	.A(\ram[148][2] ));
   OAI22X1 U4692 (.Y(n2951), 
	.B1(n8759), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6306));
   INVX1 U4693 (.Y(n8759), 
	.A(\ram[148][1] ));
   OAI22X1 U4694 (.Y(n2950), 
	.B1(n8760), 
	.B0(n8744), 
	.A1(n8743), 
	.A0(n6309));
   INVX1 U4695 (.Y(n8760), 
	.A(\ram[148][0] ));
   NOR2BX1 U4696 (.Y(n8744), 
	.B(n8743), 
	.AN(mem_write_en));
   NAND2X1 U4697 (.Y(n8743), 
	.B(n6438), 
	.A(n8562));
   OAI22X1 U4698 (.Y(n2949), 
	.B1(n8763), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6311));
   INVX1 U4699 (.Y(n8763), 
	.A(\ram[147][15] ));
   OAI22X1 U4700 (.Y(n2948), 
	.B1(n8764), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6314));
   INVX1 U4701 (.Y(n8764), 
	.A(\ram[147][14] ));
   OAI22X1 U4702 (.Y(n2947), 
	.B1(n8765), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6316));
   INVX1 U4703 (.Y(n8765), 
	.A(\ram[147][13] ));
   OAI22X1 U4704 (.Y(n2946), 
	.B1(n8766), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6318));
   INVX1 U4705 (.Y(n8766), 
	.A(\ram[147][12] ));
   OAI22X1 U4706 (.Y(n2945), 
	.B1(n8767), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6320));
   INVX1 U4707 (.Y(n8767), 
	.A(\ram[147][11] ));
   OAI22X1 U4708 (.Y(n2944), 
	.B1(n8768), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6322));
   INVX1 U4709 (.Y(n8768), 
	.A(\ram[147][10] ));
   OAI22X1 U4710 (.Y(n2943), 
	.B1(n8769), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6324));
   INVX1 U4711 (.Y(n8769), 
	.A(\ram[147][9] ));
   OAI22X1 U4712 (.Y(n2942), 
	.B1(n8770), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6326));
   INVX1 U4713 (.Y(n8770), 
	.A(\ram[147][8] ));
   OAI22X1 U4714 (.Y(n2941), 
	.B1(n8771), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6328));
   INVX1 U4715 (.Y(n8771), 
	.A(\ram[147][7] ));
   OAI22X1 U4716 (.Y(n2940), 
	.B1(n8772), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6330));
   INVX1 U4717 (.Y(n8772), 
	.A(\ram[147][6] ));
   OAI22X1 U4718 (.Y(n2939), 
	.B1(n8773), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6332));
   INVX1 U4719 (.Y(n8773), 
	.A(\ram[147][5] ));
   OAI22X1 U4720 (.Y(n2938), 
	.B1(n8774), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6334));
   INVX1 U4721 (.Y(n8774), 
	.A(\ram[147][4] ));
   OAI22X1 U4722 (.Y(n2937), 
	.B1(n8775), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6336));
   INVX1 U4723 (.Y(n8775), 
	.A(\ram[147][3] ));
   OAI22X1 U4724 (.Y(n2936), 
	.B1(n8776), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6338));
   INVX1 U4725 (.Y(n8776), 
	.A(\ram[147][2] ));
   OAI22X1 U4726 (.Y(n2935), 
	.B1(n8777), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6306));
   INVX1 U4727 (.Y(n8777), 
	.A(\ram[147][1] ));
   OAI22X1 U4728 (.Y(n2934), 
	.B1(n8778), 
	.B0(n8762), 
	.A1(n8761), 
	.A0(n6309));
   INVX1 U4729 (.Y(n8778), 
	.A(\ram[147][0] ));
   NOR2BX1 U4730 (.Y(n8762), 
	.B(n8761), 
	.AN(mem_write_en));
   NAND2X1 U4731 (.Y(n8761), 
	.B(n6457), 
	.A(n8562));
   OAI22X1 U4732 (.Y(n2933), 
	.B1(n8781), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6311));
   INVX1 U4733 (.Y(n8781), 
	.A(\ram[146][15] ));
   OAI22X1 U4734 (.Y(n2932), 
	.B1(n8782), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6314));
   INVX1 U4735 (.Y(n8782), 
	.A(\ram[146][14] ));
   OAI22X1 U4736 (.Y(n2931), 
	.B1(n8783), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6316));
   INVX1 U4737 (.Y(n8783), 
	.A(\ram[146][13] ));
   OAI22X1 U4738 (.Y(n2930), 
	.B1(n8784), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6318));
   INVX1 U4739 (.Y(n8784), 
	.A(\ram[146][12] ));
   OAI22X1 U4740 (.Y(n2929), 
	.B1(n8785), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6320));
   INVX1 U4741 (.Y(n8785), 
	.A(\ram[146][11] ));
   OAI22X1 U4742 (.Y(n2928), 
	.B1(n8786), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6322));
   INVX1 U4743 (.Y(n8786), 
	.A(\ram[146][10] ));
   OAI22X1 U4744 (.Y(n2927), 
	.B1(n8787), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6324));
   INVX1 U4745 (.Y(n8787), 
	.A(\ram[146][9] ));
   OAI22X1 U4746 (.Y(n2926), 
	.B1(n8788), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6326));
   INVX1 U4747 (.Y(n8788), 
	.A(\ram[146][8] ));
   OAI22X1 U4748 (.Y(n2925), 
	.B1(n8789), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6328));
   INVX1 U4749 (.Y(n8789), 
	.A(\ram[146][7] ));
   OAI22X1 U4750 (.Y(n2924), 
	.B1(n8790), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6330));
   INVX1 U4751 (.Y(n8790), 
	.A(\ram[146][6] ));
   OAI22X1 U4752 (.Y(n2923), 
	.B1(n8791), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6332));
   INVX1 U4753 (.Y(n8791), 
	.A(\ram[146][5] ));
   OAI22X1 U4754 (.Y(n2922), 
	.B1(n8792), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6334));
   INVX1 U4755 (.Y(n8792), 
	.A(\ram[146][4] ));
   OAI22X1 U4756 (.Y(n2921), 
	.B1(n8793), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6336));
   INVX1 U4757 (.Y(n8793), 
	.A(\ram[146][3] ));
   OAI22X1 U4758 (.Y(n2920), 
	.B1(n8794), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6338));
   INVX1 U4759 (.Y(n8794), 
	.A(\ram[146][2] ));
   OAI22X1 U4760 (.Y(n2919), 
	.B1(n8795), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6306));
   INVX1 U4761 (.Y(n8795), 
	.A(\ram[146][1] ));
   OAI22X1 U4762 (.Y(n2918), 
	.B1(n8796), 
	.B0(n8780), 
	.A1(n8779), 
	.A0(n6309));
   INVX1 U4763 (.Y(n8796), 
	.A(\ram[146][0] ));
   NOR2BX1 U4764 (.Y(n8780), 
	.B(n8779), 
	.AN(mem_write_en));
   NAND2X1 U4765 (.Y(n8779), 
	.B(n6476), 
	.A(n8562));
   OAI22X1 U4766 (.Y(n2917), 
	.B1(n8799), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6311));
   INVX1 U4767 (.Y(n8799), 
	.A(\ram[145][15] ));
   OAI22X1 U4768 (.Y(n2916), 
	.B1(n8800), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6314));
   INVX1 U4769 (.Y(n8800), 
	.A(\ram[145][14] ));
   OAI22X1 U4770 (.Y(n2915), 
	.B1(n8801), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6316));
   INVX1 U4771 (.Y(n8801), 
	.A(\ram[145][13] ));
   OAI22X1 U4772 (.Y(n2914), 
	.B1(n8802), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6318));
   INVX1 U4773 (.Y(n8802), 
	.A(\ram[145][12] ));
   OAI22X1 U4774 (.Y(n2913), 
	.B1(n8803), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6320));
   INVX1 U4775 (.Y(n8803), 
	.A(\ram[145][11] ));
   OAI22X1 U4776 (.Y(n2912), 
	.B1(n8804), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6322));
   INVX1 U4777 (.Y(n8804), 
	.A(\ram[145][10] ));
   OAI22X1 U4778 (.Y(n2911), 
	.B1(n8805), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6324));
   INVX1 U4779 (.Y(n8805), 
	.A(\ram[145][9] ));
   OAI22X1 U4780 (.Y(n2910), 
	.B1(n8806), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6326));
   INVX1 U4781 (.Y(n8806), 
	.A(\ram[145][8] ));
   OAI22X1 U4782 (.Y(n2909), 
	.B1(n8807), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6328));
   INVX1 U4783 (.Y(n8807), 
	.A(\ram[145][7] ));
   OAI22X1 U4784 (.Y(n2908), 
	.B1(n8808), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6330));
   INVX1 U4785 (.Y(n8808), 
	.A(\ram[145][6] ));
   OAI22X1 U4786 (.Y(n2907), 
	.B1(n8809), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6332));
   INVX1 U4787 (.Y(n8809), 
	.A(\ram[145][5] ));
   OAI22X1 U4788 (.Y(n2906), 
	.B1(n8810), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6334));
   INVX1 U4789 (.Y(n8810), 
	.A(\ram[145][4] ));
   OAI22X1 U4790 (.Y(n2905), 
	.B1(n8811), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6336));
   INVX1 U4791 (.Y(n8811), 
	.A(\ram[145][3] ));
   OAI22X1 U4792 (.Y(n2904), 
	.B1(n8812), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6338));
   INVX1 U4793 (.Y(n8812), 
	.A(\ram[145][2] ));
   OAI22X1 U4794 (.Y(n2903), 
	.B1(n8813), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6306));
   INVX1 U4795 (.Y(n8813), 
	.A(\ram[145][1] ));
   OAI22X1 U4796 (.Y(n2902), 
	.B1(n8814), 
	.B0(n8798), 
	.A1(n8797), 
	.A0(n6309));
   INVX1 U4797 (.Y(n8814), 
	.A(\ram[145][0] ));
   NOR2BX1 U4798 (.Y(n8798), 
	.B(n8797), 
	.AN(mem_write_en));
   NAND2X1 U4799 (.Y(n8797), 
	.B(n6495), 
	.A(n8562));
   OAI22X1 U4800 (.Y(n2901), 
	.B1(n8817), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6311));
   INVX1 U4801 (.Y(n8817), 
	.A(\ram[144][15] ));
   OAI22X1 U4802 (.Y(n2900), 
	.B1(n8818), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6314));
   INVX1 U4803 (.Y(n8818), 
	.A(\ram[144][14] ));
   OAI22X1 U4804 (.Y(n2899), 
	.B1(n8819), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6316));
   INVX1 U4805 (.Y(n8819), 
	.A(\ram[144][13] ));
   OAI22X1 U4806 (.Y(n2898), 
	.B1(n8820), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6318));
   INVX1 U4807 (.Y(n8820), 
	.A(\ram[144][12] ));
   OAI22X1 U4808 (.Y(n2897), 
	.B1(n8821), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6320));
   INVX1 U4809 (.Y(n8821), 
	.A(\ram[144][11] ));
   OAI22X1 U4810 (.Y(n2896), 
	.B1(n8822), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6322));
   INVX1 U4811 (.Y(n8822), 
	.A(\ram[144][10] ));
   OAI22X1 U4812 (.Y(n2895), 
	.B1(n8823), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6324));
   INVX1 U4813 (.Y(n8823), 
	.A(\ram[144][9] ));
   OAI22X1 U4814 (.Y(n2894), 
	.B1(n8824), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6326));
   INVX1 U4815 (.Y(n8824), 
	.A(\ram[144][8] ));
   OAI22X1 U4816 (.Y(n2893), 
	.B1(n8825), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6328));
   INVX1 U4817 (.Y(n8825), 
	.A(\ram[144][7] ));
   OAI22X1 U4818 (.Y(n2892), 
	.B1(n8826), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6330));
   INVX1 U4819 (.Y(n8826), 
	.A(\ram[144][6] ));
   OAI22X1 U4820 (.Y(n2891), 
	.B1(n8827), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6332));
   INVX1 U4821 (.Y(n8827), 
	.A(\ram[144][5] ));
   OAI22X1 U4822 (.Y(n2890), 
	.B1(n8828), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6334));
   INVX1 U4823 (.Y(n8828), 
	.A(\ram[144][4] ));
   OAI22X1 U4824 (.Y(n2889), 
	.B1(n8829), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6336));
   INVX1 U4825 (.Y(n8829), 
	.A(\ram[144][3] ));
   OAI22X1 U4826 (.Y(n2888), 
	.B1(n8830), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6338));
   INVX1 U4827 (.Y(n8830), 
	.A(\ram[144][2] ));
   OAI22X1 U4828 (.Y(n2887), 
	.B1(n8831), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6306));
   INVX1 U4829 (.Y(n8831), 
	.A(\ram[144][1] ));
   OAI22X1 U4830 (.Y(n2886), 
	.B1(n8832), 
	.B0(n8816), 
	.A1(n8815), 
	.A0(n6309));
   INVX1 U4831 (.Y(n8832), 
	.A(\ram[144][0] ));
   NOR2BX1 U4832 (.Y(n8816), 
	.B(n8815), 
	.AN(mem_write_en));
   NAND2X1 U4833 (.Y(n8815), 
	.B(n6514), 
	.A(n8562));
   OAI22X1 U4834 (.Y(n2885), 
	.B1(n8835), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6311));
   INVX1 U4835 (.Y(n8835), 
	.A(\ram[143][15] ));
   OAI22X1 U4836 (.Y(n2884), 
	.B1(n8836), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6314));
   INVX1 U4837 (.Y(n8836), 
	.A(\ram[143][14] ));
   OAI22X1 U4838 (.Y(n2883), 
	.B1(n8837), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6316));
   INVX1 U4839 (.Y(n8837), 
	.A(\ram[143][13] ));
   OAI22X1 U4840 (.Y(n2882), 
	.B1(n8838), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6318));
   INVX1 U4841 (.Y(n8838), 
	.A(\ram[143][12] ));
   OAI22X1 U4842 (.Y(n2881), 
	.B1(n8839), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6320));
   INVX1 U4843 (.Y(n8839), 
	.A(\ram[143][11] ));
   OAI22X1 U4844 (.Y(n2880), 
	.B1(n8840), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6322));
   INVX1 U4845 (.Y(n8840), 
	.A(\ram[143][10] ));
   OAI22X1 U4846 (.Y(n2879), 
	.B1(n8841), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6324));
   INVX1 U4847 (.Y(n8841), 
	.A(\ram[143][9] ));
   OAI22X1 U4848 (.Y(n2878), 
	.B1(n8842), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6326));
   INVX1 U4849 (.Y(n8842), 
	.A(\ram[143][8] ));
   OAI22X1 U4850 (.Y(n2877), 
	.B1(n8843), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6328));
   INVX1 U4851 (.Y(n8843), 
	.A(\ram[143][7] ));
   OAI22X1 U4852 (.Y(n2876), 
	.B1(n8844), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6330));
   INVX1 U4853 (.Y(n8844), 
	.A(\ram[143][6] ));
   OAI22X1 U4854 (.Y(n2875), 
	.B1(n8845), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6332));
   INVX1 U4855 (.Y(n8845), 
	.A(\ram[143][5] ));
   OAI22X1 U4856 (.Y(n2874), 
	.B1(n8846), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6334));
   INVX1 U4857 (.Y(n8846), 
	.A(\ram[143][4] ));
   OAI22X1 U4858 (.Y(n2873), 
	.B1(n8847), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6336));
   INVX1 U4859 (.Y(n8847), 
	.A(\ram[143][3] ));
   OAI22X1 U4860 (.Y(n2872), 
	.B1(n8848), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6338));
   INVX1 U4861 (.Y(n8848), 
	.A(\ram[143][2] ));
   OAI22X1 U4862 (.Y(n2871), 
	.B1(n8849), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6306));
   INVX1 U4863 (.Y(n8849), 
	.A(\ram[143][1] ));
   OAI22X1 U4864 (.Y(n2870), 
	.B1(n8850), 
	.B0(n8834), 
	.A1(n8833), 
	.A0(n6309));
   INVX1 U4865 (.Y(n8850), 
	.A(\ram[143][0] ));
   NOR2BX1 U4866 (.Y(n8834), 
	.B(n8833), 
	.AN(mem_write_en));
   NAND2X1 U4867 (.Y(n8833), 
	.B(n6533), 
	.A(n8851));
   OAI22X1 U4868 (.Y(n2869), 
	.B1(n8854), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6311));
   INVX1 U4869 (.Y(n8854), 
	.A(\ram[142][15] ));
   OAI22X1 U4870 (.Y(n2868), 
	.B1(n8855), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6314));
   INVX1 U4871 (.Y(n8855), 
	.A(\ram[142][14] ));
   OAI22X1 U4872 (.Y(n2867), 
	.B1(n8856), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6316));
   INVX1 U4873 (.Y(n8856), 
	.A(\ram[142][13] ));
   OAI22X1 U4874 (.Y(n2866), 
	.B1(n8857), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6318));
   INVX1 U4875 (.Y(n8857), 
	.A(\ram[142][12] ));
   OAI22X1 U4876 (.Y(n2865), 
	.B1(n8858), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6320));
   INVX1 U4877 (.Y(n8858), 
	.A(\ram[142][11] ));
   OAI22X1 U4878 (.Y(n2864), 
	.B1(n8859), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6322));
   INVX1 U4879 (.Y(n8859), 
	.A(\ram[142][10] ));
   OAI22X1 U4880 (.Y(n2863), 
	.B1(n8860), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6324));
   INVX1 U4881 (.Y(n8860), 
	.A(\ram[142][9] ));
   OAI22X1 U4882 (.Y(n2862), 
	.B1(n8861), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6326));
   INVX1 U4883 (.Y(n8861), 
	.A(\ram[142][8] ));
   OAI22X1 U4884 (.Y(n2861), 
	.B1(n8862), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6328));
   INVX1 U4885 (.Y(n8862), 
	.A(\ram[142][7] ));
   OAI22X1 U4886 (.Y(n2860), 
	.B1(n8863), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6330));
   INVX1 U4887 (.Y(n8863), 
	.A(\ram[142][6] ));
   OAI22X1 U4888 (.Y(n2859), 
	.B1(n8864), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6332));
   INVX1 U4889 (.Y(n8864), 
	.A(\ram[142][5] ));
   OAI22X1 U4890 (.Y(n2858), 
	.B1(n8865), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6334));
   INVX1 U4891 (.Y(n8865), 
	.A(\ram[142][4] ));
   OAI22X1 U4892 (.Y(n2857), 
	.B1(n8866), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6336));
   INVX1 U4893 (.Y(n8866), 
	.A(\ram[142][3] ));
   OAI22X1 U4894 (.Y(n2856), 
	.B1(n8867), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6338));
   INVX1 U4895 (.Y(n8867), 
	.A(\ram[142][2] ));
   OAI22X1 U4896 (.Y(n2855), 
	.B1(n8868), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6306));
   INVX1 U4897 (.Y(n8868), 
	.A(\ram[142][1] ));
   OAI22X1 U4898 (.Y(n2854), 
	.B1(n8869), 
	.B0(n8853), 
	.A1(n8852), 
	.A0(n6309));
   INVX1 U4899 (.Y(n8869), 
	.A(\ram[142][0] ));
   NOR2BX1 U4900 (.Y(n8853), 
	.B(n8852), 
	.AN(mem_write_en));
   NAND2X1 U4901 (.Y(n8852), 
	.B(n6553), 
	.A(n8851));
   OAI22X1 U4902 (.Y(n2853), 
	.B1(n8872), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6311));
   INVX1 U4903 (.Y(n8872), 
	.A(\ram[141][15] ));
   OAI22X1 U4904 (.Y(n2852), 
	.B1(n8873), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6314));
   INVX1 U4905 (.Y(n8873), 
	.A(\ram[141][14] ));
   OAI22X1 U4906 (.Y(n2851), 
	.B1(n8874), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6316));
   INVX1 U4907 (.Y(n8874), 
	.A(\ram[141][13] ));
   OAI22X1 U4908 (.Y(n2850), 
	.B1(n8875), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6318));
   INVX1 U4909 (.Y(n8875), 
	.A(\ram[141][12] ));
   OAI22X1 U4910 (.Y(n2849), 
	.B1(n8876), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6320));
   INVX1 U4911 (.Y(n8876), 
	.A(\ram[141][11] ));
   OAI22X1 U4912 (.Y(n2848), 
	.B1(n8877), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6322));
   INVX1 U4913 (.Y(n8877), 
	.A(\ram[141][10] ));
   OAI22X1 U4914 (.Y(n2847), 
	.B1(n8878), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6324));
   INVX1 U4915 (.Y(n8878), 
	.A(\ram[141][9] ));
   OAI22X1 U4916 (.Y(n2846), 
	.B1(n8879), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6326));
   INVX1 U4917 (.Y(n8879), 
	.A(\ram[141][8] ));
   OAI22X1 U4918 (.Y(n2845), 
	.B1(n8880), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6328));
   INVX1 U4919 (.Y(n8880), 
	.A(\ram[141][7] ));
   OAI22X1 U4920 (.Y(n2844), 
	.B1(n8881), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6330));
   INVX1 U4921 (.Y(n8881), 
	.A(\ram[141][6] ));
   OAI22X1 U4922 (.Y(n2843), 
	.B1(n8882), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6332));
   INVX1 U4923 (.Y(n8882), 
	.A(\ram[141][5] ));
   OAI22X1 U4924 (.Y(n2842), 
	.B1(n8883), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6334));
   INVX1 U4925 (.Y(n8883), 
	.A(\ram[141][4] ));
   OAI22X1 U4926 (.Y(n2841), 
	.B1(n8884), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6336));
   INVX1 U4927 (.Y(n8884), 
	.A(\ram[141][3] ));
   OAI22X1 U4928 (.Y(n2840), 
	.B1(n8885), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6338));
   INVX1 U4929 (.Y(n8885), 
	.A(\ram[141][2] ));
   OAI22X1 U4930 (.Y(n2839), 
	.B1(n8886), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6306));
   INVX1 U4931 (.Y(n8886), 
	.A(\ram[141][1] ));
   OAI22X1 U4932 (.Y(n2838), 
	.B1(n8887), 
	.B0(n8871), 
	.A1(n8870), 
	.A0(n6309));
   INVX1 U4933 (.Y(n8887), 
	.A(\ram[141][0] ));
   NOR2BX1 U4934 (.Y(n8871), 
	.B(n8870), 
	.AN(mem_write_en));
   NAND2X1 U4935 (.Y(n8870), 
	.B(n6572), 
	.A(n8851));
   OAI22X1 U4936 (.Y(n2837), 
	.B1(n8890), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6311));
   INVX1 U4937 (.Y(n8890), 
	.A(\ram[140][15] ));
   OAI22X1 U4938 (.Y(n2836), 
	.B1(n8891), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6314));
   INVX1 U4939 (.Y(n8891), 
	.A(\ram[140][14] ));
   OAI22X1 U4940 (.Y(n2835), 
	.B1(n8892), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6316));
   INVX1 U4941 (.Y(n8892), 
	.A(\ram[140][13] ));
   OAI22X1 U4942 (.Y(n2834), 
	.B1(n8893), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6318));
   INVX1 U4943 (.Y(n8893), 
	.A(\ram[140][12] ));
   OAI22X1 U4944 (.Y(n2833), 
	.B1(n8894), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6320));
   INVX1 U4945 (.Y(n8894), 
	.A(\ram[140][11] ));
   OAI22X1 U4946 (.Y(n2832), 
	.B1(n8895), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6322));
   INVX1 U4947 (.Y(n8895), 
	.A(\ram[140][10] ));
   OAI22X1 U4948 (.Y(n2831), 
	.B1(n8896), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6324));
   INVX1 U4949 (.Y(n8896), 
	.A(\ram[140][9] ));
   OAI22X1 U4950 (.Y(n2830), 
	.B1(n8897), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6326));
   INVX1 U4951 (.Y(n8897), 
	.A(\ram[140][8] ));
   OAI22X1 U4952 (.Y(n2829), 
	.B1(n8898), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6328));
   INVX1 U4953 (.Y(n8898), 
	.A(\ram[140][7] ));
   OAI22X1 U4954 (.Y(n2828), 
	.B1(n8899), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6330));
   INVX1 U4955 (.Y(n8899), 
	.A(\ram[140][6] ));
   OAI22X1 U4956 (.Y(n2827), 
	.B1(n8900), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6332));
   INVX1 U4957 (.Y(n8900), 
	.A(\ram[140][5] ));
   OAI22X1 U4958 (.Y(n2826), 
	.B1(n8901), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6334));
   INVX1 U4959 (.Y(n8901), 
	.A(\ram[140][4] ));
   OAI22X1 U4960 (.Y(n2825), 
	.B1(n8902), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6336));
   INVX1 U4961 (.Y(n8902), 
	.A(\ram[140][3] ));
   OAI22X1 U4962 (.Y(n2824), 
	.B1(n8903), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6338));
   INVX1 U4963 (.Y(n8903), 
	.A(\ram[140][2] ));
   OAI22X1 U4964 (.Y(n2823), 
	.B1(n8904), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6306));
   INVX1 U4965 (.Y(n8904), 
	.A(\ram[140][1] ));
   OAI22X1 U4966 (.Y(n2822), 
	.B1(n8905), 
	.B0(n8889), 
	.A1(n8888), 
	.A0(n6309));
   INVX1 U4967 (.Y(n8905), 
	.A(\ram[140][0] ));
   NOR2BX1 U4968 (.Y(n8889), 
	.B(n8888), 
	.AN(mem_write_en));
   NAND2X1 U4969 (.Y(n8888), 
	.B(n6591), 
	.A(n8851));
   OAI22X1 U4970 (.Y(n2821), 
	.B1(n8908), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6311));
   INVX1 U4971 (.Y(n8908), 
	.A(\ram[139][15] ));
   OAI22X1 U4972 (.Y(n2820), 
	.B1(n8909), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6314));
   INVX1 U4973 (.Y(n8909), 
	.A(\ram[139][14] ));
   OAI22X1 U4974 (.Y(n2819), 
	.B1(n8910), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6316));
   INVX1 U4975 (.Y(n8910), 
	.A(\ram[139][13] ));
   OAI22X1 U4976 (.Y(n2818), 
	.B1(n8911), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6318));
   INVX1 U4977 (.Y(n8911), 
	.A(\ram[139][12] ));
   OAI22X1 U4978 (.Y(n2817), 
	.B1(n8912), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6320));
   INVX1 U4979 (.Y(n8912), 
	.A(\ram[139][11] ));
   OAI22X1 U4980 (.Y(n2816), 
	.B1(n8913), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6322));
   INVX1 U4981 (.Y(n8913), 
	.A(\ram[139][10] ));
   OAI22X1 U4982 (.Y(n2815), 
	.B1(n8914), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6324));
   INVX1 U4983 (.Y(n8914), 
	.A(\ram[139][9] ));
   OAI22X1 U4984 (.Y(n2814), 
	.B1(n8915), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6326));
   INVX1 U4985 (.Y(n8915), 
	.A(\ram[139][8] ));
   OAI22X1 U4986 (.Y(n2813), 
	.B1(n8916), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6328));
   INVX1 U4987 (.Y(n8916), 
	.A(\ram[139][7] ));
   OAI22X1 U4988 (.Y(n2812), 
	.B1(n8917), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6330));
   INVX1 U4989 (.Y(n8917), 
	.A(\ram[139][6] ));
   OAI22X1 U4990 (.Y(n2811), 
	.B1(n8918), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6332));
   INVX1 U4991 (.Y(n8918), 
	.A(\ram[139][5] ));
   OAI22X1 U4992 (.Y(n2810), 
	.B1(n8919), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6334));
   INVX1 U4993 (.Y(n8919), 
	.A(\ram[139][4] ));
   OAI22X1 U4994 (.Y(n2809), 
	.B1(n8920), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6336));
   INVX1 U4995 (.Y(n8920), 
	.A(\ram[139][3] ));
   OAI22X1 U4996 (.Y(n2808), 
	.B1(n8921), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6338));
   INVX1 U4997 (.Y(n8921), 
	.A(\ram[139][2] ));
   OAI22X1 U4998 (.Y(n2807), 
	.B1(n8922), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6306));
   INVX1 U4999 (.Y(n8922), 
	.A(\ram[139][1] ));
   OAI22X1 U5000 (.Y(n2806), 
	.B1(n8923), 
	.B0(n8907), 
	.A1(n8906), 
	.A0(n6309));
   INVX1 U5001 (.Y(n8923), 
	.A(\ram[139][0] ));
   NOR2BX1 U5002 (.Y(n8907), 
	.B(n8906), 
	.AN(mem_write_en));
   NAND2X1 U5003 (.Y(n8906), 
	.B(n6610), 
	.A(n8851));
   OAI22X1 U5004 (.Y(n2805), 
	.B1(n8926), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6311));
   INVX1 U5005 (.Y(n8926), 
	.A(\ram[138][15] ));
   OAI22X1 U5006 (.Y(n2804), 
	.B1(n8927), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6314));
   INVX1 U5007 (.Y(n8927), 
	.A(\ram[138][14] ));
   OAI22X1 U5008 (.Y(n2803), 
	.B1(n8928), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6316));
   INVX1 U5009 (.Y(n8928), 
	.A(\ram[138][13] ));
   OAI22X1 U5010 (.Y(n2802), 
	.B1(n8929), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6318));
   INVX1 U5011 (.Y(n8929), 
	.A(\ram[138][12] ));
   OAI22X1 U5012 (.Y(n2801), 
	.B1(n8930), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6320));
   INVX1 U5013 (.Y(n8930), 
	.A(\ram[138][11] ));
   OAI22X1 U5014 (.Y(n2800), 
	.B1(n8931), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6322));
   INVX1 U5015 (.Y(n8931), 
	.A(\ram[138][10] ));
   OAI22X1 U5016 (.Y(n2799), 
	.B1(n8932), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6324));
   INVX1 U5017 (.Y(n8932), 
	.A(\ram[138][9] ));
   OAI22X1 U5018 (.Y(n2798), 
	.B1(n8933), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6326));
   INVX1 U5019 (.Y(n8933), 
	.A(\ram[138][8] ));
   OAI22X1 U5020 (.Y(n2797), 
	.B1(n8934), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6328));
   INVX1 U5021 (.Y(n8934), 
	.A(\ram[138][7] ));
   OAI22X1 U5022 (.Y(n2796), 
	.B1(n8935), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6330));
   INVX1 U5023 (.Y(n8935), 
	.A(\ram[138][6] ));
   OAI22X1 U5024 (.Y(n2795), 
	.B1(n8936), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6332));
   INVX1 U5025 (.Y(n8936), 
	.A(\ram[138][5] ));
   OAI22X1 U5026 (.Y(n2794), 
	.B1(n8937), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6334));
   INVX1 U5027 (.Y(n8937), 
	.A(\ram[138][4] ));
   OAI22X1 U5028 (.Y(n2793), 
	.B1(n8938), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6336));
   INVX1 U5029 (.Y(n8938), 
	.A(\ram[138][3] ));
   OAI22X1 U5030 (.Y(n2792), 
	.B1(n8939), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6338));
   INVX1 U5031 (.Y(n8939), 
	.A(\ram[138][2] ));
   OAI22X1 U5032 (.Y(n2791), 
	.B1(n8940), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6306));
   INVX1 U5033 (.Y(n8940), 
	.A(\ram[138][1] ));
   OAI22X1 U5034 (.Y(n2790), 
	.B1(n8941), 
	.B0(n8925), 
	.A1(n8924), 
	.A0(n6309));
   INVX1 U5035 (.Y(n8941), 
	.A(\ram[138][0] ));
   NOR2BX1 U5036 (.Y(n8925), 
	.B(n8924), 
	.AN(mem_write_en));
   NAND2X1 U5037 (.Y(n8924), 
	.B(n6629), 
	.A(n8851));
   OAI22X1 U5038 (.Y(n2789), 
	.B1(n8944), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6311));
   INVX1 U5039 (.Y(n8944), 
	.A(\ram[137][15] ));
   OAI22X1 U5040 (.Y(n2788), 
	.B1(n8945), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6314));
   INVX1 U5041 (.Y(n8945), 
	.A(\ram[137][14] ));
   OAI22X1 U5042 (.Y(n2787), 
	.B1(n8946), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6316));
   INVX1 U5043 (.Y(n8946), 
	.A(\ram[137][13] ));
   OAI22X1 U5044 (.Y(n2786), 
	.B1(n8947), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6318));
   INVX1 U5045 (.Y(n8947), 
	.A(\ram[137][12] ));
   OAI22X1 U5046 (.Y(n2785), 
	.B1(n8948), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6320));
   INVX1 U5047 (.Y(n8948), 
	.A(\ram[137][11] ));
   OAI22X1 U5048 (.Y(n2784), 
	.B1(n8949), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6322));
   INVX1 U5049 (.Y(n8949), 
	.A(\ram[137][10] ));
   OAI22X1 U5050 (.Y(n2783), 
	.B1(n8950), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6324));
   INVX1 U5051 (.Y(n8950), 
	.A(\ram[137][9] ));
   OAI22X1 U5052 (.Y(n2782), 
	.B1(n8951), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6326));
   INVX1 U5053 (.Y(n8951), 
	.A(\ram[137][8] ));
   OAI22X1 U5054 (.Y(n2781), 
	.B1(n8952), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6328));
   INVX1 U5055 (.Y(n8952), 
	.A(\ram[137][7] ));
   OAI22X1 U5056 (.Y(n2780), 
	.B1(n8953), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6330));
   INVX1 U5057 (.Y(n8953), 
	.A(\ram[137][6] ));
   OAI22X1 U5058 (.Y(n2779), 
	.B1(n8954), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6332));
   INVX1 U5059 (.Y(n8954), 
	.A(\ram[137][5] ));
   OAI22X1 U5060 (.Y(n2778), 
	.B1(n8955), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6334));
   INVX1 U5061 (.Y(n8955), 
	.A(\ram[137][4] ));
   OAI22X1 U5062 (.Y(n2777), 
	.B1(n8956), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6336));
   INVX1 U5063 (.Y(n8956), 
	.A(\ram[137][3] ));
   OAI22X1 U5064 (.Y(n2776), 
	.B1(n8957), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6338));
   INVX1 U5065 (.Y(n8957), 
	.A(\ram[137][2] ));
   OAI22X1 U5066 (.Y(n2775), 
	.B1(n8958), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6306));
   INVX1 U5067 (.Y(n8958), 
	.A(\ram[137][1] ));
   OAI22X1 U5068 (.Y(n2774), 
	.B1(n8959), 
	.B0(n8943), 
	.A1(n8942), 
	.A0(n6309));
   INVX1 U5069 (.Y(n8959), 
	.A(\ram[137][0] ));
   NOR2BX1 U5070 (.Y(n8943), 
	.B(n8942), 
	.AN(mem_write_en));
   NAND2X1 U5071 (.Y(n8942), 
	.B(n6342), 
	.A(n8851));
   OAI22X1 U5072 (.Y(n2773), 
	.B1(n8962), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6311));
   INVX1 U5073 (.Y(n8962), 
	.A(\ram[136][15] ));
   OAI22X1 U5074 (.Y(n2772), 
	.B1(n8963), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6314));
   INVX1 U5075 (.Y(n8963), 
	.A(\ram[136][14] ));
   OAI22X1 U5076 (.Y(n2771), 
	.B1(n8964), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6316));
   INVX1 U5077 (.Y(n8964), 
	.A(\ram[136][13] ));
   OAI22X1 U5078 (.Y(n2770), 
	.B1(n8965), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6318));
   INVX1 U5079 (.Y(n8965), 
	.A(\ram[136][12] ));
   OAI22X1 U5080 (.Y(n2769), 
	.B1(n8966), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6320));
   INVX1 U5081 (.Y(n8966), 
	.A(\ram[136][11] ));
   OAI22X1 U5082 (.Y(n2768), 
	.B1(n8967), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6322));
   INVX1 U5083 (.Y(n8967), 
	.A(\ram[136][10] ));
   OAI22X1 U5084 (.Y(n2767), 
	.B1(n8968), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6324));
   INVX1 U5085 (.Y(n8968), 
	.A(\ram[136][9] ));
   OAI22X1 U5086 (.Y(n2766), 
	.B1(n8969), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6326));
   INVX1 U5087 (.Y(n8969), 
	.A(\ram[136][8] ));
   OAI22X1 U5088 (.Y(n2765), 
	.B1(n8970), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6328));
   INVX1 U5089 (.Y(n8970), 
	.A(\ram[136][7] ));
   OAI22X1 U5090 (.Y(n2764), 
	.B1(n8971), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6330));
   INVX1 U5091 (.Y(n8971), 
	.A(\ram[136][6] ));
   OAI22X1 U5092 (.Y(n2763), 
	.B1(n8972), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6332));
   INVX1 U5093 (.Y(n8972), 
	.A(\ram[136][5] ));
   OAI22X1 U5094 (.Y(n2762), 
	.B1(n8973), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6334));
   INVX1 U5095 (.Y(n8973), 
	.A(\ram[136][4] ));
   OAI22X1 U5096 (.Y(n2761), 
	.B1(n8974), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6336));
   INVX1 U5097 (.Y(n8974), 
	.A(\ram[136][3] ));
   OAI22X1 U5098 (.Y(n2760), 
	.B1(n8975), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6338));
   INVX1 U5099 (.Y(n8975), 
	.A(\ram[136][2] ));
   OAI22X1 U5100 (.Y(n2759), 
	.B1(n8976), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6306));
   INVX1 U5101 (.Y(n8976), 
	.A(\ram[136][1] ));
   OAI22X1 U5102 (.Y(n2758), 
	.B1(n8977), 
	.B0(n8961), 
	.A1(n8960), 
	.A0(n6309));
   INVX1 U5103 (.Y(n8977), 
	.A(\ram[136][0] ));
   NOR2BX1 U5104 (.Y(n8961), 
	.B(n8960), 
	.AN(mem_write_en));
   NAND2X1 U5105 (.Y(n8960), 
	.B(n6362), 
	.A(n8851));
   OAI22X1 U5106 (.Y(n2757), 
	.B1(n8980), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6311));
   INVX1 U5107 (.Y(n8980), 
	.A(\ram[135][15] ));
   OAI22X1 U5108 (.Y(n2756), 
	.B1(n8981), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6314));
   INVX1 U5109 (.Y(n8981), 
	.A(\ram[135][14] ));
   OAI22X1 U5110 (.Y(n2755), 
	.B1(n8982), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6316));
   INVX1 U5111 (.Y(n8982), 
	.A(\ram[135][13] ));
   OAI22X1 U5112 (.Y(n2754), 
	.B1(n8983), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6318));
   INVX1 U5113 (.Y(n8983), 
	.A(\ram[135][12] ));
   OAI22X1 U5114 (.Y(n2753), 
	.B1(n8984), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6320));
   INVX1 U5115 (.Y(n8984), 
	.A(\ram[135][11] ));
   OAI22X1 U5116 (.Y(n2752), 
	.B1(n8985), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6322));
   INVX1 U5117 (.Y(n8985), 
	.A(\ram[135][10] ));
   OAI22X1 U5118 (.Y(n2751), 
	.B1(n8986), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6324));
   INVX1 U5119 (.Y(n8986), 
	.A(\ram[135][9] ));
   OAI22X1 U5120 (.Y(n2750), 
	.B1(n8987), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6326));
   INVX1 U5121 (.Y(n8987), 
	.A(\ram[135][8] ));
   OAI22X1 U5122 (.Y(n2749), 
	.B1(n8988), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6328));
   INVX1 U5123 (.Y(n8988), 
	.A(\ram[135][7] ));
   OAI22X1 U5124 (.Y(n2748), 
	.B1(n8989), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6330));
   INVX1 U5125 (.Y(n8989), 
	.A(\ram[135][6] ));
   OAI22X1 U5126 (.Y(n2747), 
	.B1(n8990), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6332));
   INVX1 U5127 (.Y(n8990), 
	.A(\ram[135][5] ));
   OAI22X1 U5128 (.Y(n2746), 
	.B1(n8991), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6334));
   INVX1 U5129 (.Y(n8991), 
	.A(\ram[135][4] ));
   OAI22X1 U5130 (.Y(n2745), 
	.B1(n8992), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6336));
   INVX1 U5131 (.Y(n8992), 
	.A(\ram[135][3] ));
   OAI22X1 U5132 (.Y(n2744), 
	.B1(n8993), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6338));
   INVX1 U5133 (.Y(n8993), 
	.A(\ram[135][2] ));
   OAI22X1 U5134 (.Y(n2743), 
	.B1(n8994), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6306));
   INVX1 U5135 (.Y(n8994), 
	.A(\ram[135][1] ));
   OAI22X1 U5136 (.Y(n2742), 
	.B1(n8995), 
	.B0(n8979), 
	.A1(n8978), 
	.A0(n6309));
   INVX1 U5137 (.Y(n8995), 
	.A(\ram[135][0] ));
   NOR2BX1 U5138 (.Y(n8979), 
	.B(n8978), 
	.AN(mem_write_en));
   NAND2X1 U5139 (.Y(n8978), 
	.B(n6381), 
	.A(n8851));
   OAI22X1 U5140 (.Y(n2741), 
	.B1(n8998), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6311));
   INVX1 U5141 (.Y(n8998), 
	.A(\ram[134][15] ));
   OAI22X1 U5142 (.Y(n2740), 
	.B1(n8999), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6314));
   INVX1 U5143 (.Y(n8999), 
	.A(\ram[134][14] ));
   OAI22X1 U5144 (.Y(n2739), 
	.B1(n9000), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6316));
   INVX1 U5145 (.Y(n9000), 
	.A(\ram[134][13] ));
   OAI22X1 U5146 (.Y(n2738), 
	.B1(n9001), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6318));
   INVX1 U5147 (.Y(n9001), 
	.A(\ram[134][12] ));
   OAI22X1 U5148 (.Y(n2737), 
	.B1(n9002), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6320));
   INVX1 U5149 (.Y(n9002), 
	.A(\ram[134][11] ));
   OAI22X1 U5150 (.Y(n2736), 
	.B1(n9003), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6322));
   INVX1 U5151 (.Y(n9003), 
	.A(\ram[134][10] ));
   OAI22X1 U5152 (.Y(n2735), 
	.B1(n9004), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6324));
   INVX1 U5153 (.Y(n9004), 
	.A(\ram[134][9] ));
   OAI22X1 U5154 (.Y(n2734), 
	.B1(n9005), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6326));
   INVX1 U5155 (.Y(n9005), 
	.A(\ram[134][8] ));
   OAI22X1 U5156 (.Y(n2733), 
	.B1(n9006), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6328));
   INVX1 U5157 (.Y(n9006), 
	.A(\ram[134][7] ));
   OAI22X1 U5158 (.Y(n2732), 
	.B1(n9007), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6330));
   INVX1 U5159 (.Y(n9007), 
	.A(\ram[134][6] ));
   OAI22X1 U5160 (.Y(n2731), 
	.B1(n9008), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6332));
   INVX1 U5161 (.Y(n9008), 
	.A(\ram[134][5] ));
   OAI22X1 U5162 (.Y(n2730), 
	.B1(n9009), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6334));
   INVX1 U5163 (.Y(n9009), 
	.A(\ram[134][4] ));
   OAI22X1 U5164 (.Y(n2729), 
	.B1(n9010), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6336));
   INVX1 U5165 (.Y(n9010), 
	.A(\ram[134][3] ));
   OAI22X1 U5166 (.Y(n2728), 
	.B1(n9011), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6338));
   INVX1 U5167 (.Y(n9011), 
	.A(\ram[134][2] ));
   OAI22X1 U5168 (.Y(n2727), 
	.B1(n9012), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6306));
   INVX1 U5169 (.Y(n9012), 
	.A(\ram[134][1] ));
   OAI22X1 U5170 (.Y(n2726), 
	.B1(n9013), 
	.B0(n8997), 
	.A1(n8996), 
	.A0(n6309));
   INVX1 U5171 (.Y(n9013), 
	.A(\ram[134][0] ));
   NOR2BX1 U5172 (.Y(n8997), 
	.B(n8996), 
	.AN(mem_write_en));
   NAND2X1 U5173 (.Y(n8996), 
	.B(n6400), 
	.A(n8851));
   OAI22X1 U5174 (.Y(n2725), 
	.B1(n9016), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6311));
   INVX1 U5175 (.Y(n9016), 
	.A(\ram[133][15] ));
   OAI22X1 U5176 (.Y(n2724), 
	.B1(n9017), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6314));
   INVX1 U5177 (.Y(n9017), 
	.A(\ram[133][14] ));
   OAI22X1 U5178 (.Y(n2723), 
	.B1(n9018), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6316));
   INVX1 U5179 (.Y(n9018), 
	.A(\ram[133][13] ));
   OAI22X1 U5180 (.Y(n2722), 
	.B1(n9019), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6318));
   INVX1 U5181 (.Y(n9019), 
	.A(\ram[133][12] ));
   OAI22X1 U5182 (.Y(n2721), 
	.B1(n9020), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6320));
   INVX1 U5183 (.Y(n9020), 
	.A(\ram[133][11] ));
   OAI22X1 U5184 (.Y(n2720), 
	.B1(n9021), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6322));
   INVX1 U5185 (.Y(n9021), 
	.A(\ram[133][10] ));
   OAI22X1 U5186 (.Y(n2719), 
	.B1(n9022), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6324));
   INVX1 U5187 (.Y(n9022), 
	.A(\ram[133][9] ));
   OAI22X1 U5188 (.Y(n2718), 
	.B1(n9023), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6326));
   INVX1 U5189 (.Y(n9023), 
	.A(\ram[133][8] ));
   OAI22X1 U5190 (.Y(n2717), 
	.B1(n9024), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6328));
   INVX1 U5191 (.Y(n9024), 
	.A(\ram[133][7] ));
   OAI22X1 U5192 (.Y(n2716), 
	.B1(n9025), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6330));
   INVX1 U5193 (.Y(n9025), 
	.A(\ram[133][6] ));
   OAI22X1 U5194 (.Y(n2715), 
	.B1(n9026), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6332));
   INVX1 U5195 (.Y(n9026), 
	.A(\ram[133][5] ));
   OAI22X1 U5196 (.Y(n2714), 
	.B1(n9027), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6334));
   INVX1 U5197 (.Y(n9027), 
	.A(\ram[133][4] ));
   OAI22X1 U5198 (.Y(n2713), 
	.B1(n9028), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6336));
   INVX1 U5199 (.Y(n9028), 
	.A(\ram[133][3] ));
   OAI22X1 U5200 (.Y(n2712), 
	.B1(n9029), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6338));
   INVX1 U5201 (.Y(n9029), 
	.A(\ram[133][2] ));
   OAI22X1 U5202 (.Y(n2711), 
	.B1(n9030), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6306));
   INVX1 U5203 (.Y(n9030), 
	.A(\ram[133][1] ));
   OAI22X1 U5204 (.Y(n2710), 
	.B1(n9031), 
	.B0(n9015), 
	.A1(n9014), 
	.A0(n6309));
   INVX1 U5205 (.Y(n9031), 
	.A(\ram[133][0] ));
   NOR2BX1 U5206 (.Y(n9015), 
	.B(n9014), 
	.AN(mem_write_en));
   NAND2X1 U5207 (.Y(n9014), 
	.B(n6419), 
	.A(n8851));
   OAI22X1 U5208 (.Y(n2709), 
	.B1(n9034), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6311));
   INVX1 U5209 (.Y(n9034), 
	.A(\ram[132][15] ));
   OAI22X1 U5210 (.Y(n2708), 
	.B1(n9035), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6314));
   INVX1 U5211 (.Y(n9035), 
	.A(\ram[132][14] ));
   OAI22X1 U5212 (.Y(n2707), 
	.B1(n9036), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6316));
   INVX1 U5213 (.Y(n9036), 
	.A(\ram[132][13] ));
   OAI22X1 U5214 (.Y(n2706), 
	.B1(n9037), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6318));
   INVX1 U5215 (.Y(n9037), 
	.A(\ram[132][12] ));
   OAI22X1 U5216 (.Y(n2705), 
	.B1(n9038), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6320));
   INVX1 U5217 (.Y(n9038), 
	.A(\ram[132][11] ));
   OAI22X1 U5218 (.Y(n2704), 
	.B1(n9039), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6322));
   INVX1 U5219 (.Y(n9039), 
	.A(\ram[132][10] ));
   OAI22X1 U5220 (.Y(n2703), 
	.B1(n9040), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6324));
   INVX1 U5221 (.Y(n9040), 
	.A(\ram[132][9] ));
   OAI22X1 U5222 (.Y(n2702), 
	.B1(n9041), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6326));
   INVX1 U5223 (.Y(n9041), 
	.A(\ram[132][8] ));
   OAI22X1 U5224 (.Y(n2701), 
	.B1(n9042), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6328));
   INVX1 U5225 (.Y(n9042), 
	.A(\ram[132][7] ));
   OAI22X1 U5226 (.Y(n2700), 
	.B1(n9043), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6330));
   INVX1 U5227 (.Y(n9043), 
	.A(\ram[132][6] ));
   OAI22X1 U5228 (.Y(n2699), 
	.B1(n9044), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6332));
   INVX1 U5229 (.Y(n9044), 
	.A(\ram[132][5] ));
   OAI22X1 U5230 (.Y(n2698), 
	.B1(n9045), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6334));
   INVX1 U5231 (.Y(n9045), 
	.A(\ram[132][4] ));
   OAI22X1 U5232 (.Y(n2697), 
	.B1(n9046), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6336));
   INVX1 U5233 (.Y(n9046), 
	.A(\ram[132][3] ));
   OAI22X1 U5234 (.Y(n2696), 
	.B1(n9047), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6338));
   INVX1 U5235 (.Y(n9047), 
	.A(\ram[132][2] ));
   OAI22X1 U5236 (.Y(n2695), 
	.B1(n9048), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6306));
   INVX1 U5237 (.Y(n9048), 
	.A(\ram[132][1] ));
   OAI22X1 U5238 (.Y(n2694), 
	.B1(n9049), 
	.B0(n9033), 
	.A1(n9032), 
	.A0(n6309));
   INVX1 U5239 (.Y(n9049), 
	.A(\ram[132][0] ));
   NOR2BX1 U5240 (.Y(n9033), 
	.B(n9032), 
	.AN(mem_write_en));
   NAND2X1 U5241 (.Y(n9032), 
	.B(n6438), 
	.A(n8851));
   OAI22X1 U5242 (.Y(n2693), 
	.B1(n9052), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6311));
   INVX1 U5243 (.Y(n9052), 
	.A(\ram[131][15] ));
   OAI22X1 U5244 (.Y(n2692), 
	.B1(n9053), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6314));
   INVX1 U5245 (.Y(n9053), 
	.A(\ram[131][14] ));
   OAI22X1 U5246 (.Y(n2691), 
	.B1(n9054), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6316));
   INVX1 U5247 (.Y(n9054), 
	.A(\ram[131][13] ));
   OAI22X1 U5248 (.Y(n2690), 
	.B1(n9055), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6318));
   INVX1 U5249 (.Y(n9055), 
	.A(\ram[131][12] ));
   OAI22X1 U5250 (.Y(n2689), 
	.B1(n9056), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6320));
   INVX1 U5251 (.Y(n9056), 
	.A(\ram[131][11] ));
   OAI22X1 U5252 (.Y(n2688), 
	.B1(n9057), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6322));
   INVX1 U5253 (.Y(n9057), 
	.A(\ram[131][10] ));
   OAI22X1 U5254 (.Y(n2687), 
	.B1(n9058), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6324));
   INVX1 U5255 (.Y(n9058), 
	.A(\ram[131][9] ));
   OAI22X1 U5256 (.Y(n2686), 
	.B1(n9059), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6326));
   INVX1 U5257 (.Y(n9059), 
	.A(\ram[131][8] ));
   OAI22X1 U5258 (.Y(n2685), 
	.B1(n9060), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6328));
   INVX1 U5259 (.Y(n9060), 
	.A(\ram[131][7] ));
   OAI22X1 U5260 (.Y(n2684), 
	.B1(n9061), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6330));
   INVX1 U5261 (.Y(n9061), 
	.A(\ram[131][6] ));
   OAI22X1 U5262 (.Y(n2683), 
	.B1(n9062), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6332));
   INVX1 U5263 (.Y(n9062), 
	.A(\ram[131][5] ));
   OAI22X1 U5264 (.Y(n2682), 
	.B1(n9063), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6334));
   INVX1 U5265 (.Y(n9063), 
	.A(\ram[131][4] ));
   OAI22X1 U5266 (.Y(n2681), 
	.B1(n9064), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6336));
   INVX1 U5267 (.Y(n9064), 
	.A(\ram[131][3] ));
   OAI22X1 U5268 (.Y(n2680), 
	.B1(n9065), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6338));
   INVX1 U5269 (.Y(n9065), 
	.A(\ram[131][2] ));
   OAI22X1 U5270 (.Y(n2679), 
	.B1(n9066), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6306));
   INVX1 U5271 (.Y(n9066), 
	.A(\ram[131][1] ));
   OAI22X1 U5272 (.Y(n2678), 
	.B1(n9067), 
	.B0(n9051), 
	.A1(n9050), 
	.A0(n6309));
   INVX1 U5273 (.Y(n9067), 
	.A(\ram[131][0] ));
   NOR2BX1 U5274 (.Y(n9051), 
	.B(n9050), 
	.AN(mem_write_en));
   NAND2X1 U5275 (.Y(n9050), 
	.B(n6457), 
	.A(n8851));
   OAI22X1 U5276 (.Y(n2677), 
	.B1(n9070), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6311));
   INVX1 U5277 (.Y(n9070), 
	.A(\ram[130][15] ));
   OAI22X1 U5278 (.Y(n2676), 
	.B1(n9071), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6314));
   INVX1 U5279 (.Y(n9071), 
	.A(\ram[130][14] ));
   OAI22X1 U5280 (.Y(n2675), 
	.B1(n9072), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6316));
   INVX1 U5281 (.Y(n9072), 
	.A(\ram[130][13] ));
   OAI22X1 U5282 (.Y(n2674), 
	.B1(n9073), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6318));
   INVX1 U5283 (.Y(n9073), 
	.A(\ram[130][12] ));
   OAI22X1 U5284 (.Y(n2673), 
	.B1(n9074), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6320));
   INVX1 U5285 (.Y(n9074), 
	.A(\ram[130][11] ));
   OAI22X1 U5286 (.Y(n2672), 
	.B1(n9075), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6322));
   INVX1 U5287 (.Y(n9075), 
	.A(\ram[130][10] ));
   OAI22X1 U5288 (.Y(n2671), 
	.B1(n9076), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6324));
   INVX1 U5289 (.Y(n9076), 
	.A(\ram[130][9] ));
   OAI22X1 U5290 (.Y(n2670), 
	.B1(n9077), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6326));
   INVX1 U5291 (.Y(n9077), 
	.A(\ram[130][8] ));
   OAI22X1 U5292 (.Y(n2669), 
	.B1(n9078), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6328));
   INVX1 U5293 (.Y(n9078), 
	.A(\ram[130][7] ));
   OAI22X1 U5294 (.Y(n2668), 
	.B1(n9079), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6330));
   INVX1 U5295 (.Y(n9079), 
	.A(\ram[130][6] ));
   OAI22X1 U5296 (.Y(n2667), 
	.B1(n9080), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6332));
   INVX1 U5297 (.Y(n9080), 
	.A(\ram[130][5] ));
   OAI22X1 U5298 (.Y(n2666), 
	.B1(n9081), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6334));
   INVX1 U5299 (.Y(n9081), 
	.A(\ram[130][4] ));
   OAI22X1 U5300 (.Y(n2665), 
	.B1(n9082), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6336));
   INVX1 U5301 (.Y(n9082), 
	.A(\ram[130][3] ));
   OAI22X1 U5302 (.Y(n2664), 
	.B1(n9083), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6338));
   INVX1 U5303 (.Y(n9083), 
	.A(\ram[130][2] ));
   OAI22X1 U5304 (.Y(n2663), 
	.B1(n9084), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6306));
   INVX1 U5305 (.Y(n9084), 
	.A(\ram[130][1] ));
   OAI22X1 U5306 (.Y(n2662), 
	.B1(n9085), 
	.B0(n9069), 
	.A1(n9068), 
	.A0(n6309));
   INVX1 U5307 (.Y(n9085), 
	.A(\ram[130][0] ));
   NOR2BX1 U5308 (.Y(n9069), 
	.B(n9068), 
	.AN(mem_write_en));
   NAND2X1 U5309 (.Y(n9068), 
	.B(n6476), 
	.A(n8851));
   OAI22X1 U5310 (.Y(n2661), 
	.B1(n9088), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6311));
   INVX1 U5311 (.Y(n9088), 
	.A(\ram[129][15] ));
   OAI22X1 U5312 (.Y(n2660), 
	.B1(n9089), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6314));
   INVX1 U5313 (.Y(n9089), 
	.A(\ram[129][14] ));
   OAI22X1 U5314 (.Y(n2659), 
	.B1(n9090), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6316));
   INVX1 U5315 (.Y(n9090), 
	.A(\ram[129][13] ));
   OAI22X1 U5316 (.Y(n2658), 
	.B1(n9091), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6318));
   INVX1 U5317 (.Y(n9091), 
	.A(\ram[129][12] ));
   OAI22X1 U5318 (.Y(n2657), 
	.B1(n9092), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6320));
   INVX1 U5319 (.Y(n9092), 
	.A(\ram[129][11] ));
   OAI22X1 U5320 (.Y(n2656), 
	.B1(n9093), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6322));
   INVX1 U5321 (.Y(n9093), 
	.A(\ram[129][10] ));
   OAI22X1 U5322 (.Y(n2655), 
	.B1(n9094), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6324));
   INVX1 U5323 (.Y(n9094), 
	.A(\ram[129][9] ));
   OAI22X1 U5324 (.Y(n2654), 
	.B1(n9095), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6326));
   INVX1 U5325 (.Y(n9095), 
	.A(\ram[129][8] ));
   OAI22X1 U5326 (.Y(n2653), 
	.B1(n9096), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6328));
   INVX1 U5327 (.Y(n9096), 
	.A(\ram[129][7] ));
   OAI22X1 U5328 (.Y(n2652), 
	.B1(n9097), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6330));
   INVX1 U5329 (.Y(n9097), 
	.A(\ram[129][6] ));
   OAI22X1 U5330 (.Y(n2651), 
	.B1(n9098), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6332));
   INVX1 U5331 (.Y(n9098), 
	.A(\ram[129][5] ));
   OAI22X1 U5332 (.Y(n2650), 
	.B1(n9099), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6334));
   INVX1 U5333 (.Y(n9099), 
	.A(\ram[129][4] ));
   OAI22X1 U5334 (.Y(n2649), 
	.B1(n9100), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6336));
   INVX1 U5335 (.Y(n9100), 
	.A(\ram[129][3] ));
   OAI22X1 U5336 (.Y(n2648), 
	.B1(n9101), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6338));
   INVX1 U5337 (.Y(n9101), 
	.A(\ram[129][2] ));
   OAI22X1 U5338 (.Y(n2647), 
	.B1(n9102), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6306));
   INVX1 U5339 (.Y(n9102), 
	.A(\ram[129][1] ));
   OAI22X1 U5340 (.Y(n2646), 
	.B1(n9103), 
	.B0(n9087), 
	.A1(n9086), 
	.A0(n6309));
   INVX1 U5341 (.Y(n9103), 
	.A(\ram[129][0] ));
   NOR2BX1 U5342 (.Y(n9087), 
	.B(n9086), 
	.AN(mem_write_en));
   NAND2X1 U5343 (.Y(n9086), 
	.B(n6495), 
	.A(n8851));
   OAI22X1 U5344 (.Y(n2645), 
	.B1(n9106), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6311));
   INVX1 U5345 (.Y(n9106), 
	.A(\ram[128][15] ));
   OAI22X1 U5346 (.Y(n2644), 
	.B1(n9107), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6314));
   INVX1 U5347 (.Y(n9107), 
	.A(\ram[128][14] ));
   OAI22X1 U5348 (.Y(n2643), 
	.B1(n9108), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6316));
   INVX1 U5349 (.Y(n9108), 
	.A(\ram[128][13] ));
   OAI22X1 U5350 (.Y(n2642), 
	.B1(n9109), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6318));
   INVX1 U5351 (.Y(n9109), 
	.A(\ram[128][12] ));
   OAI22X1 U5352 (.Y(n2641), 
	.B1(n9110), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6320));
   INVX1 U5353 (.Y(n9110), 
	.A(\ram[128][11] ));
   OAI22X1 U5354 (.Y(n2640), 
	.B1(n9111), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6322));
   INVX1 U5355 (.Y(n9111), 
	.A(\ram[128][10] ));
   OAI22X1 U5356 (.Y(n2639), 
	.B1(n9112), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6324));
   INVX1 U5357 (.Y(n9112), 
	.A(\ram[128][9] ));
   OAI22X1 U5358 (.Y(n2638), 
	.B1(n9113), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6326));
   INVX1 U5359 (.Y(n9113), 
	.A(\ram[128][8] ));
   OAI22X1 U5360 (.Y(n2637), 
	.B1(n9114), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6328));
   INVX1 U5361 (.Y(n9114), 
	.A(\ram[128][7] ));
   OAI22X1 U5362 (.Y(n2636), 
	.B1(n9115), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6330));
   INVX1 U5363 (.Y(n9115), 
	.A(\ram[128][6] ));
   OAI22X1 U5364 (.Y(n2635), 
	.B1(n9116), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6332));
   INVX1 U5365 (.Y(n9116), 
	.A(\ram[128][5] ));
   OAI22X1 U5366 (.Y(n2634), 
	.B1(n9117), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6334));
   INVX1 U5367 (.Y(n9117), 
	.A(\ram[128][4] ));
   OAI22X1 U5368 (.Y(n2633), 
	.B1(n9118), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6336));
   INVX1 U5369 (.Y(n9118), 
	.A(\ram[128][3] ));
   OAI22X1 U5370 (.Y(n2632), 
	.B1(n9119), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6338));
   INVX1 U5371 (.Y(n9119), 
	.A(\ram[128][2] ));
   OAI22X1 U5372 (.Y(n2631), 
	.B1(n9120), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6306));
   INVX1 U5373 (.Y(n9120), 
	.A(\ram[128][1] ));
   OAI22X1 U5374 (.Y(n2630), 
	.B1(n9121), 
	.B0(n9105), 
	.A1(n9104), 
	.A0(n6309));
   INVX1 U5375 (.Y(n9121), 
	.A(\ram[128][0] ));
   NOR2BX1 U5376 (.Y(n9105), 
	.B(n9104), 
	.AN(mem_write_en));
   NAND2X1 U5377 (.Y(n9104), 
	.B(n6514), 
	.A(n8851));
   OAI22X1 U5378 (.Y(n2629), 
	.B1(n9124), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6311));
   INVX1 U5379 (.Y(n9124), 
	.A(\ram[127][15] ));
   OAI22X1 U5380 (.Y(n2628), 
	.B1(n9125), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6314));
   INVX1 U5381 (.Y(n9125), 
	.A(\ram[127][14] ));
   OAI22X1 U5382 (.Y(n2627), 
	.B1(n9126), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6316));
   INVX1 U5383 (.Y(n9126), 
	.A(\ram[127][13] ));
   OAI22X1 U5384 (.Y(n2626), 
	.B1(n9127), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6318));
   INVX1 U5385 (.Y(n9127), 
	.A(\ram[127][12] ));
   OAI22X1 U5386 (.Y(n2625), 
	.B1(n9128), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6320));
   INVX1 U5387 (.Y(n9128), 
	.A(\ram[127][11] ));
   OAI22X1 U5388 (.Y(n2624), 
	.B1(n9129), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6322));
   INVX1 U5389 (.Y(n9129), 
	.A(\ram[127][10] ));
   OAI22X1 U5390 (.Y(n2623), 
	.B1(n9130), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6324));
   INVX1 U5391 (.Y(n9130), 
	.A(\ram[127][9] ));
   OAI22X1 U5392 (.Y(n2622), 
	.B1(n9131), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6326));
   INVX1 U5393 (.Y(n9131), 
	.A(\ram[127][8] ));
   OAI22X1 U5394 (.Y(n2621), 
	.B1(n9132), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6328));
   INVX1 U5395 (.Y(n9132), 
	.A(\ram[127][7] ));
   OAI22X1 U5396 (.Y(n2620), 
	.B1(n9133), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6330));
   INVX1 U5397 (.Y(n9133), 
	.A(\ram[127][6] ));
   OAI22X1 U5398 (.Y(n2619), 
	.B1(n9134), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6332));
   INVX1 U5399 (.Y(n9134), 
	.A(\ram[127][5] ));
   OAI22X1 U5400 (.Y(n2618), 
	.B1(n9135), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6334));
   INVX1 U5401 (.Y(n9135), 
	.A(\ram[127][4] ));
   OAI22X1 U5402 (.Y(n2617), 
	.B1(n9136), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6336));
   INVX1 U5403 (.Y(n9136), 
	.A(\ram[127][3] ));
   OAI22X1 U5404 (.Y(n2616), 
	.B1(n9137), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6338));
   INVX1 U5405 (.Y(n9137), 
	.A(\ram[127][2] ));
   OAI22X1 U5406 (.Y(n2615), 
	.B1(n9138), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6306));
   INVX1 U5407 (.Y(n9138), 
	.A(\ram[127][1] ));
   OAI22X1 U5408 (.Y(n2614), 
	.B1(n9139), 
	.B0(n9123), 
	.A1(n9122), 
	.A0(n6309));
   INVX1 U5409 (.Y(n9139), 
	.A(\ram[127][0] ));
   NOR2BX1 U5410 (.Y(n9123), 
	.B(n9122), 
	.AN(mem_write_en));
   NAND2X1 U5411 (.Y(n9122), 
	.B(n6533), 
	.A(n9140));
   OAI22X1 U5412 (.Y(n2613), 
	.B1(n9143), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6311));
   INVX1 U5413 (.Y(n9143), 
	.A(\ram[126][15] ));
   OAI22X1 U5414 (.Y(n2612), 
	.B1(n9144), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6314));
   INVX1 U5415 (.Y(n9144), 
	.A(\ram[126][14] ));
   OAI22X1 U5416 (.Y(n2611), 
	.B1(n9145), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6316));
   INVX1 U5417 (.Y(n9145), 
	.A(\ram[126][13] ));
   OAI22X1 U5418 (.Y(n2610), 
	.B1(n9146), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6318));
   INVX1 U5419 (.Y(n9146), 
	.A(\ram[126][12] ));
   OAI22X1 U5420 (.Y(n2609), 
	.B1(n9147), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6320));
   INVX1 U5421 (.Y(n9147), 
	.A(\ram[126][11] ));
   OAI22X1 U5422 (.Y(n2608), 
	.B1(n9148), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6322));
   INVX1 U5423 (.Y(n9148), 
	.A(\ram[126][10] ));
   OAI22X1 U5424 (.Y(n2607), 
	.B1(n9149), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6324));
   INVX1 U5425 (.Y(n9149), 
	.A(\ram[126][9] ));
   OAI22X1 U5426 (.Y(n2606), 
	.B1(n9150), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6326));
   INVX1 U5427 (.Y(n9150), 
	.A(\ram[126][8] ));
   OAI22X1 U5428 (.Y(n2605), 
	.B1(n9151), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6328));
   INVX1 U5429 (.Y(n9151), 
	.A(\ram[126][7] ));
   OAI22X1 U5430 (.Y(n2604), 
	.B1(n9152), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6330));
   INVX1 U5431 (.Y(n9152), 
	.A(\ram[126][6] ));
   OAI22X1 U5432 (.Y(n2603), 
	.B1(n9153), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6332));
   INVX1 U5433 (.Y(n9153), 
	.A(\ram[126][5] ));
   OAI22X1 U5434 (.Y(n2602), 
	.B1(n9154), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6334));
   INVX1 U5435 (.Y(n9154), 
	.A(\ram[126][4] ));
   OAI22X1 U5436 (.Y(n2601), 
	.B1(n9155), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6336));
   INVX1 U5437 (.Y(n9155), 
	.A(\ram[126][3] ));
   OAI22X1 U5438 (.Y(n2600), 
	.B1(n9156), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6338));
   INVX1 U5439 (.Y(n9156), 
	.A(\ram[126][2] ));
   OAI22X1 U5440 (.Y(n2599), 
	.B1(n9157), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6306));
   INVX1 U5441 (.Y(n9157), 
	.A(\ram[126][1] ));
   OAI22X1 U5442 (.Y(n2598), 
	.B1(n9158), 
	.B0(n9142), 
	.A1(n9141), 
	.A0(n6309));
   INVX1 U5443 (.Y(n9158), 
	.A(\ram[126][0] ));
   NOR2BX1 U5444 (.Y(n9142), 
	.B(n9141), 
	.AN(mem_write_en));
   NAND2X1 U5445 (.Y(n9141), 
	.B(n6553), 
	.A(n9140));
   OAI22X1 U5446 (.Y(n2597), 
	.B1(n9161), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6311));
   INVX1 U5447 (.Y(n9161), 
	.A(\ram[125][15] ));
   OAI22X1 U5448 (.Y(n2596), 
	.B1(n9162), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6314));
   INVX1 U5449 (.Y(n9162), 
	.A(\ram[125][14] ));
   OAI22X1 U5450 (.Y(n2595), 
	.B1(n9163), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6316));
   INVX1 U5451 (.Y(n9163), 
	.A(\ram[125][13] ));
   OAI22X1 U5452 (.Y(n2594), 
	.B1(n9164), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6318));
   INVX1 U5453 (.Y(n9164), 
	.A(\ram[125][12] ));
   OAI22X1 U5454 (.Y(n2593), 
	.B1(n9165), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6320));
   INVX1 U5455 (.Y(n9165), 
	.A(\ram[125][11] ));
   OAI22X1 U5456 (.Y(n2592), 
	.B1(n9166), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6322));
   INVX1 U5457 (.Y(n9166), 
	.A(\ram[125][10] ));
   OAI22X1 U5458 (.Y(n2591), 
	.B1(n9167), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6324));
   INVX1 U5459 (.Y(n9167), 
	.A(\ram[125][9] ));
   OAI22X1 U5460 (.Y(n2590), 
	.B1(n9168), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6326));
   INVX1 U5461 (.Y(n9168), 
	.A(\ram[125][8] ));
   OAI22X1 U5462 (.Y(n2589), 
	.B1(n9169), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6328));
   INVX1 U5463 (.Y(n9169), 
	.A(\ram[125][7] ));
   OAI22X1 U5464 (.Y(n2588), 
	.B1(n9170), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6330));
   INVX1 U5465 (.Y(n9170), 
	.A(\ram[125][6] ));
   OAI22X1 U5466 (.Y(n2587), 
	.B1(n9171), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6332));
   INVX1 U5467 (.Y(n9171), 
	.A(\ram[125][5] ));
   OAI22X1 U5468 (.Y(n2586), 
	.B1(n9172), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6334));
   INVX1 U5469 (.Y(n9172), 
	.A(\ram[125][4] ));
   OAI22X1 U5470 (.Y(n2585), 
	.B1(n9173), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6336));
   INVX1 U5471 (.Y(n9173), 
	.A(\ram[125][3] ));
   OAI22X1 U5472 (.Y(n2584), 
	.B1(n9174), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6338));
   INVX1 U5473 (.Y(n9174), 
	.A(\ram[125][2] ));
   OAI22X1 U5474 (.Y(n2583), 
	.B1(n9175), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6306));
   INVX1 U5475 (.Y(n9175), 
	.A(\ram[125][1] ));
   OAI22X1 U5476 (.Y(n2582), 
	.B1(n9176), 
	.B0(n9160), 
	.A1(n9159), 
	.A0(n6309));
   INVX1 U5477 (.Y(n9176), 
	.A(\ram[125][0] ));
   NOR2BX1 U5478 (.Y(n9160), 
	.B(n9159), 
	.AN(mem_write_en));
   NAND2X1 U5479 (.Y(n9159), 
	.B(n6572), 
	.A(n9140));
   OAI22X1 U5480 (.Y(n2581), 
	.B1(n9179), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6311));
   INVX1 U5481 (.Y(n9179), 
	.A(\ram[124][15] ));
   OAI22X1 U5482 (.Y(n2580), 
	.B1(n9180), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6314));
   INVX1 U5483 (.Y(n9180), 
	.A(\ram[124][14] ));
   OAI22X1 U5484 (.Y(n2579), 
	.B1(n9181), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6316));
   INVX1 U5485 (.Y(n9181), 
	.A(\ram[124][13] ));
   OAI22X1 U5486 (.Y(n2578), 
	.B1(n9182), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6318));
   INVX1 U5487 (.Y(n9182), 
	.A(\ram[124][12] ));
   OAI22X1 U5488 (.Y(n2577), 
	.B1(n9183), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6320));
   INVX1 U5489 (.Y(n9183), 
	.A(\ram[124][11] ));
   OAI22X1 U5490 (.Y(n2576), 
	.B1(n9184), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6322));
   INVX1 U5491 (.Y(n9184), 
	.A(\ram[124][10] ));
   OAI22X1 U5492 (.Y(n2575), 
	.B1(n9185), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6324));
   INVX1 U5493 (.Y(n9185), 
	.A(\ram[124][9] ));
   OAI22X1 U5494 (.Y(n2574), 
	.B1(n9186), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6326));
   INVX1 U5495 (.Y(n9186), 
	.A(\ram[124][8] ));
   OAI22X1 U5496 (.Y(n2573), 
	.B1(n9187), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6328));
   INVX1 U5497 (.Y(n9187), 
	.A(\ram[124][7] ));
   OAI22X1 U5498 (.Y(n2572), 
	.B1(n9188), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6330));
   INVX1 U5499 (.Y(n9188), 
	.A(\ram[124][6] ));
   OAI22X1 U5500 (.Y(n2571), 
	.B1(n9189), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6332));
   INVX1 U5501 (.Y(n9189), 
	.A(\ram[124][5] ));
   OAI22X1 U5502 (.Y(n2570), 
	.B1(n9190), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6334));
   INVX1 U5503 (.Y(n9190), 
	.A(\ram[124][4] ));
   OAI22X1 U5504 (.Y(n2569), 
	.B1(n9191), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6336));
   INVX1 U5505 (.Y(n9191), 
	.A(\ram[124][3] ));
   OAI22X1 U5506 (.Y(n2568), 
	.B1(n9192), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6338));
   INVX1 U5507 (.Y(n9192), 
	.A(\ram[124][2] ));
   OAI22X1 U5508 (.Y(n2567), 
	.B1(n9193), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6306));
   INVX1 U5509 (.Y(n9193), 
	.A(\ram[124][1] ));
   OAI22X1 U5510 (.Y(n2566), 
	.B1(n9194), 
	.B0(n9178), 
	.A1(n9177), 
	.A0(n6309));
   INVX1 U5511 (.Y(n9194), 
	.A(\ram[124][0] ));
   NOR2BX1 U5512 (.Y(n9178), 
	.B(n9177), 
	.AN(mem_write_en));
   NAND2X1 U5513 (.Y(n9177), 
	.B(n6591), 
	.A(n9140));
   OAI22X1 U5514 (.Y(n2565), 
	.B1(n9197), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6311));
   INVX1 U5515 (.Y(n9197), 
	.A(\ram[123][15] ));
   OAI22X1 U5516 (.Y(n2564), 
	.B1(n9198), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6314));
   INVX1 U5517 (.Y(n9198), 
	.A(\ram[123][14] ));
   OAI22X1 U5518 (.Y(n2563), 
	.B1(n9199), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6316));
   INVX1 U5519 (.Y(n9199), 
	.A(\ram[123][13] ));
   OAI22X1 U5520 (.Y(n2562), 
	.B1(n9200), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6318));
   INVX1 U5521 (.Y(n9200), 
	.A(\ram[123][12] ));
   OAI22X1 U5522 (.Y(n2561), 
	.B1(n9201), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6320));
   INVX1 U5523 (.Y(n9201), 
	.A(\ram[123][11] ));
   OAI22X1 U5524 (.Y(n2560), 
	.B1(n9202), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6322));
   INVX1 U5525 (.Y(n9202), 
	.A(\ram[123][10] ));
   OAI22X1 U5526 (.Y(n2559), 
	.B1(n9203), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6324));
   INVX1 U5527 (.Y(n9203), 
	.A(\ram[123][9] ));
   OAI22X1 U5528 (.Y(n2558), 
	.B1(n9204), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6326));
   INVX1 U5529 (.Y(n9204), 
	.A(\ram[123][8] ));
   OAI22X1 U5530 (.Y(n2557), 
	.B1(n9205), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6328));
   INVX1 U5531 (.Y(n9205), 
	.A(\ram[123][7] ));
   OAI22X1 U5532 (.Y(n2556), 
	.B1(n9206), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6330));
   INVX1 U5533 (.Y(n9206), 
	.A(\ram[123][6] ));
   OAI22X1 U5534 (.Y(n2555), 
	.B1(n9207), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6332));
   INVX1 U5535 (.Y(n9207), 
	.A(\ram[123][5] ));
   OAI22X1 U5536 (.Y(n2554), 
	.B1(n9208), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6334));
   INVX1 U5537 (.Y(n9208), 
	.A(\ram[123][4] ));
   OAI22X1 U5538 (.Y(n2553), 
	.B1(n9209), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6336));
   INVX1 U5539 (.Y(n9209), 
	.A(\ram[123][3] ));
   OAI22X1 U5540 (.Y(n2552), 
	.B1(n9210), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6338));
   INVX1 U5541 (.Y(n9210), 
	.A(\ram[123][2] ));
   OAI22X1 U5542 (.Y(n2551), 
	.B1(n9211), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6306));
   INVX1 U5543 (.Y(n9211), 
	.A(\ram[123][1] ));
   OAI22X1 U5544 (.Y(n2550), 
	.B1(n9212), 
	.B0(n9196), 
	.A1(n9195), 
	.A0(n6309));
   INVX1 U5545 (.Y(n9212), 
	.A(\ram[123][0] ));
   NOR2BX1 U5546 (.Y(n9196), 
	.B(n9195), 
	.AN(mem_write_en));
   NAND2X1 U5547 (.Y(n9195), 
	.B(n6610), 
	.A(n9140));
   OAI22X1 U5548 (.Y(n2549), 
	.B1(n9215), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6311));
   INVX1 U5549 (.Y(n9215), 
	.A(\ram[122][15] ));
   OAI22X1 U5550 (.Y(n2548), 
	.B1(n9216), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6314));
   INVX1 U5551 (.Y(n9216), 
	.A(\ram[122][14] ));
   OAI22X1 U5552 (.Y(n2547), 
	.B1(n9217), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6316));
   INVX1 U5553 (.Y(n9217), 
	.A(\ram[122][13] ));
   OAI22X1 U5554 (.Y(n2546), 
	.B1(n9218), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6318));
   INVX1 U5555 (.Y(n9218), 
	.A(\ram[122][12] ));
   OAI22X1 U5556 (.Y(n2545), 
	.B1(n9219), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6320));
   INVX1 U5557 (.Y(n9219), 
	.A(\ram[122][11] ));
   OAI22X1 U5558 (.Y(n2544), 
	.B1(n9220), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6322));
   INVX1 U5559 (.Y(n9220), 
	.A(\ram[122][10] ));
   OAI22X1 U5560 (.Y(n2543), 
	.B1(n9221), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6324));
   INVX1 U5561 (.Y(n9221), 
	.A(\ram[122][9] ));
   OAI22X1 U5562 (.Y(n2542), 
	.B1(n9222), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6326));
   INVX1 U5563 (.Y(n9222), 
	.A(\ram[122][8] ));
   OAI22X1 U5564 (.Y(n2541), 
	.B1(n9223), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6328));
   INVX1 U5565 (.Y(n9223), 
	.A(\ram[122][7] ));
   OAI22X1 U5566 (.Y(n2540), 
	.B1(n9224), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6330));
   INVX1 U5567 (.Y(n9224), 
	.A(\ram[122][6] ));
   OAI22X1 U5568 (.Y(n2539), 
	.B1(n9225), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6332));
   INVX1 U5569 (.Y(n9225), 
	.A(\ram[122][5] ));
   OAI22X1 U5570 (.Y(n2538), 
	.B1(n9226), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6334));
   INVX1 U5571 (.Y(n9226), 
	.A(\ram[122][4] ));
   OAI22X1 U5572 (.Y(n2537), 
	.B1(n9227), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6336));
   INVX1 U5573 (.Y(n9227), 
	.A(\ram[122][3] ));
   OAI22X1 U5574 (.Y(n2536), 
	.B1(n9228), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6338));
   INVX1 U5575 (.Y(n9228), 
	.A(\ram[122][2] ));
   OAI22X1 U5576 (.Y(n2535), 
	.B1(n9229), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6306));
   INVX1 U5577 (.Y(n9229), 
	.A(\ram[122][1] ));
   OAI22X1 U5578 (.Y(n2534), 
	.B1(n9230), 
	.B0(n9214), 
	.A1(n9213), 
	.A0(n6309));
   INVX1 U5579 (.Y(n9230), 
	.A(\ram[122][0] ));
   NOR2BX1 U5580 (.Y(n9214), 
	.B(n9213), 
	.AN(mem_write_en));
   NAND2X1 U5581 (.Y(n9213), 
	.B(n6629), 
	.A(n9140));
   OAI22X1 U5582 (.Y(n2533), 
	.B1(n9233), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6311));
   INVX1 U5583 (.Y(n9233), 
	.A(\ram[121][15] ));
   OAI22X1 U5584 (.Y(n2532), 
	.B1(n9234), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6314));
   INVX1 U5585 (.Y(n9234), 
	.A(\ram[121][14] ));
   OAI22X1 U5586 (.Y(n2531), 
	.B1(n9235), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6316));
   INVX1 U5587 (.Y(n9235), 
	.A(\ram[121][13] ));
   OAI22X1 U5588 (.Y(n2530), 
	.B1(n9236), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6318));
   INVX1 U5589 (.Y(n9236), 
	.A(\ram[121][12] ));
   OAI22X1 U5590 (.Y(n2529), 
	.B1(n9237), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6320));
   INVX1 U5591 (.Y(n9237), 
	.A(\ram[121][11] ));
   OAI22X1 U5592 (.Y(n2528), 
	.B1(n9238), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6322));
   INVX1 U5593 (.Y(n9238), 
	.A(\ram[121][10] ));
   OAI22X1 U5594 (.Y(n2527), 
	.B1(n9239), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6324));
   INVX1 U5595 (.Y(n9239), 
	.A(\ram[121][9] ));
   OAI22X1 U5596 (.Y(n2526), 
	.B1(n9240), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6326));
   INVX1 U5597 (.Y(n9240), 
	.A(\ram[121][8] ));
   OAI22X1 U5598 (.Y(n2525), 
	.B1(n9241), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6328));
   INVX1 U5599 (.Y(n9241), 
	.A(\ram[121][7] ));
   OAI22X1 U5600 (.Y(n2524), 
	.B1(n9242), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6330));
   INVX1 U5601 (.Y(n9242), 
	.A(\ram[121][6] ));
   OAI22X1 U5602 (.Y(n2523), 
	.B1(n9243), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6332));
   INVX1 U5603 (.Y(n9243), 
	.A(\ram[121][5] ));
   OAI22X1 U5604 (.Y(n2522), 
	.B1(n9244), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6334));
   INVX1 U5605 (.Y(n9244), 
	.A(\ram[121][4] ));
   OAI22X1 U5606 (.Y(n2521), 
	.B1(n9245), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6336));
   INVX1 U5607 (.Y(n9245), 
	.A(\ram[121][3] ));
   OAI22X1 U5608 (.Y(n2520), 
	.B1(n9246), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6338));
   INVX1 U5609 (.Y(n9246), 
	.A(\ram[121][2] ));
   OAI22X1 U5610 (.Y(n2519), 
	.B1(n9247), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6306));
   INVX1 U5611 (.Y(n9247), 
	.A(\ram[121][1] ));
   OAI22X1 U5612 (.Y(n2518), 
	.B1(n9248), 
	.B0(n9232), 
	.A1(n9231), 
	.A0(n6309));
   INVX1 U5613 (.Y(n9248), 
	.A(\ram[121][0] ));
   NOR2BX1 U5614 (.Y(n9232), 
	.B(n9231), 
	.AN(mem_write_en));
   NAND2X1 U5615 (.Y(n9231), 
	.B(n6342), 
	.A(n9140));
   OAI22X1 U5616 (.Y(n2517), 
	.B1(n9251), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6311));
   INVX1 U5617 (.Y(n9251), 
	.A(\ram[120][15] ));
   OAI22X1 U5618 (.Y(n2516), 
	.B1(n9252), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6314));
   INVX1 U5619 (.Y(n9252), 
	.A(\ram[120][14] ));
   OAI22X1 U5620 (.Y(n2515), 
	.B1(n9253), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6316));
   INVX1 U5621 (.Y(n9253), 
	.A(\ram[120][13] ));
   OAI22X1 U5622 (.Y(n2514), 
	.B1(n9254), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6318));
   INVX1 U5623 (.Y(n9254), 
	.A(\ram[120][12] ));
   OAI22X1 U5624 (.Y(n2513), 
	.B1(n9255), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6320));
   INVX1 U5625 (.Y(n9255), 
	.A(\ram[120][11] ));
   OAI22X1 U5626 (.Y(n2512), 
	.B1(n9256), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6322));
   INVX1 U5627 (.Y(n9256), 
	.A(\ram[120][10] ));
   OAI22X1 U5628 (.Y(n2511), 
	.B1(n9257), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6324));
   INVX1 U5629 (.Y(n9257), 
	.A(\ram[120][9] ));
   OAI22X1 U5630 (.Y(n2510), 
	.B1(n9258), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6326));
   INVX1 U5631 (.Y(n9258), 
	.A(\ram[120][8] ));
   OAI22X1 U5632 (.Y(n2509), 
	.B1(n9259), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6328));
   INVX1 U5633 (.Y(n9259), 
	.A(\ram[120][7] ));
   OAI22X1 U5634 (.Y(n2508), 
	.B1(n9260), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6330));
   INVX1 U5635 (.Y(n9260), 
	.A(\ram[120][6] ));
   OAI22X1 U5636 (.Y(n2507), 
	.B1(n9261), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6332));
   INVX1 U5637 (.Y(n9261), 
	.A(\ram[120][5] ));
   OAI22X1 U5638 (.Y(n2506), 
	.B1(n9262), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6334));
   INVX1 U5639 (.Y(n9262), 
	.A(\ram[120][4] ));
   OAI22X1 U5640 (.Y(n2505), 
	.B1(n9263), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6336));
   INVX1 U5641 (.Y(n9263), 
	.A(\ram[120][3] ));
   OAI22X1 U5642 (.Y(n2504), 
	.B1(n9264), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6338));
   INVX1 U5643 (.Y(n9264), 
	.A(\ram[120][2] ));
   OAI22X1 U5644 (.Y(n2503), 
	.B1(n9265), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6306));
   INVX1 U5645 (.Y(n9265), 
	.A(\ram[120][1] ));
   OAI22X1 U5646 (.Y(n2502), 
	.B1(n9266), 
	.B0(n9250), 
	.A1(n9249), 
	.A0(n6309));
   INVX1 U5647 (.Y(n9266), 
	.A(\ram[120][0] ));
   NOR2BX1 U5648 (.Y(n9250), 
	.B(n9249), 
	.AN(mem_write_en));
   NAND2X1 U5649 (.Y(n9249), 
	.B(n6362), 
	.A(n9140));
   OAI22X1 U5650 (.Y(n2501), 
	.B1(n9269), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6311));
   INVX1 U5651 (.Y(n9269), 
	.A(\ram[119][15] ));
   OAI22X1 U5652 (.Y(n2500), 
	.B1(n9270), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6314));
   INVX1 U5653 (.Y(n9270), 
	.A(\ram[119][14] ));
   OAI22X1 U5654 (.Y(n2499), 
	.B1(n9271), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6316));
   INVX1 U5655 (.Y(n9271), 
	.A(\ram[119][13] ));
   OAI22X1 U5656 (.Y(n2498), 
	.B1(n9272), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6318));
   INVX1 U5657 (.Y(n9272), 
	.A(\ram[119][12] ));
   OAI22X1 U5658 (.Y(n2497), 
	.B1(n9273), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6320));
   INVX1 U5659 (.Y(n9273), 
	.A(\ram[119][11] ));
   OAI22X1 U5660 (.Y(n2496), 
	.B1(n9274), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6322));
   INVX1 U5661 (.Y(n9274), 
	.A(\ram[119][10] ));
   OAI22X1 U5662 (.Y(n2495), 
	.B1(n9275), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6324));
   INVX1 U5663 (.Y(n9275), 
	.A(\ram[119][9] ));
   OAI22X1 U5664 (.Y(n2494), 
	.B1(n9276), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6326));
   INVX1 U5665 (.Y(n9276), 
	.A(\ram[119][8] ));
   OAI22X1 U5666 (.Y(n2493), 
	.B1(n9277), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6328));
   INVX1 U5667 (.Y(n9277), 
	.A(\ram[119][7] ));
   OAI22X1 U5668 (.Y(n2492), 
	.B1(n9278), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6330));
   INVX1 U5669 (.Y(n9278), 
	.A(\ram[119][6] ));
   OAI22X1 U5670 (.Y(n2491), 
	.B1(n9279), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6332));
   INVX1 U5671 (.Y(n9279), 
	.A(\ram[119][5] ));
   OAI22X1 U5672 (.Y(n2490), 
	.B1(n9280), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6334));
   INVX1 U5673 (.Y(n9280), 
	.A(\ram[119][4] ));
   OAI22X1 U5674 (.Y(n2489), 
	.B1(n9281), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6336));
   INVX1 U5675 (.Y(n9281), 
	.A(\ram[119][3] ));
   OAI22X1 U5676 (.Y(n2488), 
	.B1(n9282), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6338));
   INVX1 U5677 (.Y(n9282), 
	.A(\ram[119][2] ));
   OAI22X1 U5678 (.Y(n2487), 
	.B1(n9283), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6306));
   INVX1 U5679 (.Y(n9283), 
	.A(\ram[119][1] ));
   OAI22X1 U5680 (.Y(n2486), 
	.B1(n9284), 
	.B0(n9268), 
	.A1(n9267), 
	.A0(n6309));
   INVX1 U5681 (.Y(n9284), 
	.A(\ram[119][0] ));
   NOR2BX1 U5682 (.Y(n9268), 
	.B(n9267), 
	.AN(mem_write_en));
   NAND2X1 U5683 (.Y(n9267), 
	.B(n6381), 
	.A(n9140));
   OAI22X1 U5684 (.Y(n2485), 
	.B1(n9287), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6311));
   INVX1 U5685 (.Y(n9287), 
	.A(\ram[118][15] ));
   OAI22X1 U5686 (.Y(n2484), 
	.B1(n9288), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6314));
   INVX1 U5687 (.Y(n9288), 
	.A(\ram[118][14] ));
   OAI22X1 U5688 (.Y(n2483), 
	.B1(n9289), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6316));
   INVX1 U5689 (.Y(n9289), 
	.A(\ram[118][13] ));
   OAI22X1 U5690 (.Y(n2482), 
	.B1(n9290), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6318));
   INVX1 U5691 (.Y(n9290), 
	.A(\ram[118][12] ));
   OAI22X1 U5692 (.Y(n2481), 
	.B1(n9291), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6320));
   INVX1 U5693 (.Y(n9291), 
	.A(\ram[118][11] ));
   OAI22X1 U5694 (.Y(n2480), 
	.B1(n9292), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6322));
   INVX1 U5695 (.Y(n9292), 
	.A(\ram[118][10] ));
   OAI22X1 U5696 (.Y(n2479), 
	.B1(n9293), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6324));
   INVX1 U5697 (.Y(n9293), 
	.A(\ram[118][9] ));
   OAI22X1 U5698 (.Y(n2478), 
	.B1(n9294), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6326));
   INVX1 U5699 (.Y(n9294), 
	.A(\ram[118][8] ));
   OAI22X1 U5700 (.Y(n2477), 
	.B1(n9295), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6328));
   INVX1 U5701 (.Y(n9295), 
	.A(\ram[118][7] ));
   OAI22X1 U5702 (.Y(n2476), 
	.B1(n9296), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6330));
   INVX1 U5703 (.Y(n9296), 
	.A(\ram[118][6] ));
   OAI22X1 U5704 (.Y(n2475), 
	.B1(n9297), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6332));
   INVX1 U5705 (.Y(n9297), 
	.A(\ram[118][5] ));
   OAI22X1 U5706 (.Y(n2474), 
	.B1(n9298), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6334));
   INVX1 U5707 (.Y(n9298), 
	.A(\ram[118][4] ));
   OAI22X1 U5708 (.Y(n2473), 
	.B1(n9299), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6336));
   INVX1 U5709 (.Y(n9299), 
	.A(\ram[118][3] ));
   OAI22X1 U5710 (.Y(n2472), 
	.B1(n9300), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6338));
   INVX1 U5711 (.Y(n9300), 
	.A(\ram[118][2] ));
   OAI22X1 U5712 (.Y(n2471), 
	.B1(n9301), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6306));
   INVX1 U5713 (.Y(n9301), 
	.A(\ram[118][1] ));
   OAI22X1 U5714 (.Y(n2470), 
	.B1(n9302), 
	.B0(n9286), 
	.A1(n9285), 
	.A0(n6309));
   INVX1 U5715 (.Y(n9302), 
	.A(\ram[118][0] ));
   NOR2BX1 U5716 (.Y(n9286), 
	.B(n9285), 
	.AN(mem_write_en));
   NAND2X1 U5717 (.Y(n9285), 
	.B(n6400), 
	.A(n9140));
   OAI22X1 U5718 (.Y(n2469), 
	.B1(n9305), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6311));
   INVX1 U5719 (.Y(n9305), 
	.A(\ram[117][15] ));
   OAI22X1 U5720 (.Y(n2468), 
	.B1(n9306), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6314));
   INVX1 U5721 (.Y(n9306), 
	.A(\ram[117][14] ));
   OAI22X1 U5722 (.Y(n2467), 
	.B1(n9307), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6316));
   INVX1 U5723 (.Y(n9307), 
	.A(\ram[117][13] ));
   OAI22X1 U5724 (.Y(n2466), 
	.B1(n9308), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6318));
   INVX1 U5725 (.Y(n9308), 
	.A(\ram[117][12] ));
   OAI22X1 U5726 (.Y(n2465), 
	.B1(n9309), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6320));
   INVX1 U5727 (.Y(n9309), 
	.A(\ram[117][11] ));
   OAI22X1 U5728 (.Y(n2464), 
	.B1(n9310), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6322));
   INVX1 U5729 (.Y(n9310), 
	.A(\ram[117][10] ));
   OAI22X1 U5730 (.Y(n2463), 
	.B1(n9311), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6324));
   INVX1 U5731 (.Y(n9311), 
	.A(\ram[117][9] ));
   OAI22X1 U5732 (.Y(n2462), 
	.B1(n9312), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6326));
   INVX1 U5733 (.Y(n9312), 
	.A(\ram[117][8] ));
   OAI22X1 U5734 (.Y(n2461), 
	.B1(n9313), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6328));
   INVX1 U5735 (.Y(n9313), 
	.A(\ram[117][7] ));
   OAI22X1 U5736 (.Y(n2460), 
	.B1(n9314), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6330));
   INVX1 U5737 (.Y(n9314), 
	.A(\ram[117][6] ));
   OAI22X1 U5738 (.Y(n2459), 
	.B1(n9315), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6332));
   INVX1 U5739 (.Y(n9315), 
	.A(\ram[117][5] ));
   OAI22X1 U5740 (.Y(n2458), 
	.B1(n9316), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6334));
   INVX1 U5741 (.Y(n9316), 
	.A(\ram[117][4] ));
   OAI22X1 U5742 (.Y(n2457), 
	.B1(n9317), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6336));
   INVX1 U5743 (.Y(n9317), 
	.A(\ram[117][3] ));
   OAI22X1 U5744 (.Y(n2456), 
	.B1(n9318), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6338));
   INVX1 U5745 (.Y(n9318), 
	.A(\ram[117][2] ));
   OAI22X1 U5746 (.Y(n2455), 
	.B1(n9319), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6306));
   INVX1 U5747 (.Y(n9319), 
	.A(\ram[117][1] ));
   OAI22X1 U5748 (.Y(n2454), 
	.B1(n9320), 
	.B0(n9304), 
	.A1(n9303), 
	.A0(n6309));
   INVX1 U5749 (.Y(n9320), 
	.A(\ram[117][0] ));
   NOR2BX1 U5750 (.Y(n9304), 
	.B(n9303), 
	.AN(mem_write_en));
   NAND2X1 U5751 (.Y(n9303), 
	.B(n6419), 
	.A(n9140));
   OAI22X1 U5752 (.Y(n2453), 
	.B1(n9323), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6311));
   INVX1 U5753 (.Y(n9323), 
	.A(\ram[116][15] ));
   OAI22X1 U5754 (.Y(n2452), 
	.B1(n9324), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6314));
   INVX1 U5755 (.Y(n9324), 
	.A(\ram[116][14] ));
   OAI22X1 U5756 (.Y(n2451), 
	.B1(n9325), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6316));
   INVX1 U5757 (.Y(n9325), 
	.A(\ram[116][13] ));
   OAI22X1 U5758 (.Y(n2450), 
	.B1(n9326), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6318));
   INVX1 U5759 (.Y(n9326), 
	.A(\ram[116][12] ));
   OAI22X1 U5760 (.Y(n2449), 
	.B1(n9327), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6320));
   INVX1 U5761 (.Y(n9327), 
	.A(\ram[116][11] ));
   OAI22X1 U5762 (.Y(n2448), 
	.B1(n9328), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6322));
   INVX1 U5763 (.Y(n9328), 
	.A(\ram[116][10] ));
   OAI22X1 U5764 (.Y(n2447), 
	.B1(n9329), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6324));
   INVX1 U5765 (.Y(n9329), 
	.A(\ram[116][9] ));
   OAI22X1 U5766 (.Y(n2446), 
	.B1(n9330), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6326));
   INVX1 U5767 (.Y(n9330), 
	.A(\ram[116][8] ));
   OAI22X1 U5768 (.Y(n2445), 
	.B1(n9331), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6328));
   INVX1 U5769 (.Y(n9331), 
	.A(\ram[116][7] ));
   OAI22X1 U5770 (.Y(n2444), 
	.B1(n9332), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6330));
   INVX1 U5771 (.Y(n9332), 
	.A(\ram[116][6] ));
   OAI22X1 U5772 (.Y(n2443), 
	.B1(n9333), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6332));
   INVX1 U5773 (.Y(n9333), 
	.A(\ram[116][5] ));
   OAI22X1 U5774 (.Y(n2442), 
	.B1(n9334), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6334));
   INVX1 U5775 (.Y(n9334), 
	.A(\ram[116][4] ));
   OAI22X1 U5776 (.Y(n2441), 
	.B1(n9335), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6336));
   INVX1 U5777 (.Y(n9335), 
	.A(\ram[116][3] ));
   OAI22X1 U5778 (.Y(n2440), 
	.B1(n9336), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6338));
   INVX1 U5779 (.Y(n9336), 
	.A(\ram[116][2] ));
   OAI22X1 U5780 (.Y(n2439), 
	.B1(n9337), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6306));
   INVX1 U5781 (.Y(n9337), 
	.A(\ram[116][1] ));
   OAI22X1 U5782 (.Y(n2438), 
	.B1(n9338), 
	.B0(n9322), 
	.A1(n9321), 
	.A0(n6309));
   INVX1 U5783 (.Y(n9338), 
	.A(\ram[116][0] ));
   NOR2BX1 U5784 (.Y(n9322), 
	.B(n9321), 
	.AN(mem_write_en));
   NAND2X1 U5785 (.Y(n9321), 
	.B(n6438), 
	.A(n9140));
   OAI22X1 U5786 (.Y(n2437), 
	.B1(n9341), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6311));
   INVX1 U5787 (.Y(n9341), 
	.A(\ram[115][15] ));
   OAI22X1 U5788 (.Y(n2436), 
	.B1(n9342), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6314));
   INVX1 U5789 (.Y(n9342), 
	.A(\ram[115][14] ));
   OAI22X1 U5790 (.Y(n2435), 
	.B1(n9343), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6316));
   INVX1 U5791 (.Y(n9343), 
	.A(\ram[115][13] ));
   OAI22X1 U5792 (.Y(n2434), 
	.B1(n9344), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6318));
   INVX1 U5793 (.Y(n9344), 
	.A(\ram[115][12] ));
   OAI22X1 U5794 (.Y(n2433), 
	.B1(n9345), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6320));
   INVX1 U5795 (.Y(n9345), 
	.A(\ram[115][11] ));
   OAI22X1 U5796 (.Y(n2432), 
	.B1(n9346), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6322));
   INVX1 U5797 (.Y(n9346), 
	.A(\ram[115][10] ));
   OAI22X1 U5798 (.Y(n2431), 
	.B1(n9347), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6324));
   INVX1 U5799 (.Y(n9347), 
	.A(\ram[115][9] ));
   OAI22X1 U5800 (.Y(n2430), 
	.B1(n9348), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6326));
   INVX1 U5801 (.Y(n9348), 
	.A(\ram[115][8] ));
   OAI22X1 U5802 (.Y(n2429), 
	.B1(n9349), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6328));
   INVX1 U5803 (.Y(n9349), 
	.A(\ram[115][7] ));
   OAI22X1 U5804 (.Y(n2428), 
	.B1(n9350), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6330));
   INVX1 U5805 (.Y(n9350), 
	.A(\ram[115][6] ));
   OAI22X1 U5806 (.Y(n2427), 
	.B1(n9351), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6332));
   INVX1 U5807 (.Y(n9351), 
	.A(\ram[115][5] ));
   OAI22X1 U5808 (.Y(n2426), 
	.B1(n9352), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6334));
   INVX1 U5809 (.Y(n9352), 
	.A(\ram[115][4] ));
   OAI22X1 U5810 (.Y(n2425), 
	.B1(n9353), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6336));
   INVX1 U5811 (.Y(n9353), 
	.A(\ram[115][3] ));
   OAI22X1 U5812 (.Y(n2424), 
	.B1(n9354), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6338));
   INVX1 U5813 (.Y(n9354), 
	.A(\ram[115][2] ));
   OAI22X1 U5814 (.Y(n2423), 
	.B1(n9355), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6306));
   INVX1 U5815 (.Y(n9355), 
	.A(\ram[115][1] ));
   OAI22X1 U5816 (.Y(n2422), 
	.B1(n9356), 
	.B0(n9340), 
	.A1(n9339), 
	.A0(n6309));
   INVX1 U5817 (.Y(n9356), 
	.A(\ram[115][0] ));
   NOR2BX1 U5818 (.Y(n9340), 
	.B(n9339), 
	.AN(mem_write_en));
   NAND2X1 U5819 (.Y(n9339), 
	.B(n6457), 
	.A(n9140));
   OAI22X1 U5820 (.Y(n2421), 
	.B1(n9359), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6311));
   INVX1 U5821 (.Y(n9359), 
	.A(\ram[114][15] ));
   OAI22X1 U5822 (.Y(n2420), 
	.B1(n9360), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6314));
   INVX1 U5823 (.Y(n9360), 
	.A(\ram[114][14] ));
   OAI22X1 U5824 (.Y(n2419), 
	.B1(n9361), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6316));
   INVX1 U5825 (.Y(n9361), 
	.A(\ram[114][13] ));
   OAI22X1 U5826 (.Y(n2418), 
	.B1(n9362), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6318));
   INVX1 U5827 (.Y(n9362), 
	.A(\ram[114][12] ));
   OAI22X1 U5828 (.Y(n2417), 
	.B1(n9363), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6320));
   INVX1 U5829 (.Y(n9363), 
	.A(\ram[114][11] ));
   OAI22X1 U5830 (.Y(n2416), 
	.B1(n9364), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6322));
   INVX1 U5831 (.Y(n9364), 
	.A(\ram[114][10] ));
   OAI22X1 U5832 (.Y(n2415), 
	.B1(n9365), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6324));
   INVX1 U5833 (.Y(n9365), 
	.A(\ram[114][9] ));
   OAI22X1 U5834 (.Y(n2414), 
	.B1(n9366), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6326));
   INVX1 U5835 (.Y(n9366), 
	.A(\ram[114][8] ));
   OAI22X1 U5836 (.Y(n2413), 
	.B1(n9367), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6328));
   INVX1 U5837 (.Y(n9367), 
	.A(\ram[114][7] ));
   OAI22X1 U5838 (.Y(n2412), 
	.B1(n9368), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6330));
   INVX1 U5839 (.Y(n9368), 
	.A(\ram[114][6] ));
   OAI22X1 U5840 (.Y(n2411), 
	.B1(n9369), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6332));
   INVX1 U5841 (.Y(n9369), 
	.A(\ram[114][5] ));
   OAI22X1 U5842 (.Y(n2410), 
	.B1(n9370), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6334));
   INVX1 U5843 (.Y(n9370), 
	.A(\ram[114][4] ));
   OAI22X1 U5844 (.Y(n2409), 
	.B1(n9371), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6336));
   INVX1 U5845 (.Y(n9371), 
	.A(\ram[114][3] ));
   OAI22X1 U5846 (.Y(n2408), 
	.B1(n9372), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6338));
   INVX1 U5847 (.Y(n9372), 
	.A(\ram[114][2] ));
   OAI22X1 U5848 (.Y(n2407), 
	.B1(n9373), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6306));
   INVX1 U5849 (.Y(n9373), 
	.A(\ram[114][1] ));
   OAI22X1 U5850 (.Y(n2406), 
	.B1(n9374), 
	.B0(n9358), 
	.A1(n9357), 
	.A0(n6309));
   INVX1 U5851 (.Y(n9374), 
	.A(\ram[114][0] ));
   NOR2BX1 U5852 (.Y(n9358), 
	.B(n9357), 
	.AN(mem_write_en));
   NAND2X1 U5853 (.Y(n9357), 
	.B(n6476), 
	.A(n9140));
   OAI22X1 U5854 (.Y(n2405), 
	.B1(n9377), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6311));
   INVX1 U5855 (.Y(n9377), 
	.A(\ram[113][15] ));
   OAI22X1 U5856 (.Y(n2404), 
	.B1(n9378), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6314));
   INVX1 U5857 (.Y(n9378), 
	.A(\ram[113][14] ));
   OAI22X1 U5858 (.Y(n2403), 
	.B1(n9379), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6316));
   INVX1 U5859 (.Y(n9379), 
	.A(\ram[113][13] ));
   OAI22X1 U5860 (.Y(n2402), 
	.B1(n9380), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6318));
   INVX1 U5861 (.Y(n9380), 
	.A(\ram[113][12] ));
   OAI22X1 U5862 (.Y(n2401), 
	.B1(n9381), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6320));
   INVX1 U5863 (.Y(n9381), 
	.A(\ram[113][11] ));
   OAI22X1 U5864 (.Y(n2400), 
	.B1(n9382), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6322));
   INVX1 U5865 (.Y(n9382), 
	.A(\ram[113][10] ));
   OAI22X1 U5866 (.Y(n2399), 
	.B1(n9383), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6324));
   INVX1 U5867 (.Y(n9383), 
	.A(\ram[113][9] ));
   OAI22X1 U5868 (.Y(n2398), 
	.B1(n9384), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6326));
   INVX1 U5869 (.Y(n9384), 
	.A(\ram[113][8] ));
   OAI22X1 U5870 (.Y(n2397), 
	.B1(n9385), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6328));
   INVX1 U5871 (.Y(n9385), 
	.A(\ram[113][7] ));
   OAI22X1 U5872 (.Y(n2396), 
	.B1(n9386), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6330));
   INVX1 U5873 (.Y(n9386), 
	.A(\ram[113][6] ));
   OAI22X1 U5874 (.Y(n2395), 
	.B1(n9387), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6332));
   INVX1 U5875 (.Y(n9387), 
	.A(\ram[113][5] ));
   OAI22X1 U5876 (.Y(n2394), 
	.B1(n9388), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6334));
   INVX1 U5877 (.Y(n9388), 
	.A(\ram[113][4] ));
   OAI22X1 U5878 (.Y(n2393), 
	.B1(n9389), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6336));
   INVX1 U5879 (.Y(n9389), 
	.A(\ram[113][3] ));
   OAI22X1 U5880 (.Y(n2392), 
	.B1(n9390), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6338));
   INVX1 U5881 (.Y(n9390), 
	.A(\ram[113][2] ));
   OAI22X1 U5882 (.Y(n2391), 
	.B1(n9391), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6306));
   INVX1 U5883 (.Y(n9391), 
	.A(\ram[113][1] ));
   OAI22X1 U5884 (.Y(n2390), 
	.B1(n9392), 
	.B0(n9376), 
	.A1(n9375), 
	.A0(n6309));
   INVX1 U5885 (.Y(n9392), 
	.A(\ram[113][0] ));
   NOR2BX1 U5886 (.Y(n9376), 
	.B(n9375), 
	.AN(mem_write_en));
   NAND2X1 U5887 (.Y(n9375), 
	.B(n6495), 
	.A(n9140));
   OAI22X1 U5888 (.Y(n2389), 
	.B1(n9395), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6311));
   INVX1 U5889 (.Y(n9395), 
	.A(\ram[112][15] ));
   OAI22X1 U5890 (.Y(n2388), 
	.B1(n9396), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6314));
   INVX1 U5891 (.Y(n9396), 
	.A(\ram[112][14] ));
   OAI22X1 U5892 (.Y(n2387), 
	.B1(n9397), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6316));
   INVX1 U5893 (.Y(n9397), 
	.A(\ram[112][13] ));
   OAI22X1 U5894 (.Y(n2386), 
	.B1(n9398), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6318));
   INVX1 U5895 (.Y(n9398), 
	.A(\ram[112][12] ));
   OAI22X1 U5896 (.Y(n2385), 
	.B1(n9399), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6320));
   INVX1 U5897 (.Y(n9399), 
	.A(\ram[112][11] ));
   OAI22X1 U5898 (.Y(n2384), 
	.B1(n9400), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6322));
   INVX1 U5899 (.Y(n9400), 
	.A(\ram[112][10] ));
   OAI22X1 U5900 (.Y(n2383), 
	.B1(n9401), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6324));
   INVX1 U5901 (.Y(n9401), 
	.A(\ram[112][9] ));
   OAI22X1 U5902 (.Y(n2382), 
	.B1(n9402), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6326));
   INVX1 U5903 (.Y(n9402), 
	.A(\ram[112][8] ));
   OAI22X1 U5904 (.Y(n2381), 
	.B1(n9403), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6328));
   INVX1 U5905 (.Y(n9403), 
	.A(\ram[112][7] ));
   OAI22X1 U5906 (.Y(n2380), 
	.B1(n9404), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6330));
   INVX1 U5907 (.Y(n9404), 
	.A(\ram[112][6] ));
   OAI22X1 U5908 (.Y(n2379), 
	.B1(n9405), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6332));
   INVX1 U5909 (.Y(n9405), 
	.A(\ram[112][5] ));
   OAI22X1 U5910 (.Y(n2378), 
	.B1(n9406), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6334));
   INVX1 U5911 (.Y(n9406), 
	.A(\ram[112][4] ));
   OAI22X1 U5912 (.Y(n2377), 
	.B1(n9407), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6336));
   INVX1 U5913 (.Y(n9407), 
	.A(\ram[112][3] ));
   OAI22X1 U5914 (.Y(n2376), 
	.B1(n9408), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6338));
   INVX1 U5915 (.Y(n9408), 
	.A(\ram[112][2] ));
   OAI22X1 U5916 (.Y(n2375), 
	.B1(n9409), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6306));
   INVX1 U5917 (.Y(n9409), 
	.A(\ram[112][1] ));
   OAI22X1 U5918 (.Y(n2374), 
	.B1(n9410), 
	.B0(n9394), 
	.A1(n9393), 
	.A0(n6309));
   INVX1 U5919 (.Y(n9410), 
	.A(\ram[112][0] ));
   NOR2BX1 U5920 (.Y(n9394), 
	.B(n9393), 
	.AN(mem_write_en));
   NAND2X1 U5921 (.Y(n9393), 
	.B(n6514), 
	.A(n9140));
   OAI22X1 U5922 (.Y(n2373), 
	.B1(n9413), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6311));
   INVX1 U5923 (.Y(n9413), 
	.A(\ram[111][15] ));
   OAI22X1 U5924 (.Y(n2372), 
	.B1(n9414), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6314));
   INVX1 U5925 (.Y(n9414), 
	.A(\ram[111][14] ));
   OAI22X1 U5926 (.Y(n2371), 
	.B1(n9415), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6316));
   INVX1 U5927 (.Y(n9415), 
	.A(\ram[111][13] ));
   OAI22X1 U5928 (.Y(n2370), 
	.B1(n9416), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6318));
   INVX1 U5929 (.Y(n9416), 
	.A(\ram[111][12] ));
   OAI22X1 U5930 (.Y(n2369), 
	.B1(n9417), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6320));
   INVX1 U5931 (.Y(n9417), 
	.A(\ram[111][11] ));
   OAI22X1 U5932 (.Y(n2368), 
	.B1(n9418), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6322));
   INVX1 U5933 (.Y(n9418), 
	.A(\ram[111][10] ));
   OAI22X1 U5934 (.Y(n2367), 
	.B1(n9419), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6324));
   INVX1 U5935 (.Y(n9419), 
	.A(\ram[111][9] ));
   OAI22X1 U5936 (.Y(n2366), 
	.B1(n9420), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6326));
   INVX1 U5937 (.Y(n9420), 
	.A(\ram[111][8] ));
   OAI22X1 U5938 (.Y(n2365), 
	.B1(n9421), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6328));
   INVX1 U5939 (.Y(n9421), 
	.A(\ram[111][7] ));
   OAI22X1 U5940 (.Y(n2364), 
	.B1(n9422), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6330));
   INVX1 U5941 (.Y(n9422), 
	.A(\ram[111][6] ));
   OAI22X1 U5942 (.Y(n2363), 
	.B1(n9423), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6332));
   INVX1 U5943 (.Y(n9423), 
	.A(\ram[111][5] ));
   OAI22X1 U5944 (.Y(n2362), 
	.B1(n9424), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6334));
   INVX1 U5945 (.Y(n9424), 
	.A(\ram[111][4] ));
   OAI22X1 U5946 (.Y(n2361), 
	.B1(n9425), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6336));
   INVX1 U5947 (.Y(n9425), 
	.A(\ram[111][3] ));
   OAI22X1 U5948 (.Y(n2360), 
	.B1(n9426), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6338));
   INVX1 U5949 (.Y(n9426), 
	.A(\ram[111][2] ));
   OAI22X1 U5950 (.Y(n2359), 
	.B1(n9427), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6306));
   INVX1 U5951 (.Y(n9427), 
	.A(\ram[111][1] ));
   OAI22X1 U5952 (.Y(n2358), 
	.B1(n9428), 
	.B0(n9412), 
	.A1(n9411), 
	.A0(n6309));
   INVX1 U5953 (.Y(n9428), 
	.A(\ram[111][0] ));
   NOR2BX1 U5954 (.Y(n9412), 
	.B(n9411), 
	.AN(mem_write_en));
   NAND2X1 U5955 (.Y(n9411), 
	.B(n6533), 
	.A(n9429));
   OAI22X1 U5956 (.Y(n2357), 
	.B1(n9432), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6311));
   INVX1 U5957 (.Y(n9432), 
	.A(\ram[110][15] ));
   OAI22X1 U5958 (.Y(n2356), 
	.B1(n9433), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6314));
   INVX1 U5959 (.Y(n9433), 
	.A(\ram[110][14] ));
   OAI22X1 U5960 (.Y(n2355), 
	.B1(n9434), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6316));
   INVX1 U5961 (.Y(n9434), 
	.A(\ram[110][13] ));
   OAI22X1 U5962 (.Y(n2354), 
	.B1(n9435), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6318));
   INVX1 U5963 (.Y(n9435), 
	.A(\ram[110][12] ));
   OAI22X1 U5964 (.Y(n2353), 
	.B1(n9436), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6320));
   INVX1 U5965 (.Y(n9436), 
	.A(\ram[110][11] ));
   OAI22X1 U5966 (.Y(n2352), 
	.B1(n9437), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6322));
   INVX1 U5967 (.Y(n9437), 
	.A(\ram[110][10] ));
   OAI22X1 U5968 (.Y(n2351), 
	.B1(n9438), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6324));
   INVX1 U5969 (.Y(n9438), 
	.A(\ram[110][9] ));
   OAI22X1 U5970 (.Y(n2350), 
	.B1(n9439), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6326));
   INVX1 U5971 (.Y(n9439), 
	.A(\ram[110][8] ));
   OAI22X1 U5972 (.Y(n2349), 
	.B1(n9440), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6328));
   INVX1 U5973 (.Y(n9440), 
	.A(\ram[110][7] ));
   OAI22X1 U5974 (.Y(n2348), 
	.B1(n9441), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6330));
   INVX1 U5975 (.Y(n9441), 
	.A(\ram[110][6] ));
   OAI22X1 U5976 (.Y(n2347), 
	.B1(n9442), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6332));
   INVX1 U5977 (.Y(n9442), 
	.A(\ram[110][5] ));
   OAI22X1 U5978 (.Y(n2346), 
	.B1(n9443), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6334));
   INVX1 U5979 (.Y(n9443), 
	.A(\ram[110][4] ));
   OAI22X1 U5980 (.Y(n2345), 
	.B1(n9444), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6336));
   INVX1 U5981 (.Y(n9444), 
	.A(\ram[110][3] ));
   OAI22X1 U5982 (.Y(n2344), 
	.B1(n9445), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6338));
   INVX1 U5983 (.Y(n9445), 
	.A(\ram[110][2] ));
   OAI22X1 U5984 (.Y(n2343), 
	.B1(n9446), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6306));
   INVX1 U5985 (.Y(n9446), 
	.A(\ram[110][1] ));
   OAI22X1 U5986 (.Y(n2342), 
	.B1(n9447), 
	.B0(n9431), 
	.A1(n9430), 
	.A0(n6309));
   INVX1 U5987 (.Y(n9447), 
	.A(\ram[110][0] ));
   NOR2BX1 U5988 (.Y(n9431), 
	.B(n9430), 
	.AN(mem_write_en));
   NAND2X1 U5989 (.Y(n9430), 
	.B(n6553), 
	.A(n9429));
   OAI22X1 U5990 (.Y(n2341), 
	.B1(n9450), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6311));
   INVX1 U5991 (.Y(n9450), 
	.A(\ram[109][15] ));
   OAI22X1 U5992 (.Y(n2340), 
	.B1(n9451), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6314));
   INVX1 U5993 (.Y(n9451), 
	.A(\ram[109][14] ));
   OAI22X1 U5994 (.Y(n2339), 
	.B1(n9452), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6316));
   INVX1 U5995 (.Y(n9452), 
	.A(\ram[109][13] ));
   OAI22X1 U5996 (.Y(n2338), 
	.B1(n9453), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6318));
   INVX1 U5997 (.Y(n9453), 
	.A(\ram[109][12] ));
   OAI22X1 U5998 (.Y(n2337), 
	.B1(n9454), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6320));
   INVX1 U5999 (.Y(n9454), 
	.A(\ram[109][11] ));
   OAI22X1 U6000 (.Y(n2336), 
	.B1(n9455), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6322));
   INVX1 U6001 (.Y(n9455), 
	.A(\ram[109][10] ));
   OAI22X1 U6002 (.Y(n2335), 
	.B1(n9456), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6324));
   INVX1 U6003 (.Y(n9456), 
	.A(\ram[109][9] ));
   OAI22X1 U6004 (.Y(n2334), 
	.B1(n9457), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6326));
   INVX1 U6005 (.Y(n9457), 
	.A(\ram[109][8] ));
   OAI22X1 U6006 (.Y(n2333), 
	.B1(n9458), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6328));
   INVX1 U6007 (.Y(n9458), 
	.A(\ram[109][7] ));
   OAI22X1 U6008 (.Y(n2332), 
	.B1(n9459), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6330));
   INVX1 U6009 (.Y(n9459), 
	.A(\ram[109][6] ));
   OAI22X1 U6010 (.Y(n2331), 
	.B1(n9460), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6332));
   INVX1 U6011 (.Y(n9460), 
	.A(\ram[109][5] ));
   OAI22X1 U6012 (.Y(n2330), 
	.B1(n9461), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6334));
   INVX1 U6013 (.Y(n9461), 
	.A(\ram[109][4] ));
   OAI22X1 U6014 (.Y(n2329), 
	.B1(n9462), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6336));
   INVX1 U6015 (.Y(n9462), 
	.A(\ram[109][3] ));
   OAI22X1 U6016 (.Y(n2328), 
	.B1(n9463), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6338));
   INVX1 U6017 (.Y(n9463), 
	.A(\ram[109][2] ));
   OAI22X1 U6018 (.Y(n2327), 
	.B1(n9464), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6306));
   INVX1 U6019 (.Y(n9464), 
	.A(\ram[109][1] ));
   OAI22X1 U6020 (.Y(n2326), 
	.B1(n9465), 
	.B0(n9449), 
	.A1(n9448), 
	.A0(n6309));
   INVX1 U6021 (.Y(n9465), 
	.A(\ram[109][0] ));
   NOR2BX1 U6022 (.Y(n9449), 
	.B(n9448), 
	.AN(mem_write_en));
   NAND2X1 U6023 (.Y(n9448), 
	.B(n6572), 
	.A(n9429));
   OAI22X1 U6024 (.Y(n2325), 
	.B1(n9468), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6311));
   INVX1 U6025 (.Y(n9468), 
	.A(\ram[108][15] ));
   OAI22X1 U6026 (.Y(n2324), 
	.B1(n9469), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6314));
   INVX1 U6027 (.Y(n9469), 
	.A(\ram[108][14] ));
   OAI22X1 U6028 (.Y(n2323), 
	.B1(n9470), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6316));
   INVX1 U6029 (.Y(n9470), 
	.A(\ram[108][13] ));
   OAI22X1 U6030 (.Y(n2322), 
	.B1(n9471), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6318));
   INVX1 U6031 (.Y(n9471), 
	.A(\ram[108][12] ));
   OAI22X1 U6032 (.Y(n2321), 
	.B1(n9472), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6320));
   INVX1 U6033 (.Y(n9472), 
	.A(\ram[108][11] ));
   OAI22X1 U6034 (.Y(n2320), 
	.B1(n9473), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6322));
   INVX1 U6035 (.Y(n9473), 
	.A(\ram[108][10] ));
   OAI22X1 U6036 (.Y(n2319), 
	.B1(n9474), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6324));
   INVX1 U6037 (.Y(n9474), 
	.A(\ram[108][9] ));
   OAI22X1 U6038 (.Y(n2318), 
	.B1(n9475), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6326));
   INVX1 U6039 (.Y(n9475), 
	.A(\ram[108][8] ));
   OAI22X1 U6040 (.Y(n2317), 
	.B1(n9476), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6328));
   INVX1 U6041 (.Y(n9476), 
	.A(\ram[108][7] ));
   OAI22X1 U6042 (.Y(n2316), 
	.B1(n9477), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6330));
   INVX1 U6043 (.Y(n9477), 
	.A(\ram[108][6] ));
   OAI22X1 U6044 (.Y(n2315), 
	.B1(n9478), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6332));
   INVX1 U6045 (.Y(n9478), 
	.A(\ram[108][5] ));
   OAI22X1 U6046 (.Y(n2314), 
	.B1(n9479), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6334));
   INVX1 U6047 (.Y(n9479), 
	.A(\ram[108][4] ));
   OAI22X1 U6048 (.Y(n2313), 
	.B1(n9480), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6336));
   INVX1 U6049 (.Y(n9480), 
	.A(\ram[108][3] ));
   OAI22X1 U6050 (.Y(n2312), 
	.B1(n9481), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6338));
   INVX1 U6051 (.Y(n9481), 
	.A(\ram[108][2] ));
   OAI22X1 U6052 (.Y(n2311), 
	.B1(n9482), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6306));
   INVX1 U6053 (.Y(n9482), 
	.A(\ram[108][1] ));
   OAI22X1 U6054 (.Y(n2310), 
	.B1(n9483), 
	.B0(n9467), 
	.A1(n9466), 
	.A0(n6309));
   INVX1 U6055 (.Y(n9483), 
	.A(\ram[108][0] ));
   NOR2BX1 U6056 (.Y(n9467), 
	.B(n9466), 
	.AN(mem_write_en));
   NAND2X1 U6057 (.Y(n9466), 
	.B(n6591), 
	.A(n9429));
   OAI22X1 U6058 (.Y(n2309), 
	.B1(n9486), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6311));
   INVX1 U6059 (.Y(n9486), 
	.A(\ram[107][15] ));
   OAI22X1 U6060 (.Y(n2308), 
	.B1(n9487), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6314));
   INVX1 U6061 (.Y(n9487), 
	.A(\ram[107][14] ));
   OAI22X1 U6062 (.Y(n2307), 
	.B1(n9488), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6316));
   INVX1 U6063 (.Y(n9488), 
	.A(\ram[107][13] ));
   OAI22X1 U6064 (.Y(n2306), 
	.B1(n9489), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6318));
   INVX1 U6065 (.Y(n9489), 
	.A(\ram[107][12] ));
   OAI22X1 U6066 (.Y(n2305), 
	.B1(n9490), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6320));
   INVX1 U6067 (.Y(n9490), 
	.A(\ram[107][11] ));
   OAI22X1 U6068 (.Y(n2304), 
	.B1(n9491), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6322));
   INVX1 U6069 (.Y(n9491), 
	.A(\ram[107][10] ));
   OAI22X1 U6070 (.Y(n2303), 
	.B1(n9492), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6324));
   INVX1 U6071 (.Y(n9492), 
	.A(\ram[107][9] ));
   OAI22X1 U6072 (.Y(n2302), 
	.B1(n9493), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6326));
   INVX1 U6073 (.Y(n9493), 
	.A(\ram[107][8] ));
   OAI22X1 U6074 (.Y(n2301), 
	.B1(n9494), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6328));
   INVX1 U6075 (.Y(n9494), 
	.A(\ram[107][7] ));
   OAI22X1 U6076 (.Y(n2300), 
	.B1(n9495), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6330));
   INVX1 U6077 (.Y(n9495), 
	.A(\ram[107][6] ));
   OAI22X1 U6078 (.Y(n2299), 
	.B1(n9496), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6332));
   INVX1 U6079 (.Y(n9496), 
	.A(\ram[107][5] ));
   OAI22X1 U6080 (.Y(n2298), 
	.B1(n9497), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6334));
   INVX1 U6081 (.Y(n9497), 
	.A(\ram[107][4] ));
   OAI22X1 U6082 (.Y(n2297), 
	.B1(n9498), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6336));
   INVX1 U6083 (.Y(n9498), 
	.A(\ram[107][3] ));
   OAI22X1 U6084 (.Y(n2296), 
	.B1(n9499), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6338));
   INVX1 U6085 (.Y(n9499), 
	.A(\ram[107][2] ));
   OAI22X1 U6086 (.Y(n2295), 
	.B1(n9500), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6306));
   INVX1 U6087 (.Y(n9500), 
	.A(\ram[107][1] ));
   OAI22X1 U6088 (.Y(n2294), 
	.B1(n9501), 
	.B0(n9485), 
	.A1(n9484), 
	.A0(n6309));
   INVX1 U6089 (.Y(n9501), 
	.A(\ram[107][0] ));
   NOR2BX1 U6090 (.Y(n9485), 
	.B(n9484), 
	.AN(mem_write_en));
   NAND2X1 U6091 (.Y(n9484), 
	.B(n6610), 
	.A(n9429));
   OAI22X1 U6092 (.Y(n2293), 
	.B1(n9504), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6311));
   INVX1 U6093 (.Y(n9504), 
	.A(\ram[106][15] ));
   OAI22X1 U6094 (.Y(n2292), 
	.B1(n9505), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6314));
   INVX1 U6095 (.Y(n9505), 
	.A(\ram[106][14] ));
   OAI22X1 U6096 (.Y(n2291), 
	.B1(n9506), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6316));
   INVX1 U6097 (.Y(n9506), 
	.A(\ram[106][13] ));
   OAI22X1 U6098 (.Y(n2290), 
	.B1(n9507), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6318));
   INVX1 U6099 (.Y(n9507), 
	.A(\ram[106][12] ));
   OAI22X1 U6100 (.Y(n2289), 
	.B1(n9508), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6320));
   INVX1 U6101 (.Y(n9508), 
	.A(\ram[106][11] ));
   OAI22X1 U6102 (.Y(n2288), 
	.B1(n9509), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6322));
   INVX1 U6103 (.Y(n9509), 
	.A(\ram[106][10] ));
   OAI22X1 U6104 (.Y(n2287), 
	.B1(n9510), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6324));
   INVX1 U6105 (.Y(n9510), 
	.A(\ram[106][9] ));
   OAI22X1 U6106 (.Y(n2286), 
	.B1(n9511), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6326));
   INVX1 U6107 (.Y(n9511), 
	.A(\ram[106][8] ));
   OAI22X1 U6108 (.Y(n2285), 
	.B1(n9512), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6328));
   INVX1 U6109 (.Y(n9512), 
	.A(\ram[106][7] ));
   OAI22X1 U6110 (.Y(n2284), 
	.B1(n9513), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6330));
   INVX1 U6111 (.Y(n9513), 
	.A(\ram[106][6] ));
   OAI22X1 U6112 (.Y(n2283), 
	.B1(n9514), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6332));
   INVX1 U6113 (.Y(n9514), 
	.A(\ram[106][5] ));
   OAI22X1 U6114 (.Y(n2282), 
	.B1(n9515), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6334));
   INVX1 U6115 (.Y(n9515), 
	.A(\ram[106][4] ));
   OAI22X1 U6116 (.Y(n2281), 
	.B1(n9516), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6336));
   INVX1 U6117 (.Y(n9516), 
	.A(\ram[106][3] ));
   OAI22X1 U6118 (.Y(n2280), 
	.B1(n9517), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6338));
   INVX1 U6119 (.Y(n9517), 
	.A(\ram[106][2] ));
   OAI22X1 U6120 (.Y(n2279), 
	.B1(n9518), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6306));
   INVX1 U6121 (.Y(n9518), 
	.A(\ram[106][1] ));
   OAI22X1 U6122 (.Y(n2278), 
	.B1(n9519), 
	.B0(n9503), 
	.A1(n9502), 
	.A0(n6309));
   INVX1 U6123 (.Y(n9519), 
	.A(\ram[106][0] ));
   NOR2BX1 U6124 (.Y(n9503), 
	.B(n9502), 
	.AN(mem_write_en));
   NAND2X1 U6125 (.Y(n9502), 
	.B(n6629), 
	.A(n9429));
   OAI22X1 U6126 (.Y(n2277), 
	.B1(n9522), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6311));
   INVX1 U6127 (.Y(n9522), 
	.A(\ram[105][15] ));
   OAI22X1 U6128 (.Y(n2276), 
	.B1(n9523), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6314));
   INVX1 U6129 (.Y(n9523), 
	.A(\ram[105][14] ));
   OAI22X1 U6130 (.Y(n2275), 
	.B1(n9524), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6316));
   INVX1 U6131 (.Y(n9524), 
	.A(\ram[105][13] ));
   OAI22X1 U6132 (.Y(n2274), 
	.B1(n9525), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6318));
   INVX1 U6133 (.Y(n9525), 
	.A(\ram[105][12] ));
   OAI22X1 U6134 (.Y(n2273), 
	.B1(n9526), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6320));
   INVX1 U6135 (.Y(n9526), 
	.A(\ram[105][11] ));
   OAI22X1 U6136 (.Y(n2272), 
	.B1(n9527), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6322));
   INVX1 U6137 (.Y(n9527), 
	.A(\ram[105][10] ));
   OAI22X1 U6138 (.Y(n2271), 
	.B1(n9528), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6324));
   INVX1 U6139 (.Y(n9528), 
	.A(\ram[105][9] ));
   OAI22X1 U6140 (.Y(n2270), 
	.B1(n9529), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6326));
   INVX1 U6141 (.Y(n9529), 
	.A(\ram[105][8] ));
   OAI22X1 U6142 (.Y(n2269), 
	.B1(n9530), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6328));
   INVX1 U6143 (.Y(n9530), 
	.A(\ram[105][7] ));
   OAI22X1 U6144 (.Y(n2268), 
	.B1(n9531), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6330));
   INVX1 U6145 (.Y(n9531), 
	.A(\ram[105][6] ));
   OAI22X1 U6146 (.Y(n2267), 
	.B1(n9532), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6332));
   INVX1 U6147 (.Y(n9532), 
	.A(\ram[105][5] ));
   OAI22X1 U6148 (.Y(n2266), 
	.B1(n9533), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6334));
   INVX1 U6149 (.Y(n9533), 
	.A(\ram[105][4] ));
   OAI22X1 U6150 (.Y(n2265), 
	.B1(n9534), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6336));
   INVX1 U6151 (.Y(n9534), 
	.A(\ram[105][3] ));
   OAI22X1 U6152 (.Y(n2264), 
	.B1(n9535), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6338));
   INVX1 U6153 (.Y(n9535), 
	.A(\ram[105][2] ));
   OAI22X1 U6154 (.Y(n2263), 
	.B1(n9536), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6306));
   INVX1 U6155 (.Y(n9536), 
	.A(\ram[105][1] ));
   OAI22X1 U6156 (.Y(n2262), 
	.B1(n9537), 
	.B0(n9521), 
	.A1(n9520), 
	.A0(n6309));
   INVX1 U6157 (.Y(n9537), 
	.A(\ram[105][0] ));
   NOR2BX1 U6158 (.Y(n9521), 
	.B(n9520), 
	.AN(mem_write_en));
   NAND2X1 U6159 (.Y(n9520), 
	.B(n6342), 
	.A(n9429));
   OAI22X1 U6160 (.Y(n2261), 
	.B1(n9540), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6311));
   INVX1 U6161 (.Y(n9540), 
	.A(\ram[104][15] ));
   OAI22X1 U6162 (.Y(n2260), 
	.B1(n9541), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6314));
   INVX1 U6163 (.Y(n9541), 
	.A(\ram[104][14] ));
   OAI22X1 U6164 (.Y(n2259), 
	.B1(n9542), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6316));
   INVX1 U6165 (.Y(n9542), 
	.A(\ram[104][13] ));
   OAI22X1 U6166 (.Y(n2258), 
	.B1(n9543), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6318));
   INVX1 U6167 (.Y(n9543), 
	.A(\ram[104][12] ));
   OAI22X1 U6168 (.Y(n2257), 
	.B1(n9544), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6320));
   INVX1 U6169 (.Y(n9544), 
	.A(\ram[104][11] ));
   OAI22X1 U6170 (.Y(n2256), 
	.B1(n9545), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6322));
   INVX1 U6171 (.Y(n9545), 
	.A(\ram[104][10] ));
   OAI22X1 U6172 (.Y(n2255), 
	.B1(n9546), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6324));
   INVX1 U6173 (.Y(n9546), 
	.A(\ram[104][9] ));
   OAI22X1 U6174 (.Y(n2254), 
	.B1(n9547), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6326));
   INVX1 U6175 (.Y(n9547), 
	.A(\ram[104][8] ));
   OAI22X1 U6176 (.Y(n2253), 
	.B1(n9548), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6328));
   INVX1 U6177 (.Y(n9548), 
	.A(\ram[104][7] ));
   OAI22X1 U6178 (.Y(n2252), 
	.B1(n9549), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6330));
   INVX1 U6179 (.Y(n9549), 
	.A(\ram[104][6] ));
   OAI22X1 U6180 (.Y(n2251), 
	.B1(n9550), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6332));
   INVX1 U6181 (.Y(n9550), 
	.A(\ram[104][5] ));
   OAI22X1 U6182 (.Y(n2250), 
	.B1(n9551), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6334));
   INVX1 U6183 (.Y(n9551), 
	.A(\ram[104][4] ));
   OAI22X1 U6184 (.Y(n2249), 
	.B1(n9552), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6336));
   INVX1 U6185 (.Y(n9552), 
	.A(\ram[104][3] ));
   OAI22X1 U6186 (.Y(n2248), 
	.B1(n9553), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6338));
   INVX1 U6187 (.Y(n9553), 
	.A(\ram[104][2] ));
   OAI22X1 U6188 (.Y(n2247), 
	.B1(n9554), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6306));
   INVX1 U6189 (.Y(n9554), 
	.A(\ram[104][1] ));
   OAI22X1 U6190 (.Y(n2246), 
	.B1(n9555), 
	.B0(n9539), 
	.A1(n9538), 
	.A0(n6309));
   INVX1 U6191 (.Y(n9555), 
	.A(\ram[104][0] ));
   NOR2BX1 U6192 (.Y(n9539), 
	.B(n9538), 
	.AN(mem_write_en));
   NAND2X1 U6193 (.Y(n9538), 
	.B(n6362), 
	.A(n9429));
   OAI22X1 U6194 (.Y(n2245), 
	.B1(n9558), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6311));
   INVX1 U6195 (.Y(n9558), 
	.A(\ram[103][15] ));
   OAI22X1 U6196 (.Y(n2244), 
	.B1(n9559), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6314));
   INVX1 U6197 (.Y(n9559), 
	.A(\ram[103][14] ));
   OAI22X1 U6198 (.Y(n2243), 
	.B1(n9560), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6316));
   INVX1 U6199 (.Y(n9560), 
	.A(\ram[103][13] ));
   OAI22X1 U6200 (.Y(n2242), 
	.B1(n9561), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6318));
   INVX1 U6201 (.Y(n9561), 
	.A(\ram[103][12] ));
   OAI22X1 U6202 (.Y(n2241), 
	.B1(n9562), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6320));
   INVX1 U6203 (.Y(n9562), 
	.A(\ram[103][11] ));
   OAI22X1 U6204 (.Y(n2240), 
	.B1(n9563), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6322));
   INVX1 U6205 (.Y(n9563), 
	.A(\ram[103][10] ));
   OAI22X1 U6206 (.Y(n2239), 
	.B1(n9564), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6324));
   INVX1 U6207 (.Y(n9564), 
	.A(\ram[103][9] ));
   OAI22X1 U6208 (.Y(n2238), 
	.B1(n9565), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6326));
   INVX1 U6209 (.Y(n9565), 
	.A(\ram[103][8] ));
   OAI22X1 U6210 (.Y(n2237), 
	.B1(n9566), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6328));
   INVX1 U6211 (.Y(n9566), 
	.A(\ram[103][7] ));
   OAI22X1 U6212 (.Y(n2236), 
	.B1(n9567), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6330));
   INVX1 U6213 (.Y(n9567), 
	.A(\ram[103][6] ));
   OAI22X1 U6214 (.Y(n2235), 
	.B1(n9568), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6332));
   INVX1 U6215 (.Y(n9568), 
	.A(\ram[103][5] ));
   OAI22X1 U6216 (.Y(n2234), 
	.B1(n9569), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6334));
   INVX1 U6217 (.Y(n9569), 
	.A(\ram[103][4] ));
   OAI22X1 U6218 (.Y(n2233), 
	.B1(n9570), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6336));
   INVX1 U6219 (.Y(n9570), 
	.A(\ram[103][3] ));
   OAI22X1 U6220 (.Y(n2232), 
	.B1(n9571), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6338));
   INVX1 U6221 (.Y(n9571), 
	.A(\ram[103][2] ));
   OAI22X1 U6222 (.Y(n2231), 
	.B1(n9572), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6306));
   INVX1 U6223 (.Y(n9572), 
	.A(\ram[103][1] ));
   OAI22X1 U6224 (.Y(n2230), 
	.B1(n9573), 
	.B0(n9557), 
	.A1(n9556), 
	.A0(n6309));
   INVX1 U6225 (.Y(n9573), 
	.A(\ram[103][0] ));
   NOR2BX1 U6226 (.Y(n9557), 
	.B(n9556), 
	.AN(mem_write_en));
   NAND2X1 U6227 (.Y(n9556), 
	.B(n6381), 
	.A(n9429));
   OAI22X1 U6228 (.Y(n2229), 
	.B1(n9576), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6311));
   INVX1 U6229 (.Y(n9576), 
	.A(\ram[102][15] ));
   OAI22X1 U6230 (.Y(n2228), 
	.B1(n9577), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6314));
   INVX1 U6231 (.Y(n9577), 
	.A(\ram[102][14] ));
   OAI22X1 U6232 (.Y(n2227), 
	.B1(n9578), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6316));
   INVX1 U6233 (.Y(n9578), 
	.A(\ram[102][13] ));
   OAI22X1 U6234 (.Y(n2226), 
	.B1(n9579), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6318));
   INVX1 U6235 (.Y(n9579), 
	.A(\ram[102][12] ));
   OAI22X1 U6236 (.Y(n2225), 
	.B1(n9580), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6320));
   INVX1 U6237 (.Y(n9580), 
	.A(\ram[102][11] ));
   OAI22X1 U6238 (.Y(n2224), 
	.B1(n9581), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6322));
   INVX1 U6239 (.Y(n9581), 
	.A(\ram[102][10] ));
   OAI22X1 U6240 (.Y(n2223), 
	.B1(n9582), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6324));
   INVX1 U6241 (.Y(n9582), 
	.A(\ram[102][9] ));
   OAI22X1 U6242 (.Y(n2222), 
	.B1(n9583), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6326));
   INVX1 U6243 (.Y(n9583), 
	.A(\ram[102][8] ));
   OAI22X1 U6244 (.Y(n2221), 
	.B1(n9584), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6328));
   INVX1 U6245 (.Y(n9584), 
	.A(\ram[102][7] ));
   OAI22X1 U6246 (.Y(n2220), 
	.B1(n9585), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6330));
   INVX1 U6247 (.Y(n9585), 
	.A(\ram[102][6] ));
   OAI22X1 U6248 (.Y(n2219), 
	.B1(n9586), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6332));
   INVX1 U6249 (.Y(n9586), 
	.A(\ram[102][5] ));
   OAI22X1 U6250 (.Y(n2218), 
	.B1(n9587), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6334));
   INVX1 U6251 (.Y(n9587), 
	.A(\ram[102][4] ));
   OAI22X1 U6252 (.Y(n2217), 
	.B1(n9588), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6336));
   INVX1 U6253 (.Y(n9588), 
	.A(\ram[102][3] ));
   OAI22X1 U6254 (.Y(n2216), 
	.B1(n9589), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6338));
   INVX1 U6255 (.Y(n9589), 
	.A(\ram[102][2] ));
   OAI22X1 U6256 (.Y(n2215), 
	.B1(n9590), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6306));
   INVX1 U6257 (.Y(n9590), 
	.A(\ram[102][1] ));
   OAI22X1 U6258 (.Y(n2214), 
	.B1(n9591), 
	.B0(n9575), 
	.A1(n9574), 
	.A0(n6309));
   INVX1 U6259 (.Y(n9591), 
	.A(\ram[102][0] ));
   NOR2BX1 U6260 (.Y(n9575), 
	.B(n9574), 
	.AN(mem_write_en));
   NAND2X1 U6261 (.Y(n9574), 
	.B(n6400), 
	.A(n9429));
   OAI22X1 U6262 (.Y(n2213), 
	.B1(n9594), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6311));
   INVX1 U6263 (.Y(n9594), 
	.A(\ram[101][15] ));
   OAI22X1 U6264 (.Y(n2212), 
	.B1(n9595), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6314));
   INVX1 U6265 (.Y(n9595), 
	.A(\ram[101][14] ));
   OAI22X1 U6266 (.Y(n2211), 
	.B1(n9596), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6316));
   INVX1 U6267 (.Y(n9596), 
	.A(\ram[101][13] ));
   OAI22X1 U6268 (.Y(n2210), 
	.B1(n9597), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6318));
   INVX1 U6269 (.Y(n9597), 
	.A(\ram[101][12] ));
   OAI22X1 U6270 (.Y(n2209), 
	.B1(n9598), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6320));
   INVX1 U6271 (.Y(n9598), 
	.A(\ram[101][11] ));
   OAI22X1 U6272 (.Y(n2208), 
	.B1(n9599), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6322));
   INVX1 U6273 (.Y(n9599), 
	.A(\ram[101][10] ));
   OAI22X1 U6274 (.Y(n2207), 
	.B1(n9600), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6324));
   INVX1 U6275 (.Y(n9600), 
	.A(\ram[101][9] ));
   OAI22X1 U6276 (.Y(n2206), 
	.B1(n9601), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6326));
   INVX1 U6277 (.Y(n9601), 
	.A(\ram[101][8] ));
   OAI22X1 U6278 (.Y(n2205), 
	.B1(n9602), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6328));
   INVX1 U6279 (.Y(n9602), 
	.A(\ram[101][7] ));
   OAI22X1 U6280 (.Y(n2204), 
	.B1(n9603), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6330));
   INVX1 U6281 (.Y(n9603), 
	.A(\ram[101][6] ));
   OAI22X1 U6282 (.Y(n2203), 
	.B1(n9604), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6332));
   INVX1 U6283 (.Y(n9604), 
	.A(\ram[101][5] ));
   OAI22X1 U6284 (.Y(n2202), 
	.B1(n9605), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6334));
   INVX1 U6285 (.Y(n9605), 
	.A(\ram[101][4] ));
   OAI22X1 U6286 (.Y(n2201), 
	.B1(n9606), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6336));
   INVX1 U6287 (.Y(n9606), 
	.A(\ram[101][3] ));
   OAI22X1 U6288 (.Y(n2200), 
	.B1(n9607), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6338));
   INVX1 U6289 (.Y(n9607), 
	.A(\ram[101][2] ));
   OAI22X1 U6290 (.Y(n2199), 
	.B1(n9608), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6306));
   INVX1 U6291 (.Y(n9608), 
	.A(\ram[101][1] ));
   OAI22X1 U6292 (.Y(n2198), 
	.B1(n9609), 
	.B0(n9593), 
	.A1(n9592), 
	.A0(n6309));
   INVX1 U6293 (.Y(n9609), 
	.A(\ram[101][0] ));
   NOR2BX1 U6294 (.Y(n9593), 
	.B(n9592), 
	.AN(mem_write_en));
   NAND2X1 U6295 (.Y(n9592), 
	.B(n6419), 
	.A(n9429));
   OAI22X1 U6296 (.Y(n2197), 
	.B1(n9612), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6311));
   INVX1 U6297 (.Y(n9612), 
	.A(\ram[100][15] ));
   OAI22X1 U6298 (.Y(n2196), 
	.B1(n9613), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6314));
   INVX1 U6299 (.Y(n9613), 
	.A(\ram[100][14] ));
   OAI22X1 U6300 (.Y(n2195), 
	.B1(n9614), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6316));
   INVX1 U6301 (.Y(n9614), 
	.A(\ram[100][13] ));
   OAI22X1 U6302 (.Y(n2194), 
	.B1(n9615), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6318));
   INVX1 U6303 (.Y(n9615), 
	.A(\ram[100][12] ));
   OAI22X1 U6304 (.Y(n2193), 
	.B1(n9616), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6320));
   INVX1 U6305 (.Y(n9616), 
	.A(\ram[100][11] ));
   OAI22X1 U6306 (.Y(n2192), 
	.B1(n9617), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6322));
   INVX1 U6307 (.Y(n9617), 
	.A(\ram[100][10] ));
   OAI22X1 U6308 (.Y(n2191), 
	.B1(n9618), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6324));
   INVX1 U6309 (.Y(n9618), 
	.A(\ram[100][9] ));
   OAI22X1 U6310 (.Y(n2190), 
	.B1(n9619), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6326));
   INVX1 U6311 (.Y(n9619), 
	.A(\ram[100][8] ));
   OAI22X1 U6312 (.Y(n2189), 
	.B1(n9620), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6328));
   INVX1 U6313 (.Y(n9620), 
	.A(\ram[100][7] ));
   OAI22X1 U6314 (.Y(n2188), 
	.B1(n9621), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6330));
   INVX1 U6315 (.Y(n9621), 
	.A(\ram[100][6] ));
   OAI22X1 U6316 (.Y(n2187), 
	.B1(n9622), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6332));
   INVX1 U6317 (.Y(n9622), 
	.A(\ram[100][5] ));
   OAI22X1 U6318 (.Y(n2186), 
	.B1(n9623), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6334));
   INVX1 U6319 (.Y(n9623), 
	.A(\ram[100][4] ));
   OAI22X1 U6320 (.Y(n2185), 
	.B1(n9624), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6336));
   INVX1 U6321 (.Y(n9624), 
	.A(\ram[100][3] ));
   OAI22X1 U6322 (.Y(n2184), 
	.B1(n9625), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6338));
   INVX1 U6323 (.Y(n9625), 
	.A(\ram[100][2] ));
   OAI22X1 U6324 (.Y(n2183), 
	.B1(n9626), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6306));
   INVX1 U6325 (.Y(n9626), 
	.A(\ram[100][1] ));
   OAI22X1 U6326 (.Y(n2182), 
	.B1(n9627), 
	.B0(n9611), 
	.A1(n9610), 
	.A0(n6309));
   INVX1 U6327 (.Y(n9627), 
	.A(\ram[100][0] ));
   NOR2BX1 U6328 (.Y(n9611), 
	.B(n9610), 
	.AN(mem_write_en));
   NAND2X1 U6329 (.Y(n9610), 
	.B(n6438), 
	.A(n9429));
   OAI22X1 U6330 (.Y(n2181), 
	.B1(n9630), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6311));
   INVX1 U6331 (.Y(n9630), 
	.A(\ram[99][15] ));
   OAI22X1 U6332 (.Y(n2180), 
	.B1(n9631), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6314));
   INVX1 U6333 (.Y(n9631), 
	.A(\ram[99][14] ));
   OAI22X1 U6334 (.Y(n2179), 
	.B1(n9632), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6316));
   INVX1 U6335 (.Y(n9632), 
	.A(\ram[99][13] ));
   OAI22X1 U6336 (.Y(n2178), 
	.B1(n9633), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6318));
   INVX1 U6337 (.Y(n9633), 
	.A(\ram[99][12] ));
   OAI22X1 U6338 (.Y(n2177), 
	.B1(n9634), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6320));
   INVX1 U6339 (.Y(n9634), 
	.A(\ram[99][11] ));
   OAI22X1 U6340 (.Y(n2176), 
	.B1(n9635), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6322));
   INVX1 U6341 (.Y(n9635), 
	.A(\ram[99][10] ));
   OAI22X1 U6342 (.Y(n2175), 
	.B1(n9636), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6324));
   INVX1 U6343 (.Y(n9636), 
	.A(\ram[99][9] ));
   OAI22X1 U6344 (.Y(n2174), 
	.B1(n9637), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6326));
   INVX1 U6345 (.Y(n9637), 
	.A(\ram[99][8] ));
   OAI22X1 U6346 (.Y(n2173), 
	.B1(n9638), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6328));
   INVX1 U6347 (.Y(n9638), 
	.A(\ram[99][7] ));
   OAI22X1 U6348 (.Y(n2172), 
	.B1(n9639), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6330));
   INVX1 U6349 (.Y(n9639), 
	.A(\ram[99][6] ));
   OAI22X1 U6350 (.Y(n2171), 
	.B1(n9640), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6332));
   INVX1 U6351 (.Y(n9640), 
	.A(\ram[99][5] ));
   OAI22X1 U6352 (.Y(n2170), 
	.B1(n9641), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6334));
   INVX1 U6353 (.Y(n9641), 
	.A(\ram[99][4] ));
   OAI22X1 U6354 (.Y(n2169), 
	.B1(n9642), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6336));
   INVX1 U6355 (.Y(n9642), 
	.A(\ram[99][3] ));
   OAI22X1 U6356 (.Y(n2168), 
	.B1(n9643), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6338));
   INVX1 U6357 (.Y(n9643), 
	.A(\ram[99][2] ));
   OAI22X1 U6358 (.Y(n2167), 
	.B1(n9644), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6306));
   INVX1 U6359 (.Y(n9644), 
	.A(\ram[99][1] ));
   OAI22X1 U6360 (.Y(n2166), 
	.B1(n9645), 
	.B0(n9629), 
	.A1(n9628), 
	.A0(n6309));
   INVX1 U6361 (.Y(n9645), 
	.A(\ram[99][0] ));
   NOR2BX1 U6362 (.Y(n9629), 
	.B(n9628), 
	.AN(mem_write_en));
   NAND2X1 U6363 (.Y(n9628), 
	.B(n6457), 
	.A(n9429));
   OAI22X1 U6364 (.Y(n2165), 
	.B1(n9648), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6311));
   INVX1 U6365 (.Y(n9648), 
	.A(\ram[98][15] ));
   OAI22X1 U6366 (.Y(n2164), 
	.B1(n9649), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6314));
   INVX1 U6367 (.Y(n9649), 
	.A(\ram[98][14] ));
   OAI22X1 U6368 (.Y(n2163), 
	.B1(n9650), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6316));
   INVX1 U6369 (.Y(n9650), 
	.A(\ram[98][13] ));
   OAI22X1 U6370 (.Y(n2162), 
	.B1(n9651), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6318));
   INVX1 U6371 (.Y(n9651), 
	.A(\ram[98][12] ));
   OAI22X1 U6372 (.Y(n2161), 
	.B1(n9652), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6320));
   INVX1 U6373 (.Y(n9652), 
	.A(\ram[98][11] ));
   OAI22X1 U6374 (.Y(n2160), 
	.B1(n9653), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6322));
   INVX1 U6375 (.Y(n9653), 
	.A(\ram[98][10] ));
   OAI22X1 U6376 (.Y(n2159), 
	.B1(n9654), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6324));
   INVX1 U6377 (.Y(n9654), 
	.A(\ram[98][9] ));
   OAI22X1 U6378 (.Y(n2158), 
	.B1(n9655), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6326));
   INVX1 U6379 (.Y(n9655), 
	.A(\ram[98][8] ));
   OAI22X1 U6380 (.Y(n2157), 
	.B1(n9656), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6328));
   INVX1 U6381 (.Y(n9656), 
	.A(\ram[98][7] ));
   OAI22X1 U6382 (.Y(n2156), 
	.B1(n9657), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6330));
   INVX1 U6383 (.Y(n9657), 
	.A(\ram[98][6] ));
   OAI22X1 U6384 (.Y(n2155), 
	.B1(n9658), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6332));
   INVX1 U6385 (.Y(n9658), 
	.A(\ram[98][5] ));
   OAI22X1 U6386 (.Y(n2154), 
	.B1(n9659), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6334));
   INVX1 U6387 (.Y(n9659), 
	.A(\ram[98][4] ));
   OAI22X1 U6388 (.Y(n2153), 
	.B1(n9660), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6336));
   INVX1 U6389 (.Y(n9660), 
	.A(\ram[98][3] ));
   OAI22X1 U6390 (.Y(n2152), 
	.B1(n9661), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6338));
   INVX1 U6391 (.Y(n9661), 
	.A(\ram[98][2] ));
   OAI22X1 U6392 (.Y(n2151), 
	.B1(n9662), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6306));
   INVX1 U6393 (.Y(n9662), 
	.A(\ram[98][1] ));
   OAI22X1 U6394 (.Y(n2150), 
	.B1(n9663), 
	.B0(n9647), 
	.A1(n9646), 
	.A0(n6309));
   INVX1 U6395 (.Y(n9663), 
	.A(\ram[98][0] ));
   NOR2BX1 U6396 (.Y(n9647), 
	.B(n9646), 
	.AN(mem_write_en));
   NAND2X1 U6397 (.Y(n9646), 
	.B(n6476), 
	.A(n9429));
   OAI22X1 U6398 (.Y(n2149), 
	.B1(n9666), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6311));
   INVX1 U6399 (.Y(n9666), 
	.A(\ram[97][15] ));
   OAI22X1 U6400 (.Y(n2148), 
	.B1(n9667), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6314));
   INVX1 U6401 (.Y(n9667), 
	.A(\ram[97][14] ));
   OAI22X1 U6402 (.Y(n2147), 
	.B1(n9668), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6316));
   INVX1 U6403 (.Y(n9668), 
	.A(\ram[97][13] ));
   OAI22X1 U6404 (.Y(n2146), 
	.B1(n9669), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6318));
   INVX1 U6405 (.Y(n9669), 
	.A(\ram[97][12] ));
   OAI22X1 U6406 (.Y(n2145), 
	.B1(n9670), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6320));
   INVX1 U6407 (.Y(n9670), 
	.A(\ram[97][11] ));
   OAI22X1 U6408 (.Y(n2144), 
	.B1(n9671), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6322));
   INVX1 U6409 (.Y(n9671), 
	.A(\ram[97][10] ));
   OAI22X1 U6410 (.Y(n2143), 
	.B1(n9672), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6324));
   INVX1 U6411 (.Y(n9672), 
	.A(\ram[97][9] ));
   OAI22X1 U6412 (.Y(n2142), 
	.B1(n9673), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6326));
   INVX1 U6413 (.Y(n9673), 
	.A(\ram[97][8] ));
   OAI22X1 U6414 (.Y(n2141), 
	.B1(n9674), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6328));
   INVX1 U6415 (.Y(n9674), 
	.A(\ram[97][7] ));
   OAI22X1 U6416 (.Y(n2140), 
	.B1(n9675), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6330));
   INVX1 U6417 (.Y(n9675), 
	.A(\ram[97][6] ));
   OAI22X1 U6418 (.Y(n2139), 
	.B1(n9676), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6332));
   INVX1 U6419 (.Y(n9676), 
	.A(\ram[97][5] ));
   OAI22X1 U6420 (.Y(n2138), 
	.B1(n9677), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6334));
   INVX1 U6421 (.Y(n9677), 
	.A(\ram[97][4] ));
   OAI22X1 U6422 (.Y(n2137), 
	.B1(n9678), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6336));
   INVX1 U6423 (.Y(n9678), 
	.A(\ram[97][3] ));
   OAI22X1 U6424 (.Y(n2136), 
	.B1(n9679), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6338));
   INVX1 U6425 (.Y(n9679), 
	.A(\ram[97][2] ));
   OAI22X1 U6426 (.Y(n2135), 
	.B1(n9680), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6306));
   INVX1 U6427 (.Y(n9680), 
	.A(\ram[97][1] ));
   OAI22X1 U6428 (.Y(n2134), 
	.B1(n9681), 
	.B0(n9665), 
	.A1(n9664), 
	.A0(n6309));
   INVX1 U6429 (.Y(n9681), 
	.A(\ram[97][0] ));
   NOR2BX1 U6430 (.Y(n9665), 
	.B(n9664), 
	.AN(mem_write_en));
   NAND2X1 U6431 (.Y(n9664), 
	.B(n6495), 
	.A(n9429));
   OAI22X1 U6432 (.Y(n2133), 
	.B1(n9684), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6311));
   INVX1 U6433 (.Y(n9684), 
	.A(\ram[96][15] ));
   OAI22X1 U6434 (.Y(n2132), 
	.B1(n9685), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6314));
   INVX1 U6435 (.Y(n9685), 
	.A(\ram[96][14] ));
   OAI22X1 U6436 (.Y(n2131), 
	.B1(n9686), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6316));
   INVX1 U6437 (.Y(n9686), 
	.A(\ram[96][13] ));
   OAI22X1 U6438 (.Y(n2130), 
	.B1(n9687), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6318));
   INVX1 U6439 (.Y(n9687), 
	.A(\ram[96][12] ));
   OAI22X1 U6440 (.Y(n2129), 
	.B1(n9688), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6320));
   INVX1 U6441 (.Y(n9688), 
	.A(\ram[96][11] ));
   OAI22X1 U6442 (.Y(n2128), 
	.B1(n9689), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6322));
   INVX1 U6443 (.Y(n9689), 
	.A(\ram[96][10] ));
   OAI22X1 U6444 (.Y(n2127), 
	.B1(n9690), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6324));
   INVX1 U6445 (.Y(n9690), 
	.A(\ram[96][9] ));
   OAI22X1 U6446 (.Y(n2126), 
	.B1(n9691), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6326));
   INVX1 U6447 (.Y(n9691), 
	.A(\ram[96][8] ));
   OAI22X1 U6448 (.Y(n2125), 
	.B1(n9692), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6328));
   INVX1 U6449 (.Y(n9692), 
	.A(\ram[96][7] ));
   OAI22X1 U6450 (.Y(n2124), 
	.B1(n9693), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6330));
   INVX1 U6451 (.Y(n9693), 
	.A(\ram[96][6] ));
   OAI22X1 U6452 (.Y(n2123), 
	.B1(n9694), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6332));
   INVX1 U6453 (.Y(n9694), 
	.A(\ram[96][5] ));
   OAI22X1 U6454 (.Y(n2122), 
	.B1(n9695), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6334));
   INVX1 U6455 (.Y(n9695), 
	.A(\ram[96][4] ));
   OAI22X1 U6456 (.Y(n2121), 
	.B1(n9696), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6336));
   INVX1 U6457 (.Y(n9696), 
	.A(\ram[96][3] ));
   OAI22X1 U6458 (.Y(n2120), 
	.B1(n9697), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6338));
   INVX1 U6459 (.Y(n9697), 
	.A(\ram[96][2] ));
   OAI22X1 U6460 (.Y(n2119), 
	.B1(n9698), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6306));
   INVX1 U6461 (.Y(n9698), 
	.A(\ram[96][1] ));
   OAI22X1 U6462 (.Y(n2118), 
	.B1(n9699), 
	.B0(n9683), 
	.A1(n9682), 
	.A0(n6309));
   INVX1 U6463 (.Y(n9699), 
	.A(\ram[96][0] ));
   NOR2BX1 U6464 (.Y(n9683), 
	.B(n9682), 
	.AN(mem_write_en));
   NAND2X1 U6465 (.Y(n9682), 
	.B(n6514), 
	.A(n9429));
   OAI22X1 U6466 (.Y(n2117), 
	.B1(n9702), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6311));
   INVX1 U6467 (.Y(n9702), 
	.A(\ram[95][15] ));
   OAI22X1 U6468 (.Y(n2116), 
	.B1(n9703), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6314));
   INVX1 U6469 (.Y(n9703), 
	.A(\ram[95][14] ));
   OAI22X1 U6470 (.Y(n2115), 
	.B1(n9704), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6316));
   INVX1 U6471 (.Y(n9704), 
	.A(\ram[95][13] ));
   OAI22X1 U6472 (.Y(n2114), 
	.B1(n9705), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6318));
   INVX1 U6473 (.Y(n9705), 
	.A(\ram[95][12] ));
   OAI22X1 U6474 (.Y(n2113), 
	.B1(n9706), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6320));
   INVX1 U6475 (.Y(n9706), 
	.A(\ram[95][11] ));
   OAI22X1 U6476 (.Y(n2112), 
	.B1(n9707), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6322));
   INVX1 U6477 (.Y(n9707), 
	.A(\ram[95][10] ));
   OAI22X1 U6478 (.Y(n2111), 
	.B1(n9708), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6324));
   INVX1 U6479 (.Y(n9708), 
	.A(\ram[95][9] ));
   OAI22X1 U6480 (.Y(n2110), 
	.B1(n9709), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6326));
   INVX1 U6481 (.Y(n9709), 
	.A(\ram[95][8] ));
   OAI22X1 U6482 (.Y(n2109), 
	.B1(n9710), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6328));
   INVX1 U6483 (.Y(n9710), 
	.A(\ram[95][7] ));
   OAI22X1 U6484 (.Y(n2108), 
	.B1(n9711), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6330));
   INVX1 U6485 (.Y(n9711), 
	.A(\ram[95][6] ));
   OAI22X1 U6486 (.Y(n2107), 
	.B1(n9712), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6332));
   INVX1 U6487 (.Y(n9712), 
	.A(\ram[95][5] ));
   OAI22X1 U6488 (.Y(n2106), 
	.B1(n9713), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6334));
   INVX1 U6489 (.Y(n9713), 
	.A(\ram[95][4] ));
   OAI22X1 U6490 (.Y(n2105), 
	.B1(n9714), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6336));
   INVX1 U6491 (.Y(n9714), 
	.A(\ram[95][3] ));
   OAI22X1 U6492 (.Y(n2104), 
	.B1(n9715), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6338));
   INVX1 U6493 (.Y(n9715), 
	.A(\ram[95][2] ));
   OAI22X1 U6494 (.Y(n2103), 
	.B1(n9716), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6306));
   INVX1 U6495 (.Y(n9716), 
	.A(\ram[95][1] ));
   OAI22X1 U6496 (.Y(n2102), 
	.B1(n9717), 
	.B0(n9701), 
	.A1(n9700), 
	.A0(n6309));
   INVX1 U6497 (.Y(n9717), 
	.A(\ram[95][0] ));
   NOR2BX1 U6498 (.Y(n9701), 
	.B(n9700), 
	.AN(mem_write_en));
   NAND2X1 U6499 (.Y(n9700), 
	.B(n6533), 
	.A(n9718));
   OAI22X1 U6500 (.Y(n2101), 
	.B1(n9721), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6311));
   INVX1 U6501 (.Y(n9721), 
	.A(\ram[94][15] ));
   OAI22X1 U6502 (.Y(n2100), 
	.B1(n9722), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6314));
   INVX1 U6503 (.Y(n9722), 
	.A(\ram[94][14] ));
   OAI22X1 U6504 (.Y(n2099), 
	.B1(n9723), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6316));
   INVX1 U6505 (.Y(n9723), 
	.A(\ram[94][13] ));
   OAI22X1 U6506 (.Y(n2098), 
	.B1(n9724), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6318));
   INVX1 U6507 (.Y(n9724), 
	.A(\ram[94][12] ));
   OAI22X1 U6508 (.Y(n2097), 
	.B1(n9725), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6320));
   INVX1 U6509 (.Y(n9725), 
	.A(\ram[94][11] ));
   OAI22X1 U6510 (.Y(n2096), 
	.B1(n9726), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6322));
   INVX1 U6511 (.Y(n9726), 
	.A(\ram[94][10] ));
   OAI22X1 U6512 (.Y(n2095), 
	.B1(n9727), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6324));
   INVX1 U6513 (.Y(n9727), 
	.A(\ram[94][9] ));
   OAI22X1 U6514 (.Y(n2094), 
	.B1(n9728), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6326));
   INVX1 U6515 (.Y(n9728), 
	.A(\ram[94][8] ));
   OAI22X1 U6516 (.Y(n2093), 
	.B1(n9729), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6328));
   INVX1 U6517 (.Y(n9729), 
	.A(\ram[94][7] ));
   OAI22X1 U6518 (.Y(n2092), 
	.B1(n9730), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6330));
   INVX1 U6519 (.Y(n9730), 
	.A(\ram[94][6] ));
   OAI22X1 U6520 (.Y(n2091), 
	.B1(n9731), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6332));
   INVX1 U6521 (.Y(n9731), 
	.A(\ram[94][5] ));
   OAI22X1 U6522 (.Y(n2090), 
	.B1(n9732), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6334));
   INVX1 U6523 (.Y(n9732), 
	.A(\ram[94][4] ));
   OAI22X1 U6524 (.Y(n2089), 
	.B1(n9733), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6336));
   INVX1 U6525 (.Y(n9733), 
	.A(\ram[94][3] ));
   OAI22X1 U6526 (.Y(n2088), 
	.B1(n9734), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6338));
   INVX1 U6527 (.Y(n9734), 
	.A(\ram[94][2] ));
   OAI22X1 U6528 (.Y(n2087), 
	.B1(n9735), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6306));
   INVX1 U6529 (.Y(n9735), 
	.A(\ram[94][1] ));
   OAI22X1 U6530 (.Y(n2086), 
	.B1(n9736), 
	.B0(n9720), 
	.A1(n9719), 
	.A0(n6309));
   INVX1 U6531 (.Y(n9736), 
	.A(\ram[94][0] ));
   NOR2BX1 U6532 (.Y(n9720), 
	.B(n9719), 
	.AN(mem_write_en));
   NAND2X1 U6533 (.Y(n9719), 
	.B(n6553), 
	.A(n9718));
   OAI22X1 U6534 (.Y(n2085), 
	.B1(n9739), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6311));
   INVX1 U6535 (.Y(n9739), 
	.A(\ram[93][15] ));
   OAI22X1 U6536 (.Y(n2084), 
	.B1(n9740), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6314));
   INVX1 U6537 (.Y(n9740), 
	.A(\ram[93][14] ));
   OAI22X1 U6538 (.Y(n2083), 
	.B1(n9741), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6316));
   INVX1 U6539 (.Y(n9741), 
	.A(\ram[93][13] ));
   OAI22X1 U6540 (.Y(n2082), 
	.B1(n9742), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6318));
   INVX1 U6541 (.Y(n9742), 
	.A(\ram[93][12] ));
   OAI22X1 U6542 (.Y(n2081), 
	.B1(n9743), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6320));
   INVX1 U6543 (.Y(n9743), 
	.A(\ram[93][11] ));
   OAI22X1 U6544 (.Y(n2080), 
	.B1(n9744), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6322));
   INVX1 U6545 (.Y(n9744), 
	.A(\ram[93][10] ));
   OAI22X1 U6546 (.Y(n2079), 
	.B1(n9745), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6324));
   INVX1 U6547 (.Y(n9745), 
	.A(\ram[93][9] ));
   OAI22X1 U6548 (.Y(n2078), 
	.B1(n9746), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6326));
   INVX1 U6549 (.Y(n9746), 
	.A(\ram[93][8] ));
   OAI22X1 U6550 (.Y(n2077), 
	.B1(n9747), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6328));
   INVX1 U6551 (.Y(n9747), 
	.A(\ram[93][7] ));
   OAI22X1 U6552 (.Y(n2076), 
	.B1(n9748), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6330));
   INVX1 U6553 (.Y(n9748), 
	.A(\ram[93][6] ));
   OAI22X1 U6554 (.Y(n2075), 
	.B1(n9749), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6332));
   INVX1 U6555 (.Y(n9749), 
	.A(\ram[93][5] ));
   OAI22X1 U6556 (.Y(n2074), 
	.B1(n9750), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6334));
   INVX1 U6557 (.Y(n9750), 
	.A(\ram[93][4] ));
   OAI22X1 U6558 (.Y(n2073), 
	.B1(n9751), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6336));
   INVX1 U6559 (.Y(n9751), 
	.A(\ram[93][3] ));
   OAI22X1 U6560 (.Y(n2072), 
	.B1(n9752), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6338));
   INVX1 U6561 (.Y(n9752), 
	.A(\ram[93][2] ));
   OAI22X1 U6562 (.Y(n2071), 
	.B1(n9753), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6306));
   INVX1 U6563 (.Y(n9753), 
	.A(\ram[93][1] ));
   OAI22X1 U6564 (.Y(n2070), 
	.B1(n9754), 
	.B0(n9738), 
	.A1(n9737), 
	.A0(n6309));
   INVX1 U6565 (.Y(n9754), 
	.A(\ram[93][0] ));
   NOR2BX1 U6566 (.Y(n9738), 
	.B(n9737), 
	.AN(mem_write_en));
   NAND2X1 U6567 (.Y(n9737), 
	.B(n6572), 
	.A(n9718));
   OAI22X1 U6568 (.Y(n2069), 
	.B1(n9757), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6311));
   INVX1 U6569 (.Y(n9757), 
	.A(\ram[92][15] ));
   OAI22X1 U6570 (.Y(n2068), 
	.B1(n9758), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6314));
   INVX1 U6571 (.Y(n9758), 
	.A(\ram[92][14] ));
   OAI22X1 U6572 (.Y(n2067), 
	.B1(n9759), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6316));
   INVX1 U6573 (.Y(n9759), 
	.A(\ram[92][13] ));
   OAI22X1 U6574 (.Y(n2066), 
	.B1(n9760), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6318));
   INVX1 U6575 (.Y(n9760), 
	.A(\ram[92][12] ));
   OAI22X1 U6576 (.Y(n2065), 
	.B1(n9761), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6320));
   INVX1 U6577 (.Y(n9761), 
	.A(\ram[92][11] ));
   OAI22X1 U6578 (.Y(n2064), 
	.B1(n9762), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6322));
   INVX1 U6579 (.Y(n9762), 
	.A(\ram[92][10] ));
   OAI22X1 U6580 (.Y(n2063), 
	.B1(n9763), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6324));
   INVX1 U6581 (.Y(n9763), 
	.A(\ram[92][9] ));
   OAI22X1 U6582 (.Y(n2062), 
	.B1(n9764), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6326));
   INVX1 U6583 (.Y(n9764), 
	.A(\ram[92][8] ));
   OAI22X1 U6584 (.Y(n2061), 
	.B1(n9765), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6328));
   INVX1 U6585 (.Y(n9765), 
	.A(\ram[92][7] ));
   OAI22X1 U6586 (.Y(n2060), 
	.B1(n9766), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6330));
   INVX1 U6587 (.Y(n9766), 
	.A(\ram[92][6] ));
   OAI22X1 U6588 (.Y(n2059), 
	.B1(n9767), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6332));
   INVX1 U6589 (.Y(n9767), 
	.A(\ram[92][5] ));
   OAI22X1 U6590 (.Y(n2058), 
	.B1(n9768), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6334));
   INVX1 U6591 (.Y(n9768), 
	.A(\ram[92][4] ));
   OAI22X1 U6592 (.Y(n2057), 
	.B1(n9769), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6336));
   INVX1 U6593 (.Y(n9769), 
	.A(\ram[92][3] ));
   OAI22X1 U6594 (.Y(n2056), 
	.B1(n9770), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6338));
   INVX1 U6595 (.Y(n9770), 
	.A(\ram[92][2] ));
   OAI22X1 U6596 (.Y(n2055), 
	.B1(n9771), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6306));
   INVX1 U6597 (.Y(n9771), 
	.A(\ram[92][1] ));
   OAI22X1 U6598 (.Y(n2054), 
	.B1(n9772), 
	.B0(n9756), 
	.A1(n9755), 
	.A0(n6309));
   INVX1 U6599 (.Y(n9772), 
	.A(\ram[92][0] ));
   NOR2BX1 U6600 (.Y(n9756), 
	.B(n9755), 
	.AN(mem_write_en));
   NAND2X1 U6601 (.Y(n9755), 
	.B(n6591), 
	.A(n9718));
   OAI22X1 U6602 (.Y(n2053), 
	.B1(n9775), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6311));
   INVX1 U6603 (.Y(n9775), 
	.A(\ram[91][15] ));
   OAI22X1 U6604 (.Y(n2052), 
	.B1(n9776), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6314));
   INVX1 U6605 (.Y(n9776), 
	.A(\ram[91][14] ));
   OAI22X1 U6606 (.Y(n2051), 
	.B1(n9777), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6316));
   INVX1 U6607 (.Y(n9777), 
	.A(\ram[91][13] ));
   OAI22X1 U6608 (.Y(n2050), 
	.B1(n9778), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6318));
   INVX1 U6609 (.Y(n9778), 
	.A(\ram[91][12] ));
   OAI22X1 U6610 (.Y(n2049), 
	.B1(n9779), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6320));
   INVX1 U6611 (.Y(n9779), 
	.A(\ram[91][11] ));
   OAI22X1 U6612 (.Y(n2048), 
	.B1(n9780), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6322));
   INVX1 U6613 (.Y(n9780), 
	.A(\ram[91][10] ));
   OAI22X1 U6614 (.Y(n2047), 
	.B1(n9781), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6324));
   INVX1 U6615 (.Y(n9781), 
	.A(\ram[91][9] ));
   OAI22X1 U6616 (.Y(n2046), 
	.B1(n9782), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6326));
   INVX1 U6617 (.Y(n9782), 
	.A(\ram[91][8] ));
   OAI22X1 U6618 (.Y(n2045), 
	.B1(n9783), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6328));
   INVX1 U6619 (.Y(n9783), 
	.A(\ram[91][7] ));
   OAI22X1 U6620 (.Y(n2044), 
	.B1(n9784), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6330));
   INVX1 U6621 (.Y(n9784), 
	.A(\ram[91][6] ));
   OAI22X1 U6622 (.Y(n2043), 
	.B1(n9785), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6332));
   INVX1 U6623 (.Y(n9785), 
	.A(\ram[91][5] ));
   OAI22X1 U6624 (.Y(n2042), 
	.B1(n9786), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6334));
   INVX1 U6625 (.Y(n9786), 
	.A(\ram[91][4] ));
   OAI22X1 U6626 (.Y(n2041), 
	.B1(n9787), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6336));
   INVX1 U6627 (.Y(n9787), 
	.A(\ram[91][3] ));
   OAI22X1 U6628 (.Y(n2040), 
	.B1(n9788), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6338));
   INVX1 U6629 (.Y(n9788), 
	.A(\ram[91][2] ));
   OAI22X1 U6630 (.Y(n2039), 
	.B1(n9789), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6306));
   INVX1 U6631 (.Y(n9789), 
	.A(\ram[91][1] ));
   OAI22X1 U6632 (.Y(n2038), 
	.B1(n9790), 
	.B0(n9774), 
	.A1(n9773), 
	.A0(n6309));
   INVX1 U6633 (.Y(n9790), 
	.A(\ram[91][0] ));
   NOR2BX1 U6634 (.Y(n9774), 
	.B(n9773), 
	.AN(mem_write_en));
   NAND2X1 U6635 (.Y(n9773), 
	.B(n6610), 
	.A(n9718));
   OAI22X1 U6636 (.Y(n2037), 
	.B1(n9793), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6311));
   INVX1 U6637 (.Y(n9793), 
	.A(\ram[90][15] ));
   OAI22X1 U6638 (.Y(n2036), 
	.B1(n9794), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6314));
   INVX1 U6639 (.Y(n9794), 
	.A(\ram[90][14] ));
   OAI22X1 U6640 (.Y(n2035), 
	.B1(n9795), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6316));
   INVX1 U6641 (.Y(n9795), 
	.A(\ram[90][13] ));
   OAI22X1 U6642 (.Y(n2034), 
	.B1(n9796), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6318));
   INVX1 U6643 (.Y(n9796), 
	.A(\ram[90][12] ));
   OAI22X1 U6644 (.Y(n2033), 
	.B1(n9797), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6320));
   INVX1 U6645 (.Y(n9797), 
	.A(\ram[90][11] ));
   OAI22X1 U6646 (.Y(n2032), 
	.B1(n9798), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6322));
   INVX1 U6647 (.Y(n9798), 
	.A(\ram[90][10] ));
   OAI22X1 U6648 (.Y(n2031), 
	.B1(n9799), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6324));
   INVX1 U6649 (.Y(n9799), 
	.A(\ram[90][9] ));
   OAI22X1 U6650 (.Y(n2030), 
	.B1(n9800), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6326));
   INVX1 U6651 (.Y(n9800), 
	.A(\ram[90][8] ));
   OAI22X1 U6652 (.Y(n2029), 
	.B1(n9801), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6328));
   INVX1 U6653 (.Y(n9801), 
	.A(\ram[90][7] ));
   OAI22X1 U6654 (.Y(n2028), 
	.B1(n9802), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6330));
   INVX1 U6655 (.Y(n9802), 
	.A(\ram[90][6] ));
   OAI22X1 U6656 (.Y(n2027), 
	.B1(n9803), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6332));
   INVX1 U6657 (.Y(n9803), 
	.A(\ram[90][5] ));
   OAI22X1 U6658 (.Y(n2026), 
	.B1(n9804), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6334));
   INVX1 U6659 (.Y(n9804), 
	.A(\ram[90][4] ));
   OAI22X1 U6660 (.Y(n2025), 
	.B1(n9805), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6336));
   INVX1 U6661 (.Y(n9805), 
	.A(\ram[90][3] ));
   OAI22X1 U6662 (.Y(n2024), 
	.B1(n9806), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6338));
   INVX1 U6663 (.Y(n9806), 
	.A(\ram[90][2] ));
   OAI22X1 U6664 (.Y(n2023), 
	.B1(n9807), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6306));
   INVX1 U6665 (.Y(n9807), 
	.A(\ram[90][1] ));
   OAI22X1 U6666 (.Y(n2022), 
	.B1(n9808), 
	.B0(n9792), 
	.A1(n9791), 
	.A0(n6309));
   INVX1 U6667 (.Y(n9808), 
	.A(\ram[90][0] ));
   NOR2BX1 U6668 (.Y(n9792), 
	.B(n9791), 
	.AN(mem_write_en));
   NAND2X1 U6669 (.Y(n9791), 
	.B(n6629), 
	.A(n9718));
   OAI22X1 U6670 (.Y(n2021), 
	.B1(n9811), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6311));
   INVX1 U6671 (.Y(n9811), 
	.A(\ram[89][15] ));
   OAI22X1 U6672 (.Y(n2020), 
	.B1(n9812), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6314));
   INVX1 U6673 (.Y(n9812), 
	.A(\ram[89][14] ));
   OAI22X1 U6674 (.Y(n2019), 
	.B1(n9813), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6316));
   INVX1 U6675 (.Y(n9813), 
	.A(\ram[89][13] ));
   OAI22X1 U6676 (.Y(n2018), 
	.B1(n9814), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6318));
   INVX1 U6677 (.Y(n9814), 
	.A(\ram[89][12] ));
   OAI22X1 U6678 (.Y(n2017), 
	.B1(n9815), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6320));
   INVX1 U6679 (.Y(n9815), 
	.A(\ram[89][11] ));
   OAI22X1 U6680 (.Y(n2016), 
	.B1(n9816), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6322));
   INVX1 U6681 (.Y(n9816), 
	.A(\ram[89][10] ));
   OAI22X1 U6682 (.Y(n2015), 
	.B1(n9817), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6324));
   INVX1 U6683 (.Y(n9817), 
	.A(\ram[89][9] ));
   OAI22X1 U6684 (.Y(n2014), 
	.B1(n9818), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6326));
   INVX1 U6685 (.Y(n9818), 
	.A(\ram[89][8] ));
   OAI22X1 U6686 (.Y(n2013), 
	.B1(n9819), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6328));
   INVX1 U6687 (.Y(n9819), 
	.A(\ram[89][7] ));
   OAI22X1 U6688 (.Y(n2012), 
	.B1(n9820), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6330));
   INVX1 U6689 (.Y(n9820), 
	.A(\ram[89][6] ));
   OAI22X1 U6690 (.Y(n2011), 
	.B1(n9821), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6332));
   INVX1 U6691 (.Y(n9821), 
	.A(\ram[89][5] ));
   OAI22X1 U6692 (.Y(n2010), 
	.B1(n9822), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6334));
   INVX1 U6693 (.Y(n9822), 
	.A(\ram[89][4] ));
   OAI22X1 U6694 (.Y(n2009), 
	.B1(n9823), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6336));
   INVX1 U6695 (.Y(n9823), 
	.A(\ram[89][3] ));
   OAI22X1 U6696 (.Y(n2008), 
	.B1(n9824), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6338));
   INVX1 U6697 (.Y(n9824), 
	.A(\ram[89][2] ));
   OAI22X1 U6698 (.Y(n2007), 
	.B1(n9825), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6306));
   INVX1 U6699 (.Y(n9825), 
	.A(\ram[89][1] ));
   OAI22X1 U6700 (.Y(n2006), 
	.B1(n9826), 
	.B0(n9810), 
	.A1(n9809), 
	.A0(n6309));
   INVX1 U6701 (.Y(n9826), 
	.A(\ram[89][0] ));
   NOR2BX1 U6702 (.Y(n9810), 
	.B(n9809), 
	.AN(mem_write_en));
   NAND2X1 U6703 (.Y(n9809), 
	.B(n6342), 
	.A(n9718));
   OAI22X1 U6704 (.Y(n2005), 
	.B1(n9829), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6311));
   INVX1 U6705 (.Y(n9829), 
	.A(\ram[88][15] ));
   OAI22X1 U6706 (.Y(n2004), 
	.B1(n9830), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6314));
   INVX1 U6707 (.Y(n9830), 
	.A(\ram[88][14] ));
   OAI22X1 U6708 (.Y(n2003), 
	.B1(n9831), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6316));
   INVX1 U6709 (.Y(n9831), 
	.A(\ram[88][13] ));
   OAI22X1 U6710 (.Y(n2002), 
	.B1(n9832), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6318));
   INVX1 U6711 (.Y(n9832), 
	.A(\ram[88][12] ));
   OAI22X1 U6712 (.Y(n2001), 
	.B1(n9833), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6320));
   INVX1 U6713 (.Y(n9833), 
	.A(\ram[88][11] ));
   OAI22X1 U6714 (.Y(n2000), 
	.B1(n9834), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6322));
   INVX1 U6715 (.Y(n9834), 
	.A(\ram[88][10] ));
   OAI22X1 U6716 (.Y(n1999), 
	.B1(n9835), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6324));
   INVX1 U6717 (.Y(n9835), 
	.A(\ram[88][9] ));
   OAI22X1 U6718 (.Y(n1998), 
	.B1(n9836), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6326));
   INVX1 U6719 (.Y(n9836), 
	.A(\ram[88][8] ));
   OAI22X1 U6720 (.Y(n1997), 
	.B1(n9837), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6328));
   INVX1 U6721 (.Y(n9837), 
	.A(\ram[88][7] ));
   OAI22X1 U6722 (.Y(n1996), 
	.B1(n9838), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6330));
   INVX1 U6723 (.Y(n9838), 
	.A(\ram[88][6] ));
   OAI22X1 U6724 (.Y(n1995), 
	.B1(n9839), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6332));
   INVX1 U6725 (.Y(n9839), 
	.A(\ram[88][5] ));
   OAI22X1 U6726 (.Y(n1994), 
	.B1(n9840), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6334));
   INVX1 U6727 (.Y(n9840), 
	.A(\ram[88][4] ));
   OAI22X1 U6728 (.Y(n1993), 
	.B1(n9841), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6336));
   INVX1 U6729 (.Y(n9841), 
	.A(\ram[88][3] ));
   OAI22X1 U6730 (.Y(n1992), 
	.B1(n9842), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6338));
   INVX1 U6731 (.Y(n9842), 
	.A(\ram[88][2] ));
   OAI22X1 U6732 (.Y(n1991), 
	.B1(n9843), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6306));
   INVX1 U6733 (.Y(n9843), 
	.A(\ram[88][1] ));
   OAI22X1 U6734 (.Y(n1990), 
	.B1(n9844), 
	.B0(n9828), 
	.A1(n9827), 
	.A0(n6309));
   INVX1 U6735 (.Y(n9844), 
	.A(\ram[88][0] ));
   NOR2BX1 U6736 (.Y(n9828), 
	.B(n9827), 
	.AN(mem_write_en));
   NAND2X1 U6737 (.Y(n9827), 
	.B(n6362), 
	.A(n9718));
   OAI22X1 U6738 (.Y(n1989), 
	.B1(n9847), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6311));
   INVX1 U6739 (.Y(n9847), 
	.A(\ram[87][15] ));
   OAI22X1 U6740 (.Y(n1988), 
	.B1(n9848), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6314));
   INVX1 U6741 (.Y(n9848), 
	.A(\ram[87][14] ));
   OAI22X1 U6742 (.Y(n1987), 
	.B1(n9849), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6316));
   INVX1 U6743 (.Y(n9849), 
	.A(\ram[87][13] ));
   OAI22X1 U6744 (.Y(n1986), 
	.B1(n9850), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6318));
   INVX1 U6745 (.Y(n9850), 
	.A(\ram[87][12] ));
   OAI22X1 U6746 (.Y(n1985), 
	.B1(n9851), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6320));
   INVX1 U6747 (.Y(n9851), 
	.A(\ram[87][11] ));
   OAI22X1 U6748 (.Y(n1984), 
	.B1(n9852), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6322));
   INVX1 U6749 (.Y(n9852), 
	.A(\ram[87][10] ));
   OAI22X1 U6750 (.Y(n1983), 
	.B1(n9853), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6324));
   INVX1 U6751 (.Y(n9853), 
	.A(\ram[87][9] ));
   OAI22X1 U6752 (.Y(n1982), 
	.B1(n9854), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6326));
   INVX1 U6753 (.Y(n9854), 
	.A(\ram[87][8] ));
   OAI22X1 U6754 (.Y(n1981), 
	.B1(n9855), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6328));
   INVX1 U6755 (.Y(n9855), 
	.A(\ram[87][7] ));
   OAI22X1 U6756 (.Y(n1980), 
	.B1(n9856), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6330));
   INVX1 U6757 (.Y(n9856), 
	.A(\ram[87][6] ));
   OAI22X1 U6758 (.Y(n1979), 
	.B1(n9857), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6332));
   INVX1 U6759 (.Y(n9857), 
	.A(\ram[87][5] ));
   OAI22X1 U6760 (.Y(n1978), 
	.B1(n9858), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6334));
   INVX1 U6761 (.Y(n9858), 
	.A(\ram[87][4] ));
   OAI22X1 U6762 (.Y(n1977), 
	.B1(n9859), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6336));
   INVX1 U6763 (.Y(n9859), 
	.A(\ram[87][3] ));
   OAI22X1 U6764 (.Y(n1976), 
	.B1(n9860), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6338));
   INVX1 U6765 (.Y(n9860), 
	.A(\ram[87][2] ));
   OAI22X1 U6766 (.Y(n1975), 
	.B1(n9861), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6306));
   INVX1 U6767 (.Y(n9861), 
	.A(\ram[87][1] ));
   OAI22X1 U6768 (.Y(n1974), 
	.B1(n9862), 
	.B0(n9846), 
	.A1(n9845), 
	.A0(n6309));
   INVX1 U6769 (.Y(n9862), 
	.A(\ram[87][0] ));
   NOR2BX1 U6770 (.Y(n9846), 
	.B(n9845), 
	.AN(mem_write_en));
   NAND2X1 U6771 (.Y(n9845), 
	.B(n6381), 
	.A(n9718));
   OAI22X1 U6772 (.Y(n1973), 
	.B1(n9865), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6311));
   INVX1 U6773 (.Y(n9865), 
	.A(\ram[86][15] ));
   OAI22X1 U6774 (.Y(n1972), 
	.B1(n9866), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6314));
   INVX1 U6775 (.Y(n9866), 
	.A(\ram[86][14] ));
   OAI22X1 U6776 (.Y(n1971), 
	.B1(n9867), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6316));
   INVX1 U6777 (.Y(n9867), 
	.A(\ram[86][13] ));
   OAI22X1 U6778 (.Y(n1970), 
	.B1(n9868), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6318));
   INVX1 U6779 (.Y(n9868), 
	.A(\ram[86][12] ));
   OAI22X1 U6780 (.Y(n1969), 
	.B1(n9869), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6320));
   INVX1 U6781 (.Y(n9869), 
	.A(\ram[86][11] ));
   OAI22X1 U6782 (.Y(n1968), 
	.B1(n9870), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6322));
   INVX1 U6783 (.Y(n9870), 
	.A(\ram[86][10] ));
   OAI22X1 U6784 (.Y(n1967), 
	.B1(n9871), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6324));
   INVX1 U6785 (.Y(n9871), 
	.A(\ram[86][9] ));
   OAI22X1 U6786 (.Y(n1966), 
	.B1(n9872), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6326));
   INVX1 U6787 (.Y(n9872), 
	.A(\ram[86][8] ));
   OAI22X1 U6788 (.Y(n1965), 
	.B1(n9873), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6328));
   INVX1 U6789 (.Y(n9873), 
	.A(\ram[86][7] ));
   OAI22X1 U6790 (.Y(n1964), 
	.B1(n9874), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6330));
   INVX1 U6791 (.Y(n9874), 
	.A(\ram[86][6] ));
   OAI22X1 U6792 (.Y(n1963), 
	.B1(n9875), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6332));
   INVX1 U6793 (.Y(n9875), 
	.A(\ram[86][5] ));
   OAI22X1 U6794 (.Y(n1962), 
	.B1(n9876), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6334));
   INVX1 U6795 (.Y(n9876), 
	.A(\ram[86][4] ));
   OAI22X1 U6796 (.Y(n1961), 
	.B1(n9877), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6336));
   INVX1 U6797 (.Y(n9877), 
	.A(\ram[86][3] ));
   OAI22X1 U6798 (.Y(n1960), 
	.B1(n9878), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6338));
   INVX1 U6799 (.Y(n9878), 
	.A(\ram[86][2] ));
   OAI22X1 U6800 (.Y(n1959), 
	.B1(n9879), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6306));
   INVX1 U6801 (.Y(n9879), 
	.A(\ram[86][1] ));
   OAI22X1 U6802 (.Y(n1958), 
	.B1(n9880), 
	.B0(n9864), 
	.A1(n9863), 
	.A0(n6309));
   INVX1 U6803 (.Y(n9880), 
	.A(\ram[86][0] ));
   NOR2BX1 U6804 (.Y(n9864), 
	.B(n9863), 
	.AN(mem_write_en));
   NAND2X1 U6805 (.Y(n9863), 
	.B(n6400), 
	.A(n9718));
   OAI22X1 U6806 (.Y(n1957), 
	.B1(n9883), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6311));
   INVX1 U6807 (.Y(n9883), 
	.A(\ram[85][15] ));
   OAI22X1 U6808 (.Y(n1956), 
	.B1(n9884), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6314));
   INVX1 U6809 (.Y(n9884), 
	.A(\ram[85][14] ));
   OAI22X1 U6810 (.Y(n1955), 
	.B1(n9885), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6316));
   INVX1 U6811 (.Y(n9885), 
	.A(\ram[85][13] ));
   OAI22X1 U6812 (.Y(n1954), 
	.B1(n9886), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6318));
   INVX1 U6813 (.Y(n9886), 
	.A(\ram[85][12] ));
   OAI22X1 U6814 (.Y(n1953), 
	.B1(n9887), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6320));
   INVX1 U6815 (.Y(n9887), 
	.A(\ram[85][11] ));
   OAI22X1 U6816 (.Y(n1952), 
	.B1(n9888), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6322));
   INVX1 U6817 (.Y(n9888), 
	.A(\ram[85][10] ));
   OAI22X1 U6818 (.Y(n1951), 
	.B1(n9889), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6324));
   INVX1 U6819 (.Y(n9889), 
	.A(\ram[85][9] ));
   OAI22X1 U6820 (.Y(n1950), 
	.B1(n9890), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6326));
   INVX1 U6821 (.Y(n9890), 
	.A(\ram[85][8] ));
   OAI22X1 U6822 (.Y(n1949), 
	.B1(n9891), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6328));
   INVX1 U6823 (.Y(n9891), 
	.A(\ram[85][7] ));
   OAI22X1 U6824 (.Y(n1948), 
	.B1(n9892), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6330));
   INVX1 U6825 (.Y(n9892), 
	.A(\ram[85][6] ));
   OAI22X1 U6826 (.Y(n1947), 
	.B1(n9893), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6332));
   INVX1 U6827 (.Y(n9893), 
	.A(\ram[85][5] ));
   OAI22X1 U6828 (.Y(n1946), 
	.B1(n9894), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6334));
   INVX1 U6829 (.Y(n9894), 
	.A(\ram[85][4] ));
   OAI22X1 U6830 (.Y(n1945), 
	.B1(n9895), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6336));
   INVX1 U6831 (.Y(n9895), 
	.A(\ram[85][3] ));
   OAI22X1 U6832 (.Y(n1944), 
	.B1(n9896), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6338));
   INVX1 U6833 (.Y(n9896), 
	.A(\ram[85][2] ));
   OAI22X1 U6834 (.Y(n1943), 
	.B1(n9897), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6306));
   INVX1 U6835 (.Y(n9897), 
	.A(\ram[85][1] ));
   OAI22X1 U6836 (.Y(n1942), 
	.B1(n9898), 
	.B0(n9882), 
	.A1(n9881), 
	.A0(n6309));
   INVX1 U6837 (.Y(n9898), 
	.A(\ram[85][0] ));
   NOR2BX1 U6838 (.Y(n9882), 
	.B(n9881), 
	.AN(mem_write_en));
   NAND2X1 U6839 (.Y(n9881), 
	.B(n6419), 
	.A(n9718));
   OAI22X1 U6840 (.Y(n1941), 
	.B1(n9901), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6311));
   INVX1 U6841 (.Y(n9901), 
	.A(\ram[84][15] ));
   OAI22X1 U6842 (.Y(n1940), 
	.B1(n9902), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6314));
   INVX1 U6843 (.Y(n9902), 
	.A(\ram[84][14] ));
   OAI22X1 U6844 (.Y(n1939), 
	.B1(n9903), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6316));
   INVX1 U6845 (.Y(n9903), 
	.A(\ram[84][13] ));
   OAI22X1 U6846 (.Y(n1938), 
	.B1(n9904), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6318));
   INVX1 U6847 (.Y(n9904), 
	.A(\ram[84][12] ));
   OAI22X1 U6848 (.Y(n1937), 
	.B1(n9905), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6320));
   INVX1 U6849 (.Y(n9905), 
	.A(\ram[84][11] ));
   OAI22X1 U6850 (.Y(n1936), 
	.B1(n9906), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6322));
   INVX1 U6851 (.Y(n9906), 
	.A(\ram[84][10] ));
   OAI22X1 U6852 (.Y(n1935), 
	.B1(n9907), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6324));
   INVX1 U6853 (.Y(n9907), 
	.A(\ram[84][9] ));
   OAI22X1 U6854 (.Y(n1934), 
	.B1(n9908), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6326));
   INVX1 U6855 (.Y(n9908), 
	.A(\ram[84][8] ));
   OAI22X1 U6856 (.Y(n1933), 
	.B1(n9909), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6328));
   INVX1 U6857 (.Y(n9909), 
	.A(\ram[84][7] ));
   OAI22X1 U6858 (.Y(n1932), 
	.B1(n9910), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6330));
   INVX1 U6859 (.Y(n9910), 
	.A(\ram[84][6] ));
   OAI22X1 U6860 (.Y(n1931), 
	.B1(n9911), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6332));
   INVX1 U6861 (.Y(n9911), 
	.A(\ram[84][5] ));
   OAI22X1 U6862 (.Y(n1930), 
	.B1(n9912), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6334));
   INVX1 U6863 (.Y(n9912), 
	.A(\ram[84][4] ));
   OAI22X1 U6864 (.Y(n1929), 
	.B1(n9913), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6336));
   INVX1 U6865 (.Y(n9913), 
	.A(\ram[84][3] ));
   OAI22X1 U6866 (.Y(n1928), 
	.B1(n9914), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6338));
   INVX1 U6867 (.Y(n9914), 
	.A(\ram[84][2] ));
   OAI22X1 U6868 (.Y(n1927), 
	.B1(n9915), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6306));
   INVX1 U6869 (.Y(n9915), 
	.A(\ram[84][1] ));
   OAI22X1 U6870 (.Y(n1926), 
	.B1(n9916), 
	.B0(n9900), 
	.A1(n9899), 
	.A0(n6309));
   INVX1 U6871 (.Y(n9916), 
	.A(\ram[84][0] ));
   NOR2BX1 U6872 (.Y(n9900), 
	.B(n9899), 
	.AN(mem_write_en));
   NAND2X1 U6873 (.Y(n9899), 
	.B(n6438), 
	.A(n9718));
   OAI22X1 U6874 (.Y(n1925), 
	.B1(n9919), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6311));
   INVX1 U6875 (.Y(n9919), 
	.A(\ram[83][15] ));
   OAI22X1 U6876 (.Y(n1924), 
	.B1(n9920), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6314));
   INVX1 U6877 (.Y(n9920), 
	.A(\ram[83][14] ));
   OAI22X1 U6878 (.Y(n1923), 
	.B1(n9921), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6316));
   INVX1 U6879 (.Y(n9921), 
	.A(\ram[83][13] ));
   OAI22X1 U6880 (.Y(n1922), 
	.B1(n9922), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6318));
   INVX1 U6881 (.Y(n9922), 
	.A(\ram[83][12] ));
   OAI22X1 U6882 (.Y(n1921), 
	.B1(n9923), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6320));
   INVX1 U6883 (.Y(n9923), 
	.A(\ram[83][11] ));
   OAI22X1 U6884 (.Y(n1920), 
	.B1(n9924), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6322));
   INVX1 U6885 (.Y(n9924), 
	.A(\ram[83][10] ));
   OAI22X1 U6886 (.Y(n1919), 
	.B1(n9925), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6324));
   INVX1 U6887 (.Y(n9925), 
	.A(\ram[83][9] ));
   OAI22X1 U6888 (.Y(n1918), 
	.B1(n9926), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6326));
   INVX1 U6889 (.Y(n9926), 
	.A(\ram[83][8] ));
   OAI22X1 U6890 (.Y(n1917), 
	.B1(n9927), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6328));
   INVX1 U6891 (.Y(n9927), 
	.A(\ram[83][7] ));
   OAI22X1 U6892 (.Y(n1916), 
	.B1(n9928), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6330));
   INVX1 U6893 (.Y(n9928), 
	.A(\ram[83][6] ));
   OAI22X1 U6894 (.Y(n1915), 
	.B1(n9929), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6332));
   INVX1 U6895 (.Y(n9929), 
	.A(\ram[83][5] ));
   OAI22X1 U6896 (.Y(n1914), 
	.B1(n9930), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6334));
   INVX1 U6897 (.Y(n9930), 
	.A(\ram[83][4] ));
   OAI22X1 U6898 (.Y(n1913), 
	.B1(n9931), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6336));
   INVX1 U6899 (.Y(n9931), 
	.A(\ram[83][3] ));
   OAI22X1 U6900 (.Y(n1912), 
	.B1(n9932), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6338));
   INVX1 U6901 (.Y(n9932), 
	.A(\ram[83][2] ));
   OAI22X1 U6902 (.Y(n1911), 
	.B1(n9933), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6306));
   INVX1 U6903 (.Y(n9933), 
	.A(\ram[83][1] ));
   OAI22X1 U6904 (.Y(n1910), 
	.B1(n9934), 
	.B0(n9918), 
	.A1(n9917), 
	.A0(n6309));
   INVX1 U6905 (.Y(n9934), 
	.A(\ram[83][0] ));
   NOR2BX1 U6906 (.Y(n9918), 
	.B(n9917), 
	.AN(mem_write_en));
   NAND2X1 U6907 (.Y(n9917), 
	.B(n6457), 
	.A(n9718));
   OAI22X1 U6908 (.Y(n1909), 
	.B1(n9937), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6311));
   INVX1 U6909 (.Y(n9937), 
	.A(\ram[82][15] ));
   OAI22X1 U6910 (.Y(n1908), 
	.B1(n9938), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6314));
   INVX1 U6911 (.Y(n9938), 
	.A(\ram[82][14] ));
   OAI22X1 U6912 (.Y(n1907), 
	.B1(n9939), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6316));
   INVX1 U6913 (.Y(n9939), 
	.A(\ram[82][13] ));
   OAI22X1 U6914 (.Y(n1906), 
	.B1(n9940), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6318));
   INVX1 U6915 (.Y(n9940), 
	.A(\ram[82][12] ));
   OAI22X1 U6916 (.Y(n1905), 
	.B1(n9941), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6320));
   INVX1 U6917 (.Y(n9941), 
	.A(\ram[82][11] ));
   OAI22X1 U6918 (.Y(n1904), 
	.B1(n9942), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6322));
   INVX1 U6919 (.Y(n9942), 
	.A(\ram[82][10] ));
   OAI22X1 U6920 (.Y(n1903), 
	.B1(n9943), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6324));
   INVX1 U6921 (.Y(n9943), 
	.A(\ram[82][9] ));
   OAI22X1 U6922 (.Y(n1902), 
	.B1(n9944), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6326));
   INVX1 U6923 (.Y(n9944), 
	.A(\ram[82][8] ));
   OAI22X1 U6924 (.Y(n1901), 
	.B1(n9945), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6328));
   INVX1 U6925 (.Y(n9945), 
	.A(\ram[82][7] ));
   OAI22X1 U6926 (.Y(n1900), 
	.B1(n9946), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6330));
   INVX1 U6927 (.Y(n9946), 
	.A(\ram[82][6] ));
   OAI22X1 U6928 (.Y(n1899), 
	.B1(n9947), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6332));
   INVX1 U6929 (.Y(n9947), 
	.A(\ram[82][5] ));
   OAI22X1 U6930 (.Y(n1898), 
	.B1(n9948), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6334));
   INVX1 U6931 (.Y(n9948), 
	.A(\ram[82][4] ));
   OAI22X1 U6932 (.Y(n1897), 
	.B1(n9949), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6336));
   INVX1 U6933 (.Y(n9949), 
	.A(\ram[82][3] ));
   OAI22X1 U6934 (.Y(n1896), 
	.B1(n9950), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6338));
   INVX1 U6935 (.Y(n9950), 
	.A(\ram[82][2] ));
   OAI22X1 U6936 (.Y(n1895), 
	.B1(n9951), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6306));
   INVX1 U6937 (.Y(n9951), 
	.A(\ram[82][1] ));
   OAI22X1 U6938 (.Y(n1894), 
	.B1(n9952), 
	.B0(n9936), 
	.A1(n9935), 
	.A0(n6309));
   INVX1 U6939 (.Y(n9952), 
	.A(\ram[82][0] ));
   NOR2BX1 U6940 (.Y(n9936), 
	.B(n9935), 
	.AN(mem_write_en));
   NAND2X1 U6941 (.Y(n9935), 
	.B(n6476), 
	.A(n9718));
   OAI22X1 U6942 (.Y(n1893), 
	.B1(n9955), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6311));
   INVX1 U6943 (.Y(n9955), 
	.A(\ram[81][15] ));
   OAI22X1 U6944 (.Y(n1892), 
	.B1(n9956), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6314));
   INVX1 U6945 (.Y(n9956), 
	.A(\ram[81][14] ));
   OAI22X1 U6946 (.Y(n1891), 
	.B1(n9957), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6316));
   INVX1 U6947 (.Y(n9957), 
	.A(\ram[81][13] ));
   OAI22X1 U6948 (.Y(n1890), 
	.B1(n9958), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6318));
   INVX1 U6949 (.Y(n9958), 
	.A(\ram[81][12] ));
   OAI22X1 U6950 (.Y(n1889), 
	.B1(n9959), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6320));
   INVX1 U6951 (.Y(n9959), 
	.A(\ram[81][11] ));
   OAI22X1 U6952 (.Y(n1888), 
	.B1(n9960), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6322));
   INVX1 U6953 (.Y(n9960), 
	.A(\ram[81][10] ));
   OAI22X1 U6954 (.Y(n1887), 
	.B1(n9961), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6324));
   INVX1 U6955 (.Y(n9961), 
	.A(\ram[81][9] ));
   OAI22X1 U6956 (.Y(n1886), 
	.B1(n9962), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6326));
   INVX1 U6957 (.Y(n9962), 
	.A(\ram[81][8] ));
   OAI22X1 U6958 (.Y(n1885), 
	.B1(n9963), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6328));
   INVX1 U6959 (.Y(n9963), 
	.A(\ram[81][7] ));
   OAI22X1 U6960 (.Y(n1884), 
	.B1(n9964), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6330));
   INVX1 U6961 (.Y(n9964), 
	.A(\ram[81][6] ));
   OAI22X1 U6962 (.Y(n1883), 
	.B1(n9965), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6332));
   INVX1 U6963 (.Y(n9965), 
	.A(\ram[81][5] ));
   OAI22X1 U6964 (.Y(n1882), 
	.B1(n9966), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6334));
   INVX1 U6965 (.Y(n9966), 
	.A(\ram[81][4] ));
   OAI22X1 U6966 (.Y(n1881), 
	.B1(n9967), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6336));
   INVX1 U6967 (.Y(n9967), 
	.A(\ram[81][3] ));
   OAI22X1 U6968 (.Y(n1880), 
	.B1(n9968), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6338));
   INVX1 U6969 (.Y(n9968), 
	.A(\ram[81][2] ));
   OAI22X1 U6970 (.Y(n1879), 
	.B1(n9969), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6306));
   INVX1 U6971 (.Y(n9969), 
	.A(\ram[81][1] ));
   OAI22X1 U6972 (.Y(n1878), 
	.B1(n9970), 
	.B0(n9954), 
	.A1(n9953), 
	.A0(n6309));
   INVX1 U6973 (.Y(n9970), 
	.A(\ram[81][0] ));
   NOR2BX1 U6974 (.Y(n9954), 
	.B(n9953), 
	.AN(mem_write_en));
   NAND2X1 U6975 (.Y(n9953), 
	.B(n6495), 
	.A(n9718));
   OAI22X1 U6976 (.Y(n1877), 
	.B1(n9973), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6311));
   INVX1 U6977 (.Y(n9973), 
	.A(\ram[80][15] ));
   OAI22X1 U6978 (.Y(n1876), 
	.B1(n9974), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6314));
   INVX1 U6979 (.Y(n9974), 
	.A(\ram[80][14] ));
   OAI22X1 U6980 (.Y(n1875), 
	.B1(n9975), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6316));
   INVX1 U6981 (.Y(n9975), 
	.A(\ram[80][13] ));
   OAI22X1 U6982 (.Y(n1874), 
	.B1(n9976), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6318));
   INVX1 U6983 (.Y(n9976), 
	.A(\ram[80][12] ));
   OAI22X1 U6984 (.Y(n1873), 
	.B1(n9977), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6320));
   INVX1 U6985 (.Y(n9977), 
	.A(\ram[80][11] ));
   OAI22X1 U6986 (.Y(n1872), 
	.B1(n9978), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6322));
   INVX1 U6987 (.Y(n9978), 
	.A(\ram[80][10] ));
   OAI22X1 U6988 (.Y(n1871), 
	.B1(n9979), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6324));
   INVX1 U6989 (.Y(n9979), 
	.A(\ram[80][9] ));
   OAI22X1 U6990 (.Y(n1870), 
	.B1(n9980), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6326));
   INVX1 U6991 (.Y(n9980), 
	.A(\ram[80][8] ));
   OAI22X1 U6992 (.Y(n1869), 
	.B1(n9981), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6328));
   INVX1 U6993 (.Y(n9981), 
	.A(\ram[80][7] ));
   OAI22X1 U6994 (.Y(n1868), 
	.B1(n9982), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6330));
   INVX1 U6995 (.Y(n9982), 
	.A(\ram[80][6] ));
   OAI22X1 U6996 (.Y(n1867), 
	.B1(n9983), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6332));
   INVX1 U6997 (.Y(n9983), 
	.A(\ram[80][5] ));
   OAI22X1 U6998 (.Y(n1866), 
	.B1(n9984), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6334));
   INVX1 U6999 (.Y(n9984), 
	.A(\ram[80][4] ));
   OAI22X1 U7000 (.Y(n1865), 
	.B1(n9985), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6336));
   INVX1 U7001 (.Y(n9985), 
	.A(\ram[80][3] ));
   OAI22X1 U7002 (.Y(n1864), 
	.B1(n9986), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6338));
   INVX1 U7003 (.Y(n9986), 
	.A(\ram[80][2] ));
   OAI22X1 U7004 (.Y(n1863), 
	.B1(n9987), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6306));
   INVX1 U7005 (.Y(n9987), 
	.A(\ram[80][1] ));
   OAI22X1 U7006 (.Y(n1862), 
	.B1(n9988), 
	.B0(n9972), 
	.A1(n9971), 
	.A0(n6309));
   INVX1 U7007 (.Y(n9988), 
	.A(\ram[80][0] ));
   NOR2BX1 U7008 (.Y(n9972), 
	.B(n9971), 
	.AN(mem_write_en));
   NAND2X1 U7009 (.Y(n9971), 
	.B(n6514), 
	.A(n9718));
   OAI22X1 U7010 (.Y(n1861), 
	.B1(n9991), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6311));
   INVX1 U7011 (.Y(n9991), 
	.A(\ram[79][15] ));
   OAI22X1 U7012 (.Y(n1860), 
	.B1(n9992), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6314));
   INVX1 U7013 (.Y(n9992), 
	.A(\ram[79][14] ));
   OAI22X1 U7014 (.Y(n1859), 
	.B1(n9993), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6316));
   INVX1 U7015 (.Y(n9993), 
	.A(\ram[79][13] ));
   OAI22X1 U7016 (.Y(n1858), 
	.B1(n9994), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6318));
   INVX1 U7017 (.Y(n9994), 
	.A(\ram[79][12] ));
   OAI22X1 U7018 (.Y(n1857), 
	.B1(n9995), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6320));
   INVX1 U7019 (.Y(n9995), 
	.A(\ram[79][11] ));
   OAI22X1 U7020 (.Y(n1856), 
	.B1(n9996), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6322));
   INVX1 U7021 (.Y(n9996), 
	.A(\ram[79][10] ));
   OAI22X1 U7022 (.Y(n1855), 
	.B1(n9997), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6324));
   INVX1 U7023 (.Y(n9997), 
	.A(\ram[79][9] ));
   OAI22X1 U7024 (.Y(n1854), 
	.B1(n9998), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6326));
   INVX1 U7025 (.Y(n9998), 
	.A(\ram[79][8] ));
   OAI22X1 U7026 (.Y(n1853), 
	.B1(n9999), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6328));
   INVX1 U7027 (.Y(n9999), 
	.A(\ram[79][7] ));
   OAI22X1 U7028 (.Y(n1852), 
	.B1(n10000), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6330));
   INVX1 U7029 (.Y(n10000), 
	.A(\ram[79][6] ));
   OAI22X1 U7030 (.Y(n1851), 
	.B1(n10001), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6332));
   INVX1 U7031 (.Y(n10001), 
	.A(\ram[79][5] ));
   OAI22X1 U7032 (.Y(n1850), 
	.B1(n10002), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6334));
   INVX1 U7033 (.Y(n10002), 
	.A(\ram[79][4] ));
   OAI22X1 U7034 (.Y(n1849), 
	.B1(n10003), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6336));
   INVX1 U7035 (.Y(n10003), 
	.A(\ram[79][3] ));
   OAI22X1 U7036 (.Y(n1848), 
	.B1(n10004), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6338));
   INVX1 U7037 (.Y(n10004), 
	.A(\ram[79][2] ));
   OAI22X1 U7038 (.Y(n1847), 
	.B1(n10005), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6306));
   INVX1 U7039 (.Y(n10005), 
	.A(\ram[79][1] ));
   OAI22X1 U7040 (.Y(n1846), 
	.B1(n10006), 
	.B0(n9990), 
	.A1(n9989), 
	.A0(n6309));
   INVX1 U7041 (.Y(n10006), 
	.A(\ram[79][0] ));
   NOR2BX1 U7042 (.Y(n9990), 
	.B(n9989), 
	.AN(mem_write_en));
   NAND2X1 U7043 (.Y(n9989), 
	.B(n6533), 
	.A(n10007));
   OAI22X1 U7044 (.Y(n1845), 
	.B1(n10010), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6311));
   INVX1 U7045 (.Y(n10010), 
	.A(\ram[78][15] ));
   OAI22X1 U7046 (.Y(n1844), 
	.B1(n10011), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6314));
   INVX1 U7047 (.Y(n10011), 
	.A(\ram[78][14] ));
   OAI22X1 U7048 (.Y(n1843), 
	.B1(n10012), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6316));
   INVX1 U7049 (.Y(n10012), 
	.A(\ram[78][13] ));
   OAI22X1 U7050 (.Y(n1842), 
	.B1(n10013), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6318));
   INVX1 U7051 (.Y(n10013), 
	.A(\ram[78][12] ));
   OAI22X1 U7052 (.Y(n1841), 
	.B1(n10014), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6320));
   INVX1 U7053 (.Y(n10014), 
	.A(\ram[78][11] ));
   OAI22X1 U7054 (.Y(n1840), 
	.B1(n10015), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6322));
   INVX1 U7055 (.Y(n10015), 
	.A(\ram[78][10] ));
   OAI22X1 U7056 (.Y(n1839), 
	.B1(n10016), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6324));
   INVX1 U7057 (.Y(n10016), 
	.A(\ram[78][9] ));
   OAI22X1 U7058 (.Y(n1838), 
	.B1(n10017), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6326));
   INVX1 U7059 (.Y(n10017), 
	.A(\ram[78][8] ));
   OAI22X1 U7060 (.Y(n1837), 
	.B1(n10018), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6328));
   INVX1 U7061 (.Y(n10018), 
	.A(\ram[78][7] ));
   OAI22X1 U7062 (.Y(n1836), 
	.B1(n10019), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6330));
   INVX1 U7063 (.Y(n10019), 
	.A(\ram[78][6] ));
   OAI22X1 U7064 (.Y(n1835), 
	.B1(n10020), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6332));
   INVX1 U7065 (.Y(n10020), 
	.A(\ram[78][5] ));
   OAI22X1 U7066 (.Y(n1834), 
	.B1(n10021), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6334));
   INVX1 U7067 (.Y(n10021), 
	.A(\ram[78][4] ));
   OAI22X1 U7068 (.Y(n1833), 
	.B1(n10022), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6336));
   INVX1 U7069 (.Y(n10022), 
	.A(\ram[78][3] ));
   OAI22X1 U7070 (.Y(n1832), 
	.B1(n10023), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6338));
   INVX1 U7071 (.Y(n10023), 
	.A(\ram[78][2] ));
   OAI22X1 U7072 (.Y(n1831), 
	.B1(n10024), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6306));
   INVX1 U7073 (.Y(n10024), 
	.A(\ram[78][1] ));
   OAI22X1 U7074 (.Y(n1830), 
	.B1(n10025), 
	.B0(n10009), 
	.A1(n10008), 
	.A0(n6309));
   INVX1 U7075 (.Y(n10025), 
	.A(\ram[78][0] ));
   NOR2BX1 U7076 (.Y(n10009), 
	.B(n10008), 
	.AN(mem_write_en));
   NAND2X1 U7077 (.Y(n10008), 
	.B(n6553), 
	.A(n10007));
   OAI22X1 U7078 (.Y(n1829), 
	.B1(n10028), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6311));
   INVX1 U7079 (.Y(n10028), 
	.A(\ram[77][15] ));
   OAI22X1 U7080 (.Y(n1828), 
	.B1(n10029), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6314));
   INVX1 U7081 (.Y(n10029), 
	.A(\ram[77][14] ));
   OAI22X1 U7082 (.Y(n1827), 
	.B1(n10030), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6316));
   INVX1 U7083 (.Y(n10030), 
	.A(\ram[77][13] ));
   OAI22X1 U7084 (.Y(n1826), 
	.B1(n10031), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6318));
   INVX1 U7085 (.Y(n10031), 
	.A(\ram[77][12] ));
   OAI22X1 U7086 (.Y(n1825), 
	.B1(n10032), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6320));
   INVX1 U7087 (.Y(n10032), 
	.A(\ram[77][11] ));
   OAI22X1 U7088 (.Y(n1824), 
	.B1(n10033), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6322));
   INVX1 U7089 (.Y(n10033), 
	.A(\ram[77][10] ));
   OAI22X1 U7090 (.Y(n1823), 
	.B1(n10034), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6324));
   INVX1 U7091 (.Y(n10034), 
	.A(\ram[77][9] ));
   OAI22X1 U7092 (.Y(n1822), 
	.B1(n10035), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6326));
   INVX1 U7093 (.Y(n10035), 
	.A(\ram[77][8] ));
   OAI22X1 U7094 (.Y(n1821), 
	.B1(n10036), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6328));
   INVX1 U7095 (.Y(n10036), 
	.A(\ram[77][7] ));
   OAI22X1 U7096 (.Y(n1820), 
	.B1(n10037), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6330));
   INVX1 U7097 (.Y(n10037), 
	.A(\ram[77][6] ));
   OAI22X1 U7098 (.Y(n1819), 
	.B1(n10038), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6332));
   INVX1 U7099 (.Y(n10038), 
	.A(\ram[77][5] ));
   OAI22X1 U7100 (.Y(n1818), 
	.B1(n10039), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6334));
   INVX1 U7101 (.Y(n10039), 
	.A(\ram[77][4] ));
   OAI22X1 U7102 (.Y(n1817), 
	.B1(n10040), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6336));
   INVX1 U7103 (.Y(n10040), 
	.A(\ram[77][3] ));
   OAI22X1 U7104 (.Y(n1816), 
	.B1(n10041), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6338));
   INVX1 U7105 (.Y(n10041), 
	.A(\ram[77][2] ));
   OAI22X1 U7106 (.Y(n1815), 
	.B1(n10042), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6306));
   INVX1 U7107 (.Y(n10042), 
	.A(\ram[77][1] ));
   OAI22X1 U7108 (.Y(n1814), 
	.B1(n10043), 
	.B0(n10027), 
	.A1(n10026), 
	.A0(n6309));
   INVX1 U7109 (.Y(n10043), 
	.A(\ram[77][0] ));
   NOR2BX1 U7110 (.Y(n10027), 
	.B(n10026), 
	.AN(mem_write_en));
   NAND2X1 U7111 (.Y(n10026), 
	.B(n6572), 
	.A(n10007));
   OAI22X1 U7112 (.Y(n1813), 
	.B1(n10046), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6311));
   INVX1 U7113 (.Y(n10046), 
	.A(\ram[76][15] ));
   OAI22X1 U7114 (.Y(n1812), 
	.B1(n10047), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6314));
   INVX1 U7115 (.Y(n10047), 
	.A(\ram[76][14] ));
   OAI22X1 U7116 (.Y(n1811), 
	.B1(n10048), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6316));
   INVX1 U7117 (.Y(n10048), 
	.A(\ram[76][13] ));
   OAI22X1 U7118 (.Y(n1810), 
	.B1(n10049), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6318));
   INVX1 U7119 (.Y(n10049), 
	.A(\ram[76][12] ));
   OAI22X1 U7120 (.Y(n1809), 
	.B1(n10050), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6320));
   INVX1 U7121 (.Y(n10050), 
	.A(\ram[76][11] ));
   OAI22X1 U7122 (.Y(n1808), 
	.B1(n10051), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6322));
   INVX1 U7123 (.Y(n10051), 
	.A(\ram[76][10] ));
   OAI22X1 U7124 (.Y(n1807), 
	.B1(n10052), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6324));
   INVX1 U7125 (.Y(n10052), 
	.A(\ram[76][9] ));
   OAI22X1 U7126 (.Y(n1806), 
	.B1(n10053), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6326));
   INVX1 U7127 (.Y(n10053), 
	.A(\ram[76][8] ));
   OAI22X1 U7128 (.Y(n1805), 
	.B1(n10054), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6328));
   INVX1 U7129 (.Y(n10054), 
	.A(\ram[76][7] ));
   OAI22X1 U7130 (.Y(n1804), 
	.B1(n10055), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6330));
   INVX1 U7131 (.Y(n10055), 
	.A(\ram[76][6] ));
   OAI22X1 U7132 (.Y(n1803), 
	.B1(n10056), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6332));
   INVX1 U7133 (.Y(n10056), 
	.A(\ram[76][5] ));
   OAI22X1 U7134 (.Y(n1802), 
	.B1(n10057), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6334));
   INVX1 U7135 (.Y(n10057), 
	.A(\ram[76][4] ));
   OAI22X1 U7136 (.Y(n1801), 
	.B1(n10058), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6336));
   INVX1 U7137 (.Y(n10058), 
	.A(\ram[76][3] ));
   OAI22X1 U7138 (.Y(n1800), 
	.B1(n10059), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6338));
   INVX1 U7139 (.Y(n10059), 
	.A(\ram[76][2] ));
   OAI22X1 U7140 (.Y(n1799), 
	.B1(n10060), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6306));
   INVX1 U7141 (.Y(n10060), 
	.A(\ram[76][1] ));
   OAI22X1 U7142 (.Y(n1798), 
	.B1(n10061), 
	.B0(n10045), 
	.A1(n10044), 
	.A0(n6309));
   INVX1 U7143 (.Y(n10061), 
	.A(\ram[76][0] ));
   NOR2BX1 U7144 (.Y(n10045), 
	.B(n10044), 
	.AN(mem_write_en));
   NAND2X1 U7145 (.Y(n10044), 
	.B(n6591), 
	.A(n10007));
   OAI22X1 U7146 (.Y(n1797), 
	.B1(n10064), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6311));
   INVX1 U7147 (.Y(n10064), 
	.A(\ram[75][15] ));
   OAI22X1 U7148 (.Y(n1796), 
	.B1(n10065), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6314));
   INVX1 U7149 (.Y(n10065), 
	.A(\ram[75][14] ));
   OAI22X1 U7150 (.Y(n1795), 
	.B1(n10066), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6316));
   INVX1 U7151 (.Y(n10066), 
	.A(\ram[75][13] ));
   OAI22X1 U7152 (.Y(n1794), 
	.B1(n10067), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6318));
   INVX1 U7153 (.Y(n10067), 
	.A(\ram[75][12] ));
   OAI22X1 U7154 (.Y(n1793), 
	.B1(n10068), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6320));
   INVX1 U7155 (.Y(n10068), 
	.A(\ram[75][11] ));
   OAI22X1 U7156 (.Y(n1792), 
	.B1(n10069), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6322));
   INVX1 U7157 (.Y(n10069), 
	.A(\ram[75][10] ));
   OAI22X1 U7158 (.Y(n1791), 
	.B1(n10070), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6324));
   INVX1 U7159 (.Y(n10070), 
	.A(\ram[75][9] ));
   OAI22X1 U7160 (.Y(n1790), 
	.B1(n10071), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6326));
   INVX1 U7161 (.Y(n10071), 
	.A(\ram[75][8] ));
   OAI22X1 U7162 (.Y(n1789), 
	.B1(n10072), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6328));
   INVX1 U7163 (.Y(n10072), 
	.A(\ram[75][7] ));
   OAI22X1 U7164 (.Y(n1788), 
	.B1(n10073), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6330));
   INVX1 U7165 (.Y(n10073), 
	.A(\ram[75][6] ));
   OAI22X1 U7166 (.Y(n1787), 
	.B1(n10074), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6332));
   INVX1 U7167 (.Y(n10074), 
	.A(\ram[75][5] ));
   OAI22X1 U7168 (.Y(n1786), 
	.B1(n10075), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6334));
   INVX1 U7169 (.Y(n10075), 
	.A(\ram[75][4] ));
   OAI22X1 U7170 (.Y(n1785), 
	.B1(n10076), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6336));
   INVX1 U7171 (.Y(n10076), 
	.A(\ram[75][3] ));
   OAI22X1 U7172 (.Y(n1784), 
	.B1(n10077), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6338));
   INVX1 U7173 (.Y(n10077), 
	.A(\ram[75][2] ));
   OAI22X1 U7174 (.Y(n1783), 
	.B1(n10078), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6306));
   INVX1 U7175 (.Y(n10078), 
	.A(\ram[75][1] ));
   OAI22X1 U7176 (.Y(n1782), 
	.B1(n10079), 
	.B0(n10063), 
	.A1(n10062), 
	.A0(n6309));
   INVX1 U7177 (.Y(n10079), 
	.A(\ram[75][0] ));
   NOR2BX1 U7178 (.Y(n10063), 
	.B(n10062), 
	.AN(mem_write_en));
   NAND2X1 U7179 (.Y(n10062), 
	.B(n6610), 
	.A(n10007));
   OAI22X1 U7180 (.Y(n1781), 
	.B1(n10082), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6311));
   INVX1 U7181 (.Y(n10082), 
	.A(\ram[74][15] ));
   OAI22X1 U7182 (.Y(n1780), 
	.B1(n10083), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6314));
   INVX1 U7183 (.Y(n10083), 
	.A(\ram[74][14] ));
   OAI22X1 U7184 (.Y(n1779), 
	.B1(n10084), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6316));
   INVX1 U7185 (.Y(n10084), 
	.A(\ram[74][13] ));
   OAI22X1 U7186 (.Y(n1778), 
	.B1(n10085), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6318));
   INVX1 U7187 (.Y(n10085), 
	.A(\ram[74][12] ));
   OAI22X1 U7188 (.Y(n1777), 
	.B1(n10086), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6320));
   INVX1 U7189 (.Y(n10086), 
	.A(\ram[74][11] ));
   OAI22X1 U7190 (.Y(n1776), 
	.B1(n10087), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6322));
   INVX1 U7191 (.Y(n10087), 
	.A(\ram[74][10] ));
   OAI22X1 U7192 (.Y(n1775), 
	.B1(n10088), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6324));
   INVX1 U7193 (.Y(n10088), 
	.A(\ram[74][9] ));
   OAI22X1 U7194 (.Y(n1774), 
	.B1(n10089), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6326));
   INVX1 U7195 (.Y(n10089), 
	.A(\ram[74][8] ));
   OAI22X1 U7196 (.Y(n1773), 
	.B1(n10090), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6328));
   INVX1 U7197 (.Y(n10090), 
	.A(\ram[74][7] ));
   OAI22X1 U7198 (.Y(n1772), 
	.B1(n10091), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6330));
   INVX1 U7199 (.Y(n10091), 
	.A(\ram[74][6] ));
   OAI22X1 U7200 (.Y(n1771), 
	.B1(n10092), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6332));
   INVX1 U7201 (.Y(n10092), 
	.A(\ram[74][5] ));
   OAI22X1 U7202 (.Y(n1770), 
	.B1(n10093), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6334));
   INVX1 U7203 (.Y(n10093), 
	.A(\ram[74][4] ));
   OAI22X1 U7204 (.Y(n1769), 
	.B1(n10094), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6336));
   INVX1 U7205 (.Y(n10094), 
	.A(\ram[74][3] ));
   OAI22X1 U7206 (.Y(n1768), 
	.B1(n10095), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6338));
   INVX1 U7207 (.Y(n10095), 
	.A(\ram[74][2] ));
   OAI22X1 U7208 (.Y(n1767), 
	.B1(n10096), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6306));
   INVX1 U7209 (.Y(n10096), 
	.A(\ram[74][1] ));
   OAI22X1 U7210 (.Y(n1766), 
	.B1(n10097), 
	.B0(n10081), 
	.A1(n10080), 
	.A0(n6309));
   INVX1 U7211 (.Y(n10097), 
	.A(\ram[74][0] ));
   NOR2BX1 U7212 (.Y(n10081), 
	.B(n10080), 
	.AN(mem_write_en));
   NAND2X1 U7213 (.Y(n10080), 
	.B(n6629), 
	.A(n10007));
   OAI22X1 U7214 (.Y(n1765), 
	.B1(n10100), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6311));
   INVX1 U7215 (.Y(n10100), 
	.A(\ram[73][15] ));
   OAI22X1 U7216 (.Y(n1764), 
	.B1(n10101), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6314));
   INVX1 U7217 (.Y(n10101), 
	.A(\ram[73][14] ));
   OAI22X1 U7218 (.Y(n1763), 
	.B1(n10102), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6316));
   INVX1 U7219 (.Y(n10102), 
	.A(\ram[73][13] ));
   OAI22X1 U7220 (.Y(n1762), 
	.B1(n10103), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6318));
   INVX1 U7221 (.Y(n10103), 
	.A(\ram[73][12] ));
   OAI22X1 U7222 (.Y(n1761), 
	.B1(n10104), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6320));
   INVX1 U7223 (.Y(n10104), 
	.A(\ram[73][11] ));
   OAI22X1 U7224 (.Y(n1760), 
	.B1(n10105), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6322));
   INVX1 U7225 (.Y(n10105), 
	.A(\ram[73][10] ));
   OAI22X1 U7226 (.Y(n1759), 
	.B1(n10106), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6324));
   INVX1 U7227 (.Y(n10106), 
	.A(\ram[73][9] ));
   OAI22X1 U7228 (.Y(n1758), 
	.B1(n10107), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6326));
   INVX1 U7229 (.Y(n10107), 
	.A(\ram[73][8] ));
   OAI22X1 U7230 (.Y(n1757), 
	.B1(n10108), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6328));
   INVX1 U7231 (.Y(n10108), 
	.A(\ram[73][7] ));
   OAI22X1 U7232 (.Y(n1756), 
	.B1(n10109), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6330));
   INVX1 U7233 (.Y(n10109), 
	.A(\ram[73][6] ));
   OAI22X1 U7234 (.Y(n1755), 
	.B1(n10110), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6332));
   INVX1 U7235 (.Y(n10110), 
	.A(\ram[73][5] ));
   OAI22X1 U7236 (.Y(n1754), 
	.B1(n10111), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6334));
   INVX1 U7237 (.Y(n10111), 
	.A(\ram[73][4] ));
   OAI22X1 U7238 (.Y(n1753), 
	.B1(n10112), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6336));
   INVX1 U7239 (.Y(n10112), 
	.A(\ram[73][3] ));
   OAI22X1 U7240 (.Y(n1752), 
	.B1(n10113), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6338));
   INVX1 U7241 (.Y(n10113), 
	.A(\ram[73][2] ));
   OAI22X1 U7242 (.Y(n1751), 
	.B1(n10114), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6306));
   INVX1 U7243 (.Y(n10114), 
	.A(\ram[73][1] ));
   OAI22X1 U7244 (.Y(n1750), 
	.B1(n10115), 
	.B0(n10099), 
	.A1(n10098), 
	.A0(n6309));
   INVX1 U7245 (.Y(n10115), 
	.A(\ram[73][0] ));
   NOR2BX1 U7246 (.Y(n10099), 
	.B(n10098), 
	.AN(mem_write_en));
   NAND2X1 U7247 (.Y(n10098), 
	.B(n6342), 
	.A(n10007));
   OAI22X1 U7248 (.Y(n1749), 
	.B1(n10118), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6311));
   INVX1 U7249 (.Y(n10118), 
	.A(\ram[72][15] ));
   OAI22X1 U7250 (.Y(n1748), 
	.B1(n10119), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6314));
   INVX1 U7251 (.Y(n10119), 
	.A(\ram[72][14] ));
   OAI22X1 U7252 (.Y(n1747), 
	.B1(n10120), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6316));
   INVX1 U7253 (.Y(n10120), 
	.A(\ram[72][13] ));
   OAI22X1 U7254 (.Y(n1746), 
	.B1(n10121), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6318));
   INVX1 U7255 (.Y(n10121), 
	.A(\ram[72][12] ));
   OAI22X1 U7256 (.Y(n1745), 
	.B1(n10122), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6320));
   INVX1 U7257 (.Y(n10122), 
	.A(\ram[72][11] ));
   OAI22X1 U7258 (.Y(n1744), 
	.B1(n10123), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6322));
   INVX1 U7259 (.Y(n10123), 
	.A(\ram[72][10] ));
   OAI22X1 U7260 (.Y(n1743), 
	.B1(n10124), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6324));
   INVX1 U7261 (.Y(n10124), 
	.A(\ram[72][9] ));
   OAI22X1 U7262 (.Y(n1742), 
	.B1(n10125), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6326));
   INVX1 U7263 (.Y(n10125), 
	.A(\ram[72][8] ));
   OAI22X1 U7264 (.Y(n1741), 
	.B1(n10126), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6328));
   INVX1 U7265 (.Y(n10126), 
	.A(\ram[72][7] ));
   OAI22X1 U7266 (.Y(n1740), 
	.B1(n10127), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6330));
   INVX1 U7267 (.Y(n10127), 
	.A(\ram[72][6] ));
   OAI22X1 U7268 (.Y(n1739), 
	.B1(n10128), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6332));
   INVX1 U7269 (.Y(n10128), 
	.A(\ram[72][5] ));
   OAI22X1 U7270 (.Y(n1738), 
	.B1(n10129), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6334));
   INVX1 U7271 (.Y(n10129), 
	.A(\ram[72][4] ));
   OAI22X1 U7272 (.Y(n1737), 
	.B1(n10130), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6336));
   INVX1 U7273 (.Y(n10130), 
	.A(\ram[72][3] ));
   OAI22X1 U7274 (.Y(n1736), 
	.B1(n10131), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6338));
   INVX1 U7275 (.Y(n10131), 
	.A(\ram[72][2] ));
   OAI22X1 U7276 (.Y(n1735), 
	.B1(n10132), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6306));
   INVX1 U7277 (.Y(n10132), 
	.A(\ram[72][1] ));
   OAI22X1 U7278 (.Y(n1734), 
	.B1(n10133), 
	.B0(n10117), 
	.A1(n10116), 
	.A0(n6309));
   INVX1 U7279 (.Y(n10133), 
	.A(\ram[72][0] ));
   NOR2BX1 U7280 (.Y(n10117), 
	.B(n10116), 
	.AN(mem_write_en));
   NAND2X1 U7281 (.Y(n10116), 
	.B(n6362), 
	.A(n10007));
   OAI22X1 U7282 (.Y(n1733), 
	.B1(n10136), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6311));
   INVX1 U7283 (.Y(n10136), 
	.A(\ram[71][15] ));
   OAI22X1 U7284 (.Y(n1732), 
	.B1(n10137), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6314));
   INVX1 U7285 (.Y(n10137), 
	.A(\ram[71][14] ));
   OAI22X1 U7286 (.Y(n1731), 
	.B1(n10138), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6316));
   INVX1 U7287 (.Y(n10138), 
	.A(\ram[71][13] ));
   OAI22X1 U7288 (.Y(n1730), 
	.B1(n10139), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6318));
   INVX1 U7289 (.Y(n10139), 
	.A(\ram[71][12] ));
   OAI22X1 U7290 (.Y(n1729), 
	.B1(n10140), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6320));
   INVX1 U7291 (.Y(n10140), 
	.A(\ram[71][11] ));
   OAI22X1 U7292 (.Y(n1728), 
	.B1(n10141), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6322));
   INVX1 U7293 (.Y(n10141), 
	.A(\ram[71][10] ));
   OAI22X1 U7294 (.Y(n1727), 
	.B1(n10142), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6324));
   INVX1 U7295 (.Y(n10142), 
	.A(\ram[71][9] ));
   OAI22X1 U7296 (.Y(n1726), 
	.B1(n10143), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6326));
   INVX1 U7297 (.Y(n10143), 
	.A(\ram[71][8] ));
   OAI22X1 U7298 (.Y(n1725), 
	.B1(n10144), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6328));
   INVX1 U7299 (.Y(n10144), 
	.A(\ram[71][7] ));
   OAI22X1 U7300 (.Y(n1724), 
	.B1(n10145), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6330));
   INVX1 U7301 (.Y(n10145), 
	.A(\ram[71][6] ));
   OAI22X1 U7302 (.Y(n1723), 
	.B1(n10146), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6332));
   INVX1 U7303 (.Y(n10146), 
	.A(\ram[71][5] ));
   OAI22X1 U7304 (.Y(n1722), 
	.B1(n10147), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6334));
   INVX1 U7305 (.Y(n10147), 
	.A(\ram[71][4] ));
   OAI22X1 U7306 (.Y(n1721), 
	.B1(n10148), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6336));
   INVX1 U7307 (.Y(n10148), 
	.A(\ram[71][3] ));
   OAI22X1 U7308 (.Y(n1720), 
	.B1(n10149), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6338));
   INVX1 U7309 (.Y(n10149), 
	.A(\ram[71][2] ));
   OAI22X1 U7310 (.Y(n1719), 
	.B1(n10150), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6306));
   INVX1 U7311 (.Y(n10150), 
	.A(\ram[71][1] ));
   OAI22X1 U7312 (.Y(n1718), 
	.B1(n10151), 
	.B0(n10135), 
	.A1(n10134), 
	.A0(n6309));
   INVX1 U7313 (.Y(n10151), 
	.A(\ram[71][0] ));
   NOR2BX1 U7314 (.Y(n10135), 
	.B(n10134), 
	.AN(mem_write_en));
   NAND2X1 U7315 (.Y(n10134), 
	.B(n6381), 
	.A(n10007));
   OAI22X1 U7316 (.Y(n1717), 
	.B1(n10154), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6311));
   INVX1 U7317 (.Y(n10154), 
	.A(\ram[70][15] ));
   OAI22X1 U7318 (.Y(n1716), 
	.B1(n10155), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6314));
   INVX1 U7319 (.Y(n10155), 
	.A(\ram[70][14] ));
   OAI22X1 U7320 (.Y(n1715), 
	.B1(n10156), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6316));
   INVX1 U7321 (.Y(n10156), 
	.A(\ram[70][13] ));
   OAI22X1 U7322 (.Y(n1714), 
	.B1(n10157), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6318));
   INVX1 U7323 (.Y(n10157), 
	.A(\ram[70][12] ));
   OAI22X1 U7324 (.Y(n1713), 
	.B1(n10158), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6320));
   INVX1 U7325 (.Y(n10158), 
	.A(\ram[70][11] ));
   OAI22X1 U7326 (.Y(n1712), 
	.B1(n10159), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6322));
   INVX1 U7327 (.Y(n10159), 
	.A(\ram[70][10] ));
   OAI22X1 U7328 (.Y(n1711), 
	.B1(n10160), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6324));
   INVX1 U7329 (.Y(n10160), 
	.A(\ram[70][9] ));
   OAI22X1 U7330 (.Y(n1710), 
	.B1(n10161), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6326));
   INVX1 U7331 (.Y(n10161), 
	.A(\ram[70][8] ));
   OAI22X1 U7332 (.Y(n1709), 
	.B1(n10162), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6328));
   INVX1 U7333 (.Y(n10162), 
	.A(\ram[70][7] ));
   OAI22X1 U7334 (.Y(n1708), 
	.B1(n10163), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6330));
   INVX1 U7335 (.Y(n10163), 
	.A(\ram[70][6] ));
   OAI22X1 U7336 (.Y(n1707), 
	.B1(n10164), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6332));
   INVX1 U7337 (.Y(n10164), 
	.A(\ram[70][5] ));
   OAI22X1 U7338 (.Y(n1706), 
	.B1(n10165), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6334));
   INVX1 U7339 (.Y(n10165), 
	.A(\ram[70][4] ));
   OAI22X1 U7340 (.Y(n1705), 
	.B1(n10166), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6336));
   INVX1 U7341 (.Y(n10166), 
	.A(\ram[70][3] ));
   OAI22X1 U7342 (.Y(n1704), 
	.B1(n10167), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6338));
   INVX1 U7343 (.Y(n10167), 
	.A(\ram[70][2] ));
   OAI22X1 U7344 (.Y(n1703), 
	.B1(n10168), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6306));
   INVX1 U7345 (.Y(n10168), 
	.A(\ram[70][1] ));
   OAI22X1 U7346 (.Y(n1702), 
	.B1(n10169), 
	.B0(n10153), 
	.A1(n10152), 
	.A0(n6309));
   INVX1 U7347 (.Y(n10169), 
	.A(\ram[70][0] ));
   NOR2BX1 U7348 (.Y(n10153), 
	.B(n10152), 
	.AN(mem_write_en));
   NAND2X1 U7349 (.Y(n10152), 
	.B(n6400), 
	.A(n10007));
   OAI22X1 U7350 (.Y(n1701), 
	.B1(n10172), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6311));
   INVX1 U7351 (.Y(n10172), 
	.A(\ram[69][15] ));
   OAI22X1 U7352 (.Y(n1700), 
	.B1(n10173), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6314));
   INVX1 U7353 (.Y(n10173), 
	.A(\ram[69][14] ));
   OAI22X1 U7354 (.Y(n1699), 
	.B1(n10174), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6316));
   INVX1 U7355 (.Y(n10174), 
	.A(\ram[69][13] ));
   OAI22X1 U7356 (.Y(n1698), 
	.B1(n10175), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6318));
   INVX1 U7357 (.Y(n10175), 
	.A(\ram[69][12] ));
   OAI22X1 U7358 (.Y(n1697), 
	.B1(n10176), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6320));
   INVX1 U7359 (.Y(n10176), 
	.A(\ram[69][11] ));
   OAI22X1 U7360 (.Y(n1696), 
	.B1(n10177), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6322));
   INVX1 U7361 (.Y(n10177), 
	.A(\ram[69][10] ));
   OAI22X1 U7362 (.Y(n1695), 
	.B1(n10178), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6324));
   INVX1 U7363 (.Y(n10178), 
	.A(\ram[69][9] ));
   OAI22X1 U7364 (.Y(n1694), 
	.B1(n10179), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6326));
   INVX1 U7365 (.Y(n10179), 
	.A(\ram[69][8] ));
   OAI22X1 U7366 (.Y(n1693), 
	.B1(n10180), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6328));
   INVX1 U7367 (.Y(n10180), 
	.A(\ram[69][7] ));
   OAI22X1 U7368 (.Y(n1692), 
	.B1(n10181), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6330));
   INVX1 U7369 (.Y(n10181), 
	.A(\ram[69][6] ));
   OAI22X1 U7370 (.Y(n1691), 
	.B1(n10182), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6332));
   INVX1 U7371 (.Y(n10182), 
	.A(\ram[69][5] ));
   OAI22X1 U7372 (.Y(n1690), 
	.B1(n10183), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6334));
   INVX1 U7373 (.Y(n10183), 
	.A(\ram[69][4] ));
   OAI22X1 U7374 (.Y(n1689), 
	.B1(n10184), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6336));
   INVX1 U7375 (.Y(n10184), 
	.A(\ram[69][3] ));
   OAI22X1 U7376 (.Y(n1688), 
	.B1(n10185), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6338));
   INVX1 U7377 (.Y(n10185), 
	.A(\ram[69][2] ));
   OAI22X1 U7378 (.Y(n1687), 
	.B1(n10186), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6306));
   INVX1 U7379 (.Y(n10186), 
	.A(\ram[69][1] ));
   OAI22X1 U7380 (.Y(n1686), 
	.B1(n10187), 
	.B0(n10171), 
	.A1(n10170), 
	.A0(n6309));
   INVX1 U7381 (.Y(n10187), 
	.A(\ram[69][0] ));
   NOR2BX1 U7382 (.Y(n10171), 
	.B(n10170), 
	.AN(mem_write_en));
   NAND2X1 U7383 (.Y(n10170), 
	.B(n6419), 
	.A(n10007));
   OAI22X1 U7384 (.Y(n1685), 
	.B1(n10190), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6311));
   INVX1 U7385 (.Y(n10190), 
	.A(\ram[68][15] ));
   OAI22X1 U7386 (.Y(n1684), 
	.B1(n10191), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6314));
   INVX1 U7387 (.Y(n10191), 
	.A(\ram[68][14] ));
   OAI22X1 U7388 (.Y(n1683), 
	.B1(n10192), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6316));
   INVX1 U7389 (.Y(n10192), 
	.A(\ram[68][13] ));
   OAI22X1 U7390 (.Y(n1682), 
	.B1(n10193), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6318));
   INVX1 U7391 (.Y(n10193), 
	.A(\ram[68][12] ));
   OAI22X1 U7392 (.Y(n1681), 
	.B1(n10194), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6320));
   INVX1 U7393 (.Y(n10194), 
	.A(\ram[68][11] ));
   OAI22X1 U7394 (.Y(n1680), 
	.B1(n10195), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6322));
   INVX1 U7395 (.Y(n10195), 
	.A(\ram[68][10] ));
   OAI22X1 U7396 (.Y(n1679), 
	.B1(n10196), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6324));
   INVX1 U7397 (.Y(n10196), 
	.A(\ram[68][9] ));
   OAI22X1 U7398 (.Y(n1678), 
	.B1(n10197), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6326));
   INVX1 U7399 (.Y(n10197), 
	.A(\ram[68][8] ));
   OAI22X1 U7400 (.Y(n1677), 
	.B1(n10198), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6328));
   INVX1 U7401 (.Y(n10198), 
	.A(\ram[68][7] ));
   OAI22X1 U7402 (.Y(n1676), 
	.B1(n10199), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6330));
   INVX1 U7403 (.Y(n10199), 
	.A(\ram[68][6] ));
   OAI22X1 U7404 (.Y(n1675), 
	.B1(n10200), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6332));
   INVX1 U7405 (.Y(n10200), 
	.A(\ram[68][5] ));
   OAI22X1 U7406 (.Y(n1674), 
	.B1(n10201), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6334));
   INVX1 U7407 (.Y(n10201), 
	.A(\ram[68][4] ));
   OAI22X1 U7408 (.Y(n1673), 
	.B1(n10202), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6336));
   INVX1 U7409 (.Y(n10202), 
	.A(\ram[68][3] ));
   OAI22X1 U7410 (.Y(n1672), 
	.B1(n10203), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6338));
   INVX1 U7411 (.Y(n10203), 
	.A(\ram[68][2] ));
   OAI22X1 U7412 (.Y(n1671), 
	.B1(n10204), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6306));
   INVX1 U7413 (.Y(n10204), 
	.A(\ram[68][1] ));
   OAI22X1 U7414 (.Y(n1670), 
	.B1(n10205), 
	.B0(n10189), 
	.A1(n10188), 
	.A0(n6309));
   INVX1 U7415 (.Y(n10205), 
	.A(\ram[68][0] ));
   NOR2BX1 U7416 (.Y(n10189), 
	.B(n10188), 
	.AN(mem_write_en));
   NAND2X1 U7417 (.Y(n10188), 
	.B(n6438), 
	.A(n10007));
   OAI22X1 U7418 (.Y(n1669), 
	.B1(n10208), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6311));
   INVX1 U7419 (.Y(n10208), 
	.A(\ram[67][15] ));
   OAI22X1 U7420 (.Y(n1668), 
	.B1(n10209), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6314));
   INVX1 U7421 (.Y(n10209), 
	.A(\ram[67][14] ));
   OAI22X1 U7422 (.Y(n1667), 
	.B1(n10210), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6316));
   INVX1 U7423 (.Y(n10210), 
	.A(\ram[67][13] ));
   OAI22X1 U7424 (.Y(n1666), 
	.B1(n10211), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6318));
   INVX1 U7425 (.Y(n10211), 
	.A(\ram[67][12] ));
   OAI22X1 U7426 (.Y(n1665), 
	.B1(n10212), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6320));
   INVX1 U7427 (.Y(n10212), 
	.A(\ram[67][11] ));
   OAI22X1 U7428 (.Y(n1664), 
	.B1(n10213), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6322));
   INVX1 U7429 (.Y(n10213), 
	.A(\ram[67][10] ));
   OAI22X1 U7430 (.Y(n1663), 
	.B1(n10214), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6324));
   INVX1 U7431 (.Y(n10214), 
	.A(\ram[67][9] ));
   OAI22X1 U7432 (.Y(n1662), 
	.B1(n10215), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6326));
   INVX1 U7433 (.Y(n10215), 
	.A(\ram[67][8] ));
   OAI22X1 U7434 (.Y(n1661), 
	.B1(n10216), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6328));
   INVX1 U7435 (.Y(n10216), 
	.A(\ram[67][7] ));
   OAI22X1 U7436 (.Y(n1660), 
	.B1(n10217), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6330));
   INVX1 U7437 (.Y(n10217), 
	.A(\ram[67][6] ));
   OAI22X1 U7438 (.Y(n1659), 
	.B1(n10218), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6332));
   INVX1 U7439 (.Y(n10218), 
	.A(\ram[67][5] ));
   OAI22X1 U7440 (.Y(n1658), 
	.B1(n10219), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6334));
   INVX1 U7441 (.Y(n10219), 
	.A(\ram[67][4] ));
   OAI22X1 U7442 (.Y(n1657), 
	.B1(n10220), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6336));
   INVX1 U7443 (.Y(n10220), 
	.A(\ram[67][3] ));
   OAI22X1 U7444 (.Y(n1656), 
	.B1(n10221), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6338));
   INVX1 U7445 (.Y(n10221), 
	.A(\ram[67][2] ));
   OAI22X1 U7446 (.Y(n1655), 
	.B1(n10222), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6306));
   INVX1 U7447 (.Y(n10222), 
	.A(\ram[67][1] ));
   OAI22X1 U7448 (.Y(n1654), 
	.B1(n10223), 
	.B0(n10207), 
	.A1(n10206), 
	.A0(n6309));
   INVX1 U7449 (.Y(n10223), 
	.A(\ram[67][0] ));
   NOR2BX1 U7450 (.Y(n10207), 
	.B(n10206), 
	.AN(mem_write_en));
   NAND2X1 U7451 (.Y(n10206), 
	.B(n6457), 
	.A(n10007));
   OAI22X1 U7452 (.Y(n1653), 
	.B1(n10226), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6311));
   INVX1 U7453 (.Y(n10226), 
	.A(\ram[66][15] ));
   OAI22X1 U7454 (.Y(n1652), 
	.B1(n10227), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6314));
   INVX1 U7455 (.Y(n10227), 
	.A(\ram[66][14] ));
   OAI22X1 U7456 (.Y(n1651), 
	.B1(n10228), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6316));
   INVX1 U7457 (.Y(n10228), 
	.A(\ram[66][13] ));
   OAI22X1 U7458 (.Y(n1650), 
	.B1(n10229), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6318));
   INVX1 U7459 (.Y(n10229), 
	.A(\ram[66][12] ));
   OAI22X1 U7460 (.Y(n1649), 
	.B1(n10230), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6320));
   INVX1 U7461 (.Y(n10230), 
	.A(\ram[66][11] ));
   OAI22X1 U7462 (.Y(n1648), 
	.B1(n10231), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6322));
   INVX1 U7463 (.Y(n10231), 
	.A(\ram[66][10] ));
   OAI22X1 U7464 (.Y(n1647), 
	.B1(n10232), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6324));
   INVX1 U7465 (.Y(n10232), 
	.A(\ram[66][9] ));
   OAI22X1 U7466 (.Y(n1646), 
	.B1(n10233), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6326));
   INVX1 U7467 (.Y(n10233), 
	.A(\ram[66][8] ));
   OAI22X1 U7468 (.Y(n1645), 
	.B1(n10234), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6328));
   INVX1 U7469 (.Y(n10234), 
	.A(\ram[66][7] ));
   OAI22X1 U7470 (.Y(n1644), 
	.B1(n10235), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6330));
   INVX1 U7471 (.Y(n10235), 
	.A(\ram[66][6] ));
   OAI22X1 U7472 (.Y(n1643), 
	.B1(n10236), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6332));
   INVX1 U7473 (.Y(n10236), 
	.A(\ram[66][5] ));
   OAI22X1 U7474 (.Y(n1642), 
	.B1(n10237), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6334));
   INVX1 U7475 (.Y(n10237), 
	.A(\ram[66][4] ));
   OAI22X1 U7476 (.Y(n1641), 
	.B1(n10238), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6336));
   INVX1 U7477 (.Y(n10238), 
	.A(\ram[66][3] ));
   OAI22X1 U7478 (.Y(n1640), 
	.B1(n10239), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6338));
   INVX1 U7479 (.Y(n10239), 
	.A(\ram[66][2] ));
   OAI22X1 U7480 (.Y(n1639), 
	.B1(n10240), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6306));
   INVX1 U7481 (.Y(n10240), 
	.A(\ram[66][1] ));
   OAI22X1 U7482 (.Y(n1638), 
	.B1(n10241), 
	.B0(n10225), 
	.A1(n10224), 
	.A0(n6309));
   INVX1 U7483 (.Y(n10241), 
	.A(\ram[66][0] ));
   NOR2BX1 U7484 (.Y(n10225), 
	.B(n10224), 
	.AN(mem_write_en));
   NAND2X1 U7485 (.Y(n10224), 
	.B(n6476), 
	.A(n10007));
   OAI22X1 U7486 (.Y(n1637), 
	.B1(n10244), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6311));
   INVX1 U7487 (.Y(n10244), 
	.A(\ram[65][15] ));
   OAI22X1 U7488 (.Y(n1636), 
	.B1(n10245), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6314));
   INVX1 U7489 (.Y(n10245), 
	.A(\ram[65][14] ));
   OAI22X1 U7490 (.Y(n1635), 
	.B1(n10246), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6316));
   INVX1 U7491 (.Y(n10246), 
	.A(\ram[65][13] ));
   OAI22X1 U7492 (.Y(n1634), 
	.B1(n10247), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6318));
   INVX1 U7493 (.Y(n10247), 
	.A(\ram[65][12] ));
   OAI22X1 U7494 (.Y(n1633), 
	.B1(n10248), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6320));
   INVX1 U7495 (.Y(n10248), 
	.A(\ram[65][11] ));
   OAI22X1 U7496 (.Y(n1632), 
	.B1(n10249), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6322));
   INVX1 U7497 (.Y(n10249), 
	.A(\ram[65][10] ));
   OAI22X1 U7498 (.Y(n1631), 
	.B1(n10250), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6324));
   INVX1 U7499 (.Y(n10250), 
	.A(\ram[65][9] ));
   OAI22X1 U7500 (.Y(n1630), 
	.B1(n10251), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6326));
   INVX1 U7501 (.Y(n10251), 
	.A(\ram[65][8] ));
   OAI22X1 U7502 (.Y(n1629), 
	.B1(n10252), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6328));
   INVX1 U7503 (.Y(n10252), 
	.A(\ram[65][7] ));
   OAI22X1 U7504 (.Y(n1628), 
	.B1(n10253), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6330));
   INVX1 U7505 (.Y(n10253), 
	.A(\ram[65][6] ));
   OAI22X1 U7506 (.Y(n1627), 
	.B1(n10254), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6332));
   INVX1 U7507 (.Y(n10254), 
	.A(\ram[65][5] ));
   OAI22X1 U7508 (.Y(n1626), 
	.B1(n10255), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6334));
   INVX1 U7509 (.Y(n10255), 
	.A(\ram[65][4] ));
   OAI22X1 U7510 (.Y(n1625), 
	.B1(n10256), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6336));
   INVX1 U7511 (.Y(n10256), 
	.A(\ram[65][3] ));
   OAI22X1 U7512 (.Y(n1624), 
	.B1(n10257), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6338));
   INVX1 U7513 (.Y(n10257), 
	.A(\ram[65][2] ));
   OAI22X1 U7514 (.Y(n1623), 
	.B1(n10258), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6306));
   INVX1 U7515 (.Y(n10258), 
	.A(\ram[65][1] ));
   OAI22X1 U7516 (.Y(n1622), 
	.B1(n10259), 
	.B0(n10243), 
	.A1(n10242), 
	.A0(n6309));
   INVX1 U7517 (.Y(n10259), 
	.A(\ram[65][0] ));
   NOR2BX1 U7518 (.Y(n10243), 
	.B(n10242), 
	.AN(mem_write_en));
   NAND2X1 U7519 (.Y(n10242), 
	.B(n6495), 
	.A(n10007));
   OAI22X1 U7520 (.Y(n1621), 
	.B1(n10262), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6311));
   INVX1 U7521 (.Y(n10262), 
	.A(\ram[64][15] ));
   OAI22X1 U7522 (.Y(n1620), 
	.B1(n10263), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6314));
   INVX1 U7523 (.Y(n10263), 
	.A(\ram[64][14] ));
   OAI22X1 U7524 (.Y(n1619), 
	.B1(n10264), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6316));
   INVX1 U7525 (.Y(n10264), 
	.A(\ram[64][13] ));
   OAI22X1 U7526 (.Y(n1618), 
	.B1(n10265), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6318));
   INVX1 U7527 (.Y(n10265), 
	.A(\ram[64][12] ));
   OAI22X1 U7528 (.Y(n1617), 
	.B1(n10266), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6320));
   INVX1 U7529 (.Y(n10266), 
	.A(\ram[64][11] ));
   OAI22X1 U7530 (.Y(n1616), 
	.B1(n10267), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6322));
   INVX1 U7531 (.Y(n10267), 
	.A(\ram[64][10] ));
   OAI22X1 U7532 (.Y(n1615), 
	.B1(n10268), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6324));
   INVX1 U7533 (.Y(n10268), 
	.A(\ram[64][9] ));
   OAI22X1 U7534 (.Y(n1614), 
	.B1(n10269), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6326));
   INVX1 U7535 (.Y(n10269), 
	.A(\ram[64][8] ));
   OAI22X1 U7536 (.Y(n1613), 
	.B1(n10270), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6328));
   INVX1 U7537 (.Y(n10270), 
	.A(\ram[64][7] ));
   OAI22X1 U7538 (.Y(n1612), 
	.B1(n10271), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6330));
   INVX1 U7539 (.Y(n10271), 
	.A(\ram[64][6] ));
   OAI22X1 U7540 (.Y(n1611), 
	.B1(n10272), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6332));
   INVX1 U7541 (.Y(n10272), 
	.A(\ram[64][5] ));
   OAI22X1 U7542 (.Y(n1610), 
	.B1(n10273), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6334));
   INVX1 U7543 (.Y(n10273), 
	.A(\ram[64][4] ));
   OAI22X1 U7544 (.Y(n1609), 
	.B1(n10274), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6336));
   INVX1 U7545 (.Y(n10274), 
	.A(\ram[64][3] ));
   OAI22X1 U7546 (.Y(n1608), 
	.B1(n10275), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6338));
   INVX1 U7547 (.Y(n10275), 
	.A(\ram[64][2] ));
   OAI22X1 U7548 (.Y(n1607), 
	.B1(n10276), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6306));
   INVX1 U7549 (.Y(n10276), 
	.A(\ram[64][1] ));
   OAI22X1 U7550 (.Y(n1606), 
	.B1(n10277), 
	.B0(n10261), 
	.A1(n10260), 
	.A0(n6309));
   INVX1 U7551 (.Y(n10277), 
	.A(\ram[64][0] ));
   NOR2BX1 U7552 (.Y(n10261), 
	.B(n10260), 
	.AN(mem_write_en));
   NAND2X1 U7553 (.Y(n10260), 
	.B(n6514), 
	.A(n10007));
   OAI22X1 U7554 (.Y(n1605), 
	.B1(n10280), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6311));
   INVX1 U7555 (.Y(n10280), 
	.A(\ram[63][15] ));
   OAI22X1 U7556 (.Y(n1604), 
	.B1(n10281), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6314));
   INVX1 U7557 (.Y(n10281), 
	.A(\ram[63][14] ));
   OAI22X1 U7558 (.Y(n1603), 
	.B1(n10282), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6316));
   INVX1 U7559 (.Y(n10282), 
	.A(\ram[63][13] ));
   OAI22X1 U7560 (.Y(n1602), 
	.B1(n10283), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6318));
   INVX1 U7561 (.Y(n10283), 
	.A(\ram[63][12] ));
   OAI22X1 U7562 (.Y(n1601), 
	.B1(n10284), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6320));
   INVX1 U7563 (.Y(n10284), 
	.A(\ram[63][11] ));
   OAI22X1 U7564 (.Y(n1600), 
	.B1(n10285), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6322));
   INVX1 U7565 (.Y(n10285), 
	.A(\ram[63][10] ));
   OAI22X1 U7566 (.Y(n1599), 
	.B1(n10286), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6324));
   INVX1 U7567 (.Y(n10286), 
	.A(\ram[63][9] ));
   OAI22X1 U7568 (.Y(n1598), 
	.B1(n10287), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6326));
   INVX1 U7569 (.Y(n10287), 
	.A(\ram[63][8] ));
   OAI22X1 U7570 (.Y(n1597), 
	.B1(n10288), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6328));
   INVX1 U7571 (.Y(n10288), 
	.A(\ram[63][7] ));
   OAI22X1 U7572 (.Y(n1596), 
	.B1(n10289), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6330));
   INVX1 U7573 (.Y(n10289), 
	.A(\ram[63][6] ));
   OAI22X1 U7574 (.Y(n1595), 
	.B1(n10290), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6332));
   INVX1 U7575 (.Y(n10290), 
	.A(\ram[63][5] ));
   OAI22X1 U7576 (.Y(n1594), 
	.B1(n10291), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6334));
   INVX1 U7577 (.Y(n10291), 
	.A(\ram[63][4] ));
   OAI22X1 U7578 (.Y(n1593), 
	.B1(n10292), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6336));
   INVX1 U7579 (.Y(n10292), 
	.A(\ram[63][3] ));
   OAI22X1 U7580 (.Y(n1592), 
	.B1(n10293), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6338));
   INVX1 U7581 (.Y(n10293), 
	.A(\ram[63][2] ));
   OAI22X1 U7582 (.Y(n1591), 
	.B1(n10294), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6306));
   INVX1 U7583 (.Y(n10294), 
	.A(\ram[63][1] ));
   OAI22X1 U7584 (.Y(n1590), 
	.B1(n10295), 
	.B0(n10279), 
	.A1(n10278), 
	.A0(n6309));
   INVX1 U7585 (.Y(n10295), 
	.A(\ram[63][0] ));
   NOR2BX1 U7586 (.Y(n10279), 
	.B(n10278), 
	.AN(mem_write_en));
   NAND2X1 U7587 (.Y(n10278), 
	.B(n6533), 
	.A(n10296));
   OAI22X1 U7588 (.Y(n1589), 
	.B1(n10299), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6311));
   INVX1 U7589 (.Y(n10299), 
	.A(\ram[62][15] ));
   OAI22X1 U7590 (.Y(n1588), 
	.B1(n10300), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6314));
   INVX1 U7591 (.Y(n10300), 
	.A(\ram[62][14] ));
   OAI22X1 U7592 (.Y(n1587), 
	.B1(n10301), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6316));
   INVX1 U7593 (.Y(n10301), 
	.A(\ram[62][13] ));
   OAI22X1 U7594 (.Y(n1586), 
	.B1(n10302), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6318));
   INVX1 U7595 (.Y(n10302), 
	.A(\ram[62][12] ));
   OAI22X1 U7596 (.Y(n1585), 
	.B1(n10303), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6320));
   INVX1 U7597 (.Y(n10303), 
	.A(\ram[62][11] ));
   OAI22X1 U7598 (.Y(n1584), 
	.B1(n10304), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6322));
   INVX1 U7599 (.Y(n10304), 
	.A(\ram[62][10] ));
   OAI22X1 U7600 (.Y(n1583), 
	.B1(n10305), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6324));
   INVX1 U7601 (.Y(n10305), 
	.A(\ram[62][9] ));
   OAI22X1 U7602 (.Y(n1582), 
	.B1(n10306), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6326));
   INVX1 U7603 (.Y(n10306), 
	.A(\ram[62][8] ));
   OAI22X1 U7604 (.Y(n1581), 
	.B1(n10307), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6328));
   INVX1 U7605 (.Y(n10307), 
	.A(\ram[62][7] ));
   OAI22X1 U7606 (.Y(n1580), 
	.B1(n10308), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6330));
   INVX1 U7607 (.Y(n10308), 
	.A(\ram[62][6] ));
   OAI22X1 U7608 (.Y(n1579), 
	.B1(n10309), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6332));
   INVX1 U7609 (.Y(n10309), 
	.A(\ram[62][5] ));
   OAI22X1 U7610 (.Y(n1578), 
	.B1(n10310), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6334));
   INVX1 U7611 (.Y(n10310), 
	.A(\ram[62][4] ));
   OAI22X1 U7612 (.Y(n1577), 
	.B1(n10311), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6336));
   INVX1 U7613 (.Y(n10311), 
	.A(\ram[62][3] ));
   OAI22X1 U7614 (.Y(n1576), 
	.B1(n10312), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6338));
   INVX1 U7615 (.Y(n10312), 
	.A(\ram[62][2] ));
   OAI22X1 U7616 (.Y(n1575), 
	.B1(n10313), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6306));
   INVX1 U7617 (.Y(n10313), 
	.A(\ram[62][1] ));
   OAI22X1 U7618 (.Y(n1574), 
	.B1(n10314), 
	.B0(n10298), 
	.A1(n10297), 
	.A0(n6309));
   INVX1 U7619 (.Y(n10314), 
	.A(\ram[62][0] ));
   NOR2BX1 U7620 (.Y(n10298), 
	.B(n10297), 
	.AN(mem_write_en));
   NAND2X1 U7621 (.Y(n10297), 
	.B(n6553), 
	.A(n10296));
   OAI22X1 U7622 (.Y(n1573), 
	.B1(n10317), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6311));
   INVX1 U7623 (.Y(n10317), 
	.A(\ram[61][15] ));
   OAI22X1 U7624 (.Y(n1572), 
	.B1(n10318), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6314));
   INVX1 U7625 (.Y(n10318), 
	.A(\ram[61][14] ));
   OAI22X1 U7626 (.Y(n1571), 
	.B1(n10319), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6316));
   INVX1 U7627 (.Y(n10319), 
	.A(\ram[61][13] ));
   OAI22X1 U7628 (.Y(n1570), 
	.B1(n10320), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6318));
   INVX1 U7629 (.Y(n10320), 
	.A(\ram[61][12] ));
   OAI22X1 U7630 (.Y(n1569), 
	.B1(n10321), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6320));
   INVX1 U7631 (.Y(n10321), 
	.A(\ram[61][11] ));
   OAI22X1 U7632 (.Y(n1568), 
	.B1(n10322), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6322));
   INVX1 U7633 (.Y(n10322), 
	.A(\ram[61][10] ));
   OAI22X1 U7634 (.Y(n1567), 
	.B1(n10323), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6324));
   INVX1 U7635 (.Y(n10323), 
	.A(\ram[61][9] ));
   OAI22X1 U7636 (.Y(n1566), 
	.B1(n10324), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6326));
   INVX1 U7637 (.Y(n10324), 
	.A(\ram[61][8] ));
   OAI22X1 U7638 (.Y(n1565), 
	.B1(n10325), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6328));
   INVX1 U7639 (.Y(n10325), 
	.A(\ram[61][7] ));
   OAI22X1 U7640 (.Y(n1564), 
	.B1(n10326), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6330));
   INVX1 U7641 (.Y(n10326), 
	.A(\ram[61][6] ));
   OAI22X1 U7642 (.Y(n1563), 
	.B1(n10327), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6332));
   INVX1 U7643 (.Y(n10327), 
	.A(\ram[61][5] ));
   OAI22X1 U7644 (.Y(n1562), 
	.B1(n10328), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6334));
   INVX1 U7645 (.Y(n10328), 
	.A(\ram[61][4] ));
   OAI22X1 U7646 (.Y(n1561), 
	.B1(n10329), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6336));
   INVX1 U7647 (.Y(n10329), 
	.A(\ram[61][3] ));
   OAI22X1 U7648 (.Y(n1560), 
	.B1(n10330), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6338));
   INVX1 U7649 (.Y(n10330), 
	.A(\ram[61][2] ));
   OAI22X1 U7650 (.Y(n1559), 
	.B1(n10331), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6306));
   INVX1 U7651 (.Y(n10331), 
	.A(\ram[61][1] ));
   OAI22X1 U7652 (.Y(n1558), 
	.B1(n10332), 
	.B0(n10316), 
	.A1(n10315), 
	.A0(n6309));
   INVX1 U7653 (.Y(n10332), 
	.A(\ram[61][0] ));
   NOR2BX1 U7654 (.Y(n10316), 
	.B(n10315), 
	.AN(mem_write_en));
   NAND2X1 U7655 (.Y(n10315), 
	.B(n6572), 
	.A(n10296));
   OAI22X1 U7656 (.Y(n1557), 
	.B1(n10335), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6311));
   INVX1 U7657 (.Y(n10335), 
	.A(\ram[60][15] ));
   OAI22X1 U7658 (.Y(n1556), 
	.B1(n10336), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6314));
   INVX1 U7659 (.Y(n10336), 
	.A(\ram[60][14] ));
   OAI22X1 U7660 (.Y(n1555), 
	.B1(n10337), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6316));
   INVX1 U7661 (.Y(n10337), 
	.A(\ram[60][13] ));
   OAI22X1 U7662 (.Y(n1554), 
	.B1(n10338), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6318));
   INVX1 U7663 (.Y(n10338), 
	.A(\ram[60][12] ));
   OAI22X1 U7664 (.Y(n1553), 
	.B1(n10339), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6320));
   INVX1 U7665 (.Y(n10339), 
	.A(\ram[60][11] ));
   OAI22X1 U7666 (.Y(n1552), 
	.B1(n10340), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6322));
   INVX1 U7667 (.Y(n10340), 
	.A(\ram[60][10] ));
   OAI22X1 U7668 (.Y(n1551), 
	.B1(n10341), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6324));
   INVX1 U7669 (.Y(n10341), 
	.A(\ram[60][9] ));
   OAI22X1 U7670 (.Y(n1550), 
	.B1(n10342), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6326));
   INVX1 U7671 (.Y(n10342), 
	.A(\ram[60][8] ));
   OAI22X1 U7672 (.Y(n1549), 
	.B1(n10343), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6328));
   INVX1 U7673 (.Y(n10343), 
	.A(\ram[60][7] ));
   OAI22X1 U7674 (.Y(n1548), 
	.B1(n10344), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6330));
   INVX1 U7675 (.Y(n10344), 
	.A(\ram[60][6] ));
   OAI22X1 U7676 (.Y(n1547), 
	.B1(n10345), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6332));
   INVX1 U7677 (.Y(n10345), 
	.A(\ram[60][5] ));
   OAI22X1 U7678 (.Y(n1546), 
	.B1(n10346), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6334));
   INVX1 U7679 (.Y(n10346), 
	.A(\ram[60][4] ));
   OAI22X1 U7680 (.Y(n1545), 
	.B1(n10347), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6336));
   INVX1 U7681 (.Y(n10347), 
	.A(\ram[60][3] ));
   OAI22X1 U7682 (.Y(n1544), 
	.B1(n10348), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6338));
   INVX1 U7683 (.Y(n10348), 
	.A(\ram[60][2] ));
   OAI22X1 U7684 (.Y(n1543), 
	.B1(n10349), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6306));
   INVX1 U7685 (.Y(n10349), 
	.A(\ram[60][1] ));
   OAI22X1 U7686 (.Y(n1542), 
	.B1(n10350), 
	.B0(n10334), 
	.A1(n10333), 
	.A0(n6309));
   INVX1 U7687 (.Y(n10350), 
	.A(\ram[60][0] ));
   NOR2BX1 U7688 (.Y(n10334), 
	.B(n10333), 
	.AN(mem_write_en));
   NAND2X1 U7689 (.Y(n10333), 
	.B(n6591), 
	.A(n10296));
   OAI22X1 U7690 (.Y(n1541), 
	.B1(n10353), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6311));
   INVX1 U7691 (.Y(n10353), 
	.A(\ram[59][15] ));
   OAI22X1 U7692 (.Y(n1540), 
	.B1(n10354), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6314));
   INVX1 U7693 (.Y(n10354), 
	.A(\ram[59][14] ));
   OAI22X1 U7694 (.Y(n1539), 
	.B1(n10355), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6316));
   INVX1 U7695 (.Y(n10355), 
	.A(\ram[59][13] ));
   OAI22X1 U7696 (.Y(n1538), 
	.B1(n10356), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6318));
   INVX1 U7697 (.Y(n10356), 
	.A(\ram[59][12] ));
   OAI22X1 U7698 (.Y(n1537), 
	.B1(n10357), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6320));
   INVX1 U7699 (.Y(n10357), 
	.A(\ram[59][11] ));
   OAI22X1 U7700 (.Y(n1536), 
	.B1(n10358), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6322));
   INVX1 U7701 (.Y(n10358), 
	.A(\ram[59][10] ));
   OAI22X1 U7702 (.Y(n1535), 
	.B1(n10359), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6324));
   INVX1 U7703 (.Y(n10359), 
	.A(\ram[59][9] ));
   OAI22X1 U7704 (.Y(n1534), 
	.B1(n10360), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6326));
   INVX1 U7705 (.Y(n10360), 
	.A(\ram[59][8] ));
   OAI22X1 U7706 (.Y(n1533), 
	.B1(n10361), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6328));
   INVX1 U7707 (.Y(n10361), 
	.A(\ram[59][7] ));
   OAI22X1 U7708 (.Y(n1532), 
	.B1(n10362), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6330));
   INVX1 U7709 (.Y(n10362), 
	.A(\ram[59][6] ));
   OAI22X1 U7710 (.Y(n1531), 
	.B1(n10363), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6332));
   INVX1 U7711 (.Y(n10363), 
	.A(\ram[59][5] ));
   OAI22X1 U7712 (.Y(n1530), 
	.B1(n10364), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6334));
   INVX1 U7713 (.Y(n10364), 
	.A(\ram[59][4] ));
   OAI22X1 U7714 (.Y(n1529), 
	.B1(n10365), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6336));
   INVX1 U7715 (.Y(n10365), 
	.A(\ram[59][3] ));
   OAI22X1 U7716 (.Y(n1528), 
	.B1(n10366), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6338));
   INVX1 U7717 (.Y(n10366), 
	.A(\ram[59][2] ));
   OAI22X1 U7718 (.Y(n1527), 
	.B1(n10367), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6306));
   INVX1 U7719 (.Y(n10367), 
	.A(\ram[59][1] ));
   OAI22X1 U7720 (.Y(n1526), 
	.B1(n10368), 
	.B0(n10352), 
	.A1(n10351), 
	.A0(n6309));
   INVX1 U7721 (.Y(n10368), 
	.A(\ram[59][0] ));
   NOR2BX1 U7722 (.Y(n10352), 
	.B(n10351), 
	.AN(mem_write_en));
   NAND2X1 U7723 (.Y(n10351), 
	.B(n6610), 
	.A(n10296));
   OAI22X1 U7724 (.Y(n1525), 
	.B1(n10371), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6311));
   INVX1 U7725 (.Y(n10371), 
	.A(\ram[58][15] ));
   OAI22X1 U7726 (.Y(n1524), 
	.B1(n10372), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6314));
   INVX1 U7727 (.Y(n10372), 
	.A(\ram[58][14] ));
   OAI22X1 U7728 (.Y(n1523), 
	.B1(n10373), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6316));
   INVX1 U7729 (.Y(n10373), 
	.A(\ram[58][13] ));
   OAI22X1 U7730 (.Y(n1522), 
	.B1(n10374), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6318));
   INVX1 U7731 (.Y(n10374), 
	.A(\ram[58][12] ));
   OAI22X1 U7732 (.Y(n1521), 
	.B1(n10375), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6320));
   INVX1 U7733 (.Y(n10375), 
	.A(\ram[58][11] ));
   OAI22X1 U7734 (.Y(n1520), 
	.B1(n10376), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6322));
   INVX1 U7735 (.Y(n10376), 
	.A(\ram[58][10] ));
   OAI22X1 U7736 (.Y(n1519), 
	.B1(n10377), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6324));
   INVX1 U7737 (.Y(n10377), 
	.A(\ram[58][9] ));
   OAI22X1 U7738 (.Y(n1518), 
	.B1(n10378), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6326));
   INVX1 U7739 (.Y(n10378), 
	.A(\ram[58][8] ));
   OAI22X1 U7740 (.Y(n1517), 
	.B1(n10379), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6328));
   INVX1 U7741 (.Y(n10379), 
	.A(\ram[58][7] ));
   OAI22X1 U7742 (.Y(n1516), 
	.B1(n10380), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6330));
   INVX1 U7743 (.Y(n10380), 
	.A(\ram[58][6] ));
   OAI22X1 U7744 (.Y(n1515), 
	.B1(n10381), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6332));
   INVX1 U7745 (.Y(n10381), 
	.A(\ram[58][5] ));
   OAI22X1 U7746 (.Y(n1514), 
	.B1(n10382), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6334));
   INVX1 U7747 (.Y(n10382), 
	.A(\ram[58][4] ));
   OAI22X1 U7748 (.Y(n1513), 
	.B1(n10383), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6336));
   INVX1 U7749 (.Y(n10383), 
	.A(\ram[58][3] ));
   OAI22X1 U7750 (.Y(n1512), 
	.B1(n10384), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6338));
   INVX1 U7751 (.Y(n10384), 
	.A(\ram[58][2] ));
   OAI22X1 U7752 (.Y(n1511), 
	.B1(n10385), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6306));
   INVX1 U7753 (.Y(n10385), 
	.A(\ram[58][1] ));
   OAI22X1 U7754 (.Y(n1510), 
	.B1(n10386), 
	.B0(n10370), 
	.A1(n10369), 
	.A0(n6309));
   INVX1 U7755 (.Y(n10386), 
	.A(\ram[58][0] ));
   NOR2BX1 U7756 (.Y(n10370), 
	.B(n10369), 
	.AN(mem_write_en));
   NAND2X1 U7757 (.Y(n10369), 
	.B(n6629), 
	.A(n10296));
   OAI22X1 U7758 (.Y(n1509), 
	.B1(n10389), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6311));
   INVX1 U7759 (.Y(n10389), 
	.A(\ram[57][15] ));
   OAI22X1 U7760 (.Y(n1508), 
	.B1(n10390), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6314));
   INVX1 U7761 (.Y(n10390), 
	.A(\ram[57][14] ));
   OAI22X1 U7762 (.Y(n1507), 
	.B1(n10391), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6316));
   INVX1 U7763 (.Y(n10391), 
	.A(\ram[57][13] ));
   OAI22X1 U7764 (.Y(n1506), 
	.B1(n10392), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6318));
   INVX1 U7765 (.Y(n10392), 
	.A(\ram[57][12] ));
   OAI22X1 U7766 (.Y(n1505), 
	.B1(n10393), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6320));
   INVX1 U7767 (.Y(n10393), 
	.A(\ram[57][11] ));
   OAI22X1 U7768 (.Y(n1504), 
	.B1(n10394), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6322));
   INVX1 U7769 (.Y(n10394), 
	.A(\ram[57][10] ));
   OAI22X1 U7770 (.Y(n1503), 
	.B1(n10395), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6324));
   INVX1 U7771 (.Y(n10395), 
	.A(\ram[57][9] ));
   OAI22X1 U7772 (.Y(n1502), 
	.B1(n10396), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6326));
   INVX1 U7773 (.Y(n10396), 
	.A(\ram[57][8] ));
   OAI22X1 U7774 (.Y(n1501), 
	.B1(n10397), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6328));
   INVX1 U7775 (.Y(n10397), 
	.A(\ram[57][7] ));
   OAI22X1 U7776 (.Y(n1500), 
	.B1(n10398), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6330));
   INVX1 U7777 (.Y(n10398), 
	.A(\ram[57][6] ));
   OAI22X1 U7778 (.Y(n1499), 
	.B1(n10399), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6332));
   INVX1 U7779 (.Y(n10399), 
	.A(\ram[57][5] ));
   OAI22X1 U7780 (.Y(n1498), 
	.B1(n10400), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6334));
   INVX1 U7781 (.Y(n10400), 
	.A(\ram[57][4] ));
   OAI22X1 U7782 (.Y(n1497), 
	.B1(n10401), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6336));
   INVX1 U7783 (.Y(n10401), 
	.A(\ram[57][3] ));
   OAI22X1 U7784 (.Y(n1496), 
	.B1(n10402), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6338));
   INVX1 U7785 (.Y(n10402), 
	.A(\ram[57][2] ));
   OAI22X1 U7786 (.Y(n1495), 
	.B1(n10403), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6306));
   INVX1 U7787 (.Y(n10403), 
	.A(\ram[57][1] ));
   OAI22X1 U7788 (.Y(n1494), 
	.B1(n10404), 
	.B0(n10388), 
	.A1(n10387), 
	.A0(n6309));
   INVX1 U7789 (.Y(n10404), 
	.A(\ram[57][0] ));
   NOR2BX1 U7790 (.Y(n10388), 
	.B(n10387), 
	.AN(mem_write_en));
   NAND2X1 U7791 (.Y(n10387), 
	.B(n6342), 
	.A(n10296));
   OAI22X1 U7792 (.Y(n1493), 
	.B1(n10407), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6311));
   INVX1 U7793 (.Y(n10407), 
	.A(\ram[56][15] ));
   OAI22X1 U7794 (.Y(n1492), 
	.B1(n10408), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6314));
   INVX1 U7795 (.Y(n10408), 
	.A(\ram[56][14] ));
   OAI22X1 U7796 (.Y(n1491), 
	.B1(n10409), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6316));
   INVX1 U7797 (.Y(n10409), 
	.A(\ram[56][13] ));
   OAI22X1 U7798 (.Y(n1490), 
	.B1(n10410), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6318));
   INVX1 U7799 (.Y(n10410), 
	.A(\ram[56][12] ));
   OAI22X1 U7800 (.Y(n1489), 
	.B1(n10411), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6320));
   INVX1 U7801 (.Y(n10411), 
	.A(\ram[56][11] ));
   OAI22X1 U7802 (.Y(n1488), 
	.B1(n10412), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6322));
   INVX1 U7803 (.Y(n10412), 
	.A(\ram[56][10] ));
   OAI22X1 U7804 (.Y(n1487), 
	.B1(n10413), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6324));
   INVX1 U7805 (.Y(n10413), 
	.A(\ram[56][9] ));
   OAI22X1 U7806 (.Y(n1486), 
	.B1(n10414), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6326));
   INVX1 U7807 (.Y(n10414), 
	.A(\ram[56][8] ));
   OAI22X1 U7808 (.Y(n1485), 
	.B1(n10415), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6328));
   INVX1 U7809 (.Y(n10415), 
	.A(\ram[56][7] ));
   OAI22X1 U7810 (.Y(n1484), 
	.B1(n10416), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6330));
   INVX1 U7811 (.Y(n10416), 
	.A(\ram[56][6] ));
   OAI22X1 U7812 (.Y(n1483), 
	.B1(n10417), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6332));
   INVX1 U7813 (.Y(n10417), 
	.A(\ram[56][5] ));
   OAI22X1 U7814 (.Y(n1482), 
	.B1(n10418), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6334));
   INVX1 U7815 (.Y(n10418), 
	.A(\ram[56][4] ));
   OAI22X1 U7816 (.Y(n1481), 
	.B1(n10419), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6336));
   INVX1 U7817 (.Y(n10419), 
	.A(\ram[56][3] ));
   OAI22X1 U7818 (.Y(n1480), 
	.B1(n10420), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6338));
   INVX1 U7819 (.Y(n10420), 
	.A(\ram[56][2] ));
   OAI22X1 U7820 (.Y(n1479), 
	.B1(n10421), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6306));
   INVX1 U7821 (.Y(n10421), 
	.A(\ram[56][1] ));
   OAI22X1 U7822 (.Y(n1478), 
	.B1(n10422), 
	.B0(n10406), 
	.A1(n10405), 
	.A0(n6309));
   INVX1 U7823 (.Y(n10422), 
	.A(\ram[56][0] ));
   NOR2BX1 U7824 (.Y(n10406), 
	.B(n10405), 
	.AN(mem_write_en));
   NAND2X1 U7825 (.Y(n10405), 
	.B(n6362), 
	.A(n10296));
   OAI22X1 U7826 (.Y(n1477), 
	.B1(n10425), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6311));
   INVX1 U7827 (.Y(n10425), 
	.A(\ram[55][15] ));
   OAI22X1 U7828 (.Y(n1476), 
	.B1(n10426), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6314));
   INVX1 U7829 (.Y(n10426), 
	.A(\ram[55][14] ));
   OAI22X1 U7830 (.Y(n1475), 
	.B1(n10427), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6316));
   INVX1 U7831 (.Y(n10427), 
	.A(\ram[55][13] ));
   OAI22X1 U7832 (.Y(n1474), 
	.B1(n10428), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6318));
   INVX1 U7833 (.Y(n10428), 
	.A(\ram[55][12] ));
   OAI22X1 U7834 (.Y(n1473), 
	.B1(n10429), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6320));
   INVX1 U7835 (.Y(n10429), 
	.A(\ram[55][11] ));
   OAI22X1 U7836 (.Y(n1472), 
	.B1(n10430), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6322));
   INVX1 U7837 (.Y(n10430), 
	.A(\ram[55][10] ));
   OAI22X1 U7838 (.Y(n1471), 
	.B1(n10431), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6324));
   INVX1 U7839 (.Y(n10431), 
	.A(\ram[55][9] ));
   OAI22X1 U7840 (.Y(n1470), 
	.B1(n10432), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6326));
   INVX1 U7841 (.Y(n10432), 
	.A(\ram[55][8] ));
   OAI22X1 U7842 (.Y(n1469), 
	.B1(n10433), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6328));
   INVX1 U7843 (.Y(n10433), 
	.A(\ram[55][7] ));
   OAI22X1 U7844 (.Y(n1468), 
	.B1(n10434), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6330));
   INVX1 U7845 (.Y(n10434), 
	.A(\ram[55][6] ));
   OAI22X1 U7846 (.Y(n1467), 
	.B1(n10435), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6332));
   INVX1 U7847 (.Y(n10435), 
	.A(\ram[55][5] ));
   OAI22X1 U7848 (.Y(n1466), 
	.B1(n10436), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6334));
   INVX1 U7849 (.Y(n10436), 
	.A(\ram[55][4] ));
   OAI22X1 U7850 (.Y(n1465), 
	.B1(n10437), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6336));
   INVX1 U7851 (.Y(n10437), 
	.A(\ram[55][3] ));
   OAI22X1 U7852 (.Y(n1464), 
	.B1(n10438), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6338));
   INVX1 U7853 (.Y(n10438), 
	.A(\ram[55][2] ));
   OAI22X1 U7854 (.Y(n1463), 
	.B1(n10439), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6306));
   INVX1 U7855 (.Y(n10439), 
	.A(\ram[55][1] ));
   OAI22X1 U7856 (.Y(n1462), 
	.B1(n10440), 
	.B0(n10424), 
	.A1(n10423), 
	.A0(n6309));
   INVX1 U7857 (.Y(n10440), 
	.A(\ram[55][0] ));
   NOR2BX1 U7858 (.Y(n10424), 
	.B(n10423), 
	.AN(mem_write_en));
   NAND2X1 U7859 (.Y(n10423), 
	.B(n6381), 
	.A(n10296));
   OAI22X1 U7860 (.Y(n1461), 
	.B1(n10443), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6311));
   INVX1 U7861 (.Y(n10443), 
	.A(\ram[54][15] ));
   OAI22X1 U7862 (.Y(n1460), 
	.B1(n10444), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6314));
   INVX1 U7863 (.Y(n10444), 
	.A(\ram[54][14] ));
   OAI22X1 U7864 (.Y(n1459), 
	.B1(n10445), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6316));
   INVX1 U7865 (.Y(n10445), 
	.A(\ram[54][13] ));
   OAI22X1 U7866 (.Y(n1458), 
	.B1(n10446), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6318));
   INVX1 U7867 (.Y(n10446), 
	.A(\ram[54][12] ));
   OAI22X1 U7868 (.Y(n1457), 
	.B1(n10447), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6320));
   INVX1 U7869 (.Y(n10447), 
	.A(\ram[54][11] ));
   OAI22X1 U7870 (.Y(n1456), 
	.B1(n10448), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6322));
   INVX1 U7871 (.Y(n10448), 
	.A(\ram[54][10] ));
   OAI22X1 U7872 (.Y(n1455), 
	.B1(n10449), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6324));
   INVX1 U7873 (.Y(n10449), 
	.A(\ram[54][9] ));
   OAI22X1 U7874 (.Y(n1454), 
	.B1(n10450), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6326));
   INVX1 U7875 (.Y(n10450), 
	.A(\ram[54][8] ));
   OAI22X1 U7876 (.Y(n1453), 
	.B1(n10451), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6328));
   INVX1 U7877 (.Y(n10451), 
	.A(\ram[54][7] ));
   OAI22X1 U7878 (.Y(n1452), 
	.B1(n10452), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6330));
   INVX1 U7879 (.Y(n10452), 
	.A(\ram[54][6] ));
   OAI22X1 U7880 (.Y(n1451), 
	.B1(n10453), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6332));
   INVX1 U7881 (.Y(n10453), 
	.A(\ram[54][5] ));
   OAI22X1 U7882 (.Y(n1450), 
	.B1(n10454), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6334));
   INVX1 U7883 (.Y(n10454), 
	.A(\ram[54][4] ));
   OAI22X1 U7884 (.Y(n1449), 
	.B1(n10455), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6336));
   INVX1 U7885 (.Y(n10455), 
	.A(\ram[54][3] ));
   OAI22X1 U7886 (.Y(n1448), 
	.B1(n10456), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6338));
   INVX1 U7887 (.Y(n10456), 
	.A(\ram[54][2] ));
   OAI22X1 U7888 (.Y(n1447), 
	.B1(n10457), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6306));
   INVX1 U7889 (.Y(n10457), 
	.A(\ram[54][1] ));
   OAI22X1 U7890 (.Y(n1446), 
	.B1(n10458), 
	.B0(n10442), 
	.A1(n10441), 
	.A0(n6309));
   INVX1 U7891 (.Y(n10458), 
	.A(\ram[54][0] ));
   NOR2BX1 U7892 (.Y(n10442), 
	.B(n10441), 
	.AN(mem_write_en));
   NAND2X1 U7893 (.Y(n10441), 
	.B(n6400), 
	.A(n10296));
   OAI22X1 U7894 (.Y(n1445), 
	.B1(n10461), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6311));
   INVX1 U7895 (.Y(n10461), 
	.A(\ram[53][15] ));
   OAI22X1 U7896 (.Y(n1444), 
	.B1(n10462), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6314));
   INVX1 U7897 (.Y(n10462), 
	.A(\ram[53][14] ));
   OAI22X1 U7898 (.Y(n1443), 
	.B1(n10463), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6316));
   INVX1 U7899 (.Y(n10463), 
	.A(\ram[53][13] ));
   OAI22X1 U7900 (.Y(n1442), 
	.B1(n10464), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6318));
   INVX1 U7901 (.Y(n10464), 
	.A(\ram[53][12] ));
   OAI22X1 U7902 (.Y(n1441), 
	.B1(n10465), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6320));
   INVX1 U7903 (.Y(n10465), 
	.A(\ram[53][11] ));
   OAI22X1 U7904 (.Y(n1440), 
	.B1(n10466), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6322));
   INVX1 U7905 (.Y(n10466), 
	.A(\ram[53][10] ));
   OAI22X1 U7906 (.Y(n1439), 
	.B1(n10467), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6324));
   INVX1 U7907 (.Y(n10467), 
	.A(\ram[53][9] ));
   OAI22X1 U7908 (.Y(n1438), 
	.B1(n10468), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6326));
   INVX1 U7909 (.Y(n10468), 
	.A(\ram[53][8] ));
   OAI22X1 U7910 (.Y(n1437), 
	.B1(n10469), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6328));
   INVX1 U7911 (.Y(n10469), 
	.A(\ram[53][7] ));
   OAI22X1 U7912 (.Y(n1436), 
	.B1(n10470), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6330));
   INVX1 U7913 (.Y(n10470), 
	.A(\ram[53][6] ));
   OAI22X1 U7914 (.Y(n1435), 
	.B1(n10471), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6332));
   INVX1 U7915 (.Y(n10471), 
	.A(\ram[53][5] ));
   OAI22X1 U7916 (.Y(n1434), 
	.B1(n10472), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6334));
   INVX1 U7917 (.Y(n10472), 
	.A(\ram[53][4] ));
   OAI22X1 U7918 (.Y(n1433), 
	.B1(n10473), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6336));
   INVX1 U7919 (.Y(n10473), 
	.A(\ram[53][3] ));
   OAI22X1 U7920 (.Y(n1432), 
	.B1(n10474), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6338));
   INVX1 U7921 (.Y(n10474), 
	.A(\ram[53][2] ));
   OAI22X1 U7922 (.Y(n1431), 
	.B1(n10475), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6306));
   INVX1 U7923 (.Y(n10475), 
	.A(\ram[53][1] ));
   OAI22X1 U7924 (.Y(n1430), 
	.B1(n10476), 
	.B0(n10460), 
	.A1(n10459), 
	.A0(n6309));
   INVX1 U7925 (.Y(n10476), 
	.A(\ram[53][0] ));
   NOR2BX1 U7926 (.Y(n10460), 
	.B(n10459), 
	.AN(mem_write_en));
   NAND2X1 U7927 (.Y(n10459), 
	.B(n6419), 
	.A(n10296));
   OAI22X1 U7928 (.Y(n1429), 
	.B1(n10479), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6311));
   INVX1 U7929 (.Y(n10479), 
	.A(\ram[52][15] ));
   OAI22X1 U7930 (.Y(n1428), 
	.B1(n10480), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6314));
   INVX1 U7931 (.Y(n10480), 
	.A(\ram[52][14] ));
   OAI22X1 U7932 (.Y(n1427), 
	.B1(n10481), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6316));
   INVX1 U7933 (.Y(n10481), 
	.A(\ram[52][13] ));
   OAI22X1 U7934 (.Y(n1426), 
	.B1(n10482), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6318));
   INVX1 U7935 (.Y(n10482), 
	.A(\ram[52][12] ));
   OAI22X1 U7936 (.Y(n1425), 
	.B1(n10483), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6320));
   INVX1 U7937 (.Y(n10483), 
	.A(\ram[52][11] ));
   OAI22X1 U7938 (.Y(n1424), 
	.B1(n10484), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6322));
   INVX1 U7939 (.Y(n10484), 
	.A(\ram[52][10] ));
   OAI22X1 U7940 (.Y(n1423), 
	.B1(n10485), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6324));
   INVX1 U7941 (.Y(n10485), 
	.A(\ram[52][9] ));
   OAI22X1 U7942 (.Y(n1422), 
	.B1(n10486), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6326));
   INVX1 U7943 (.Y(n10486), 
	.A(\ram[52][8] ));
   OAI22X1 U7944 (.Y(n1421), 
	.B1(n10487), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6328));
   INVX1 U7945 (.Y(n10487), 
	.A(\ram[52][7] ));
   OAI22X1 U7946 (.Y(n1420), 
	.B1(n10488), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6330));
   INVX1 U7947 (.Y(n10488), 
	.A(\ram[52][6] ));
   OAI22X1 U7948 (.Y(n1419), 
	.B1(n10489), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6332));
   INVX1 U7949 (.Y(n10489), 
	.A(\ram[52][5] ));
   OAI22X1 U7950 (.Y(n1418), 
	.B1(n10490), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6334));
   INVX1 U7951 (.Y(n10490), 
	.A(\ram[52][4] ));
   OAI22X1 U7952 (.Y(n1417), 
	.B1(n10491), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6336));
   INVX1 U7953 (.Y(n10491), 
	.A(\ram[52][3] ));
   OAI22X1 U7954 (.Y(n1416), 
	.B1(n10492), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6338));
   INVX1 U7955 (.Y(n10492), 
	.A(\ram[52][2] ));
   OAI22X1 U7956 (.Y(n1415), 
	.B1(n10493), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6306));
   INVX1 U7957 (.Y(n10493), 
	.A(\ram[52][1] ));
   OAI22X1 U7958 (.Y(n1414), 
	.B1(n10494), 
	.B0(n10478), 
	.A1(n10477), 
	.A0(n6309));
   INVX1 U7959 (.Y(n10494), 
	.A(\ram[52][0] ));
   NOR2BX1 U7960 (.Y(n10478), 
	.B(n10477), 
	.AN(mem_write_en));
   NAND2X1 U7961 (.Y(n10477), 
	.B(n6438), 
	.A(n10296));
   OAI22X1 U7962 (.Y(n1413), 
	.B1(n10497), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6311));
   INVX1 U7963 (.Y(n10497), 
	.A(\ram[51][15] ));
   OAI22X1 U7964 (.Y(n1412), 
	.B1(n10498), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6314));
   INVX1 U7965 (.Y(n10498), 
	.A(\ram[51][14] ));
   OAI22X1 U7966 (.Y(n1411), 
	.B1(n10499), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6316));
   INVX1 U7967 (.Y(n10499), 
	.A(\ram[51][13] ));
   OAI22X1 U7968 (.Y(n1410), 
	.B1(n10500), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6318));
   INVX1 U7969 (.Y(n10500), 
	.A(\ram[51][12] ));
   OAI22X1 U7970 (.Y(n1409), 
	.B1(n10501), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6320));
   INVX1 U7971 (.Y(n10501), 
	.A(\ram[51][11] ));
   OAI22X1 U7972 (.Y(n1408), 
	.B1(n10502), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6322));
   INVX1 U7973 (.Y(n10502), 
	.A(\ram[51][10] ));
   OAI22X1 U7974 (.Y(n1407), 
	.B1(n10503), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6324));
   INVX1 U7975 (.Y(n10503), 
	.A(\ram[51][9] ));
   OAI22X1 U7976 (.Y(n1406), 
	.B1(n10504), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6326));
   INVX1 U7977 (.Y(n10504), 
	.A(\ram[51][8] ));
   OAI22X1 U7978 (.Y(n1405), 
	.B1(n10505), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6328));
   INVX1 U7979 (.Y(n10505), 
	.A(\ram[51][7] ));
   OAI22X1 U7980 (.Y(n1404), 
	.B1(n10506), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6330));
   INVX1 U7981 (.Y(n10506), 
	.A(\ram[51][6] ));
   OAI22X1 U7982 (.Y(n1403), 
	.B1(n10507), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6332));
   INVX1 U7983 (.Y(n10507), 
	.A(\ram[51][5] ));
   OAI22X1 U7984 (.Y(n1402), 
	.B1(n10508), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6334));
   INVX1 U7985 (.Y(n10508), 
	.A(\ram[51][4] ));
   OAI22X1 U7986 (.Y(n1401), 
	.B1(n10509), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6336));
   INVX1 U7987 (.Y(n10509), 
	.A(\ram[51][3] ));
   OAI22X1 U7988 (.Y(n1400), 
	.B1(n10510), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6338));
   INVX1 U7989 (.Y(n10510), 
	.A(\ram[51][2] ));
   OAI22X1 U7990 (.Y(n1399), 
	.B1(n10511), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6306));
   INVX1 U7991 (.Y(n10511), 
	.A(\ram[51][1] ));
   OAI22X1 U7992 (.Y(n1398), 
	.B1(n10512), 
	.B0(n10496), 
	.A1(n10495), 
	.A0(n6309));
   INVX1 U7993 (.Y(n10512), 
	.A(\ram[51][0] ));
   NOR2BX1 U7994 (.Y(n10496), 
	.B(n10495), 
	.AN(mem_write_en));
   NAND2X1 U7995 (.Y(n10495), 
	.B(n6457), 
	.A(n10296));
   OAI22X1 U7996 (.Y(n1397), 
	.B1(n10515), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6311));
   INVX1 U7997 (.Y(n10515), 
	.A(\ram[50][15] ));
   OAI22X1 U7998 (.Y(n1396), 
	.B1(n10516), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6314));
   INVX1 U7999 (.Y(n10516), 
	.A(\ram[50][14] ));
   OAI22X1 U8000 (.Y(n1395), 
	.B1(n10517), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6316));
   INVX1 U8001 (.Y(n10517), 
	.A(\ram[50][13] ));
   OAI22X1 U8002 (.Y(n1394), 
	.B1(n10518), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6318));
   INVX1 U8003 (.Y(n10518), 
	.A(\ram[50][12] ));
   OAI22X1 U8004 (.Y(n1393), 
	.B1(n10519), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6320));
   INVX1 U8005 (.Y(n10519), 
	.A(\ram[50][11] ));
   OAI22X1 U8006 (.Y(n1392), 
	.B1(n10520), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6322));
   INVX1 U8007 (.Y(n10520), 
	.A(\ram[50][10] ));
   OAI22X1 U8008 (.Y(n1391), 
	.B1(n10521), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6324));
   INVX1 U8009 (.Y(n10521), 
	.A(\ram[50][9] ));
   OAI22X1 U8010 (.Y(n1390), 
	.B1(n10522), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6326));
   INVX1 U8011 (.Y(n10522), 
	.A(\ram[50][8] ));
   OAI22X1 U8012 (.Y(n1389), 
	.B1(n10523), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6328));
   INVX1 U8013 (.Y(n10523), 
	.A(\ram[50][7] ));
   OAI22X1 U8014 (.Y(n1388), 
	.B1(n10524), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6330));
   INVX1 U8015 (.Y(n10524), 
	.A(\ram[50][6] ));
   OAI22X1 U8016 (.Y(n1387), 
	.B1(n10525), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6332));
   INVX1 U8017 (.Y(n10525), 
	.A(\ram[50][5] ));
   OAI22X1 U8018 (.Y(n1386), 
	.B1(n10526), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6334));
   INVX1 U8019 (.Y(n10526), 
	.A(\ram[50][4] ));
   OAI22X1 U8020 (.Y(n1385), 
	.B1(n10527), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6336));
   INVX1 U8021 (.Y(n10527), 
	.A(\ram[50][3] ));
   OAI22X1 U8022 (.Y(n1384), 
	.B1(n10528), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6338));
   INVX1 U8023 (.Y(n10528), 
	.A(\ram[50][2] ));
   OAI22X1 U8024 (.Y(n1383), 
	.B1(n10529), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6306));
   INVX1 U8025 (.Y(n10529), 
	.A(\ram[50][1] ));
   OAI22X1 U8026 (.Y(n1382), 
	.B1(n10530), 
	.B0(n10514), 
	.A1(n10513), 
	.A0(n6309));
   INVX1 U8027 (.Y(n10530), 
	.A(\ram[50][0] ));
   NOR2BX1 U8028 (.Y(n10514), 
	.B(n10513), 
	.AN(mem_write_en));
   NAND2X1 U8029 (.Y(n10513), 
	.B(n6476), 
	.A(n10296));
   OAI22X1 U8030 (.Y(n1381), 
	.B1(n10533), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6311));
   INVX1 U8031 (.Y(n10533), 
	.A(\ram[49][15] ));
   OAI22X1 U8032 (.Y(n1380), 
	.B1(n10534), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6314));
   INVX1 U8033 (.Y(n10534), 
	.A(\ram[49][14] ));
   OAI22X1 U8034 (.Y(n1379), 
	.B1(n10535), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6316));
   INVX1 U8035 (.Y(n10535), 
	.A(\ram[49][13] ));
   OAI22X1 U8036 (.Y(n1378), 
	.B1(n10536), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6318));
   INVX1 U8037 (.Y(n10536), 
	.A(\ram[49][12] ));
   OAI22X1 U8038 (.Y(n1377), 
	.B1(n10537), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6320));
   INVX1 U8039 (.Y(n10537), 
	.A(\ram[49][11] ));
   OAI22X1 U8040 (.Y(n1376), 
	.B1(n10538), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6322));
   INVX1 U8041 (.Y(n10538), 
	.A(\ram[49][10] ));
   OAI22X1 U8042 (.Y(n1375), 
	.B1(n10539), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6324));
   INVX1 U8043 (.Y(n10539), 
	.A(\ram[49][9] ));
   OAI22X1 U8044 (.Y(n1374), 
	.B1(n10540), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6326));
   INVX1 U8045 (.Y(n10540), 
	.A(\ram[49][8] ));
   OAI22X1 U8046 (.Y(n1373), 
	.B1(n10541), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6328));
   INVX1 U8047 (.Y(n10541), 
	.A(\ram[49][7] ));
   OAI22X1 U8048 (.Y(n1372), 
	.B1(n10542), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6330));
   INVX1 U8049 (.Y(n10542), 
	.A(\ram[49][6] ));
   OAI22X1 U8050 (.Y(n1371), 
	.B1(n10543), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6332));
   INVX1 U8051 (.Y(n10543), 
	.A(\ram[49][5] ));
   OAI22X1 U8052 (.Y(n1370), 
	.B1(n10544), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6334));
   INVX1 U8053 (.Y(n10544), 
	.A(\ram[49][4] ));
   OAI22X1 U8054 (.Y(n1369), 
	.B1(n10545), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6336));
   INVX1 U8055 (.Y(n10545), 
	.A(\ram[49][3] ));
   OAI22X1 U8056 (.Y(n1368), 
	.B1(n10546), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6338));
   INVX1 U8057 (.Y(n10546), 
	.A(\ram[49][2] ));
   OAI22X1 U8058 (.Y(n1367), 
	.B1(n10547), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6306));
   INVX1 U8059 (.Y(n10547), 
	.A(\ram[49][1] ));
   OAI22X1 U8060 (.Y(n1366), 
	.B1(n10548), 
	.B0(n10532), 
	.A1(n10531), 
	.A0(n6309));
   INVX1 U8061 (.Y(n10548), 
	.A(\ram[49][0] ));
   NOR2BX1 U8062 (.Y(n10532), 
	.B(n10531), 
	.AN(mem_write_en));
   NAND2X1 U8063 (.Y(n10531), 
	.B(n6495), 
	.A(n10296));
   OAI22X1 U8064 (.Y(n1365), 
	.B1(n10551), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6311));
   INVX1 U8065 (.Y(n10551), 
	.A(\ram[48][15] ));
   OAI22X1 U8066 (.Y(n1364), 
	.B1(n10552), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6314));
   INVX1 U8067 (.Y(n10552), 
	.A(\ram[48][14] ));
   OAI22X1 U8068 (.Y(n1363), 
	.B1(n10553), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6316));
   INVX1 U8069 (.Y(n10553), 
	.A(\ram[48][13] ));
   OAI22X1 U8070 (.Y(n1362), 
	.B1(n10554), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6318));
   INVX1 U8071 (.Y(n10554), 
	.A(\ram[48][12] ));
   OAI22X1 U8072 (.Y(n1361), 
	.B1(n10555), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6320));
   INVX1 U8073 (.Y(n10555), 
	.A(\ram[48][11] ));
   OAI22X1 U8074 (.Y(n1360), 
	.B1(n10556), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6322));
   INVX1 U8075 (.Y(n10556), 
	.A(\ram[48][10] ));
   OAI22X1 U8076 (.Y(n1359), 
	.B1(n10557), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6324));
   INVX1 U8077 (.Y(n10557), 
	.A(\ram[48][9] ));
   OAI22X1 U8078 (.Y(n1358), 
	.B1(n10558), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6326));
   INVX1 U8079 (.Y(n10558), 
	.A(\ram[48][8] ));
   OAI22X1 U8080 (.Y(n1357), 
	.B1(n10559), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6328));
   INVX1 U8081 (.Y(n10559), 
	.A(\ram[48][7] ));
   OAI22X1 U8082 (.Y(n1356), 
	.B1(n10560), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6330));
   INVX1 U8083 (.Y(n10560), 
	.A(\ram[48][6] ));
   OAI22X1 U8084 (.Y(n1355), 
	.B1(n10561), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6332));
   INVX1 U8085 (.Y(n10561), 
	.A(\ram[48][5] ));
   OAI22X1 U8086 (.Y(n1354), 
	.B1(n10562), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6334));
   INVX1 U8087 (.Y(n10562), 
	.A(\ram[48][4] ));
   OAI22X1 U8088 (.Y(n1353), 
	.B1(n10563), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6336));
   INVX1 U8089 (.Y(n10563), 
	.A(\ram[48][3] ));
   OAI22X1 U8090 (.Y(n1352), 
	.B1(n10564), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6338));
   INVX1 U8091 (.Y(n10564), 
	.A(\ram[48][2] ));
   OAI22X1 U8092 (.Y(n1351), 
	.B1(n10565), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6306));
   INVX1 U8093 (.Y(n10565), 
	.A(\ram[48][1] ));
   OAI22X1 U8094 (.Y(n1350), 
	.B1(n10566), 
	.B0(n10550), 
	.A1(n10549), 
	.A0(n6309));
   INVX1 U8095 (.Y(n10566), 
	.A(\ram[48][0] ));
   NOR2BX1 U8096 (.Y(n10550), 
	.B(n10549), 
	.AN(mem_write_en));
   NAND2X1 U8097 (.Y(n10549), 
	.B(n6514), 
	.A(n10296));
   OAI22X1 U8098 (.Y(n1349), 
	.B1(n10569), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6311));
   INVX1 U8099 (.Y(n10569), 
	.A(\ram[47][15] ));
   OAI22X1 U8100 (.Y(n1348), 
	.B1(n10570), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6314));
   INVX1 U8101 (.Y(n10570), 
	.A(\ram[47][14] ));
   OAI22X1 U8102 (.Y(n1347), 
	.B1(n10571), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6316));
   INVX1 U8103 (.Y(n10571), 
	.A(\ram[47][13] ));
   OAI22X1 U8104 (.Y(n1346), 
	.B1(n10572), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6318));
   INVX1 U8105 (.Y(n10572), 
	.A(\ram[47][12] ));
   OAI22X1 U8106 (.Y(n1345), 
	.B1(n10573), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6320));
   INVX1 U8107 (.Y(n10573), 
	.A(\ram[47][11] ));
   OAI22X1 U8108 (.Y(n1344), 
	.B1(n10574), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6322));
   INVX1 U8109 (.Y(n10574), 
	.A(\ram[47][10] ));
   OAI22X1 U8110 (.Y(n1343), 
	.B1(n10575), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6324));
   INVX1 U8111 (.Y(n10575), 
	.A(\ram[47][9] ));
   OAI22X1 U8112 (.Y(n1342), 
	.B1(n10576), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6326));
   INVX1 U8113 (.Y(n10576), 
	.A(\ram[47][8] ));
   OAI22X1 U8114 (.Y(n1341), 
	.B1(n10577), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6328));
   INVX1 U8115 (.Y(n10577), 
	.A(\ram[47][7] ));
   OAI22X1 U8116 (.Y(n1340), 
	.B1(n10578), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6330));
   INVX1 U8117 (.Y(n10578), 
	.A(\ram[47][6] ));
   OAI22X1 U8118 (.Y(n1339), 
	.B1(n10579), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6332));
   INVX1 U8119 (.Y(n10579), 
	.A(\ram[47][5] ));
   OAI22X1 U8120 (.Y(n1338), 
	.B1(n10580), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6334));
   INVX1 U8121 (.Y(n10580), 
	.A(\ram[47][4] ));
   OAI22X1 U8122 (.Y(n1337), 
	.B1(n10581), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6336));
   INVX1 U8123 (.Y(n10581), 
	.A(\ram[47][3] ));
   OAI22X1 U8124 (.Y(n1336), 
	.B1(n10582), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6338));
   INVX1 U8125 (.Y(n10582), 
	.A(\ram[47][2] ));
   OAI22X1 U8126 (.Y(n1335), 
	.B1(n10583), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6306));
   INVX1 U8127 (.Y(n10583), 
	.A(\ram[47][1] ));
   OAI22X1 U8128 (.Y(n1334), 
	.B1(n10584), 
	.B0(n10568), 
	.A1(n10567), 
	.A0(n6309));
   INVX1 U8129 (.Y(n10584), 
	.A(\ram[47][0] ));
   NOR2BX1 U8130 (.Y(n10568), 
	.B(n10567), 
	.AN(mem_write_en));
   NAND2X1 U8131 (.Y(n10567), 
	.B(n6533), 
	.A(n10585));
   OAI22X1 U8132 (.Y(n1333), 
	.B1(n10588), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6311));
   INVX1 U8133 (.Y(n10588), 
	.A(\ram[46][15] ));
   OAI22X1 U8134 (.Y(n1332), 
	.B1(n10589), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6314));
   INVX1 U8135 (.Y(n10589), 
	.A(\ram[46][14] ));
   OAI22X1 U8136 (.Y(n1331), 
	.B1(n10590), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6316));
   INVX1 U8137 (.Y(n10590), 
	.A(\ram[46][13] ));
   OAI22X1 U8138 (.Y(n1330), 
	.B1(n10591), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6318));
   INVX1 U8139 (.Y(n10591), 
	.A(\ram[46][12] ));
   OAI22X1 U8140 (.Y(n1329), 
	.B1(n10592), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6320));
   INVX1 U8141 (.Y(n10592), 
	.A(\ram[46][11] ));
   OAI22X1 U8142 (.Y(n1328), 
	.B1(n10593), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6322));
   INVX1 U8143 (.Y(n10593), 
	.A(\ram[46][10] ));
   OAI22X1 U8144 (.Y(n1327), 
	.B1(n10594), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6324));
   INVX1 U8145 (.Y(n10594), 
	.A(\ram[46][9] ));
   OAI22X1 U8146 (.Y(n1326), 
	.B1(n10595), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6326));
   INVX1 U8147 (.Y(n10595), 
	.A(\ram[46][8] ));
   OAI22X1 U8148 (.Y(n1325), 
	.B1(n10596), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6328));
   INVX1 U8149 (.Y(n10596), 
	.A(\ram[46][7] ));
   OAI22X1 U8150 (.Y(n1324), 
	.B1(n10597), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6330));
   INVX1 U8151 (.Y(n10597), 
	.A(\ram[46][6] ));
   OAI22X1 U8152 (.Y(n1323), 
	.B1(n10598), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6332));
   INVX1 U8153 (.Y(n10598), 
	.A(\ram[46][5] ));
   OAI22X1 U8154 (.Y(n1322), 
	.B1(n10599), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6334));
   INVX1 U8155 (.Y(n10599), 
	.A(\ram[46][4] ));
   OAI22X1 U8156 (.Y(n1321), 
	.B1(n10600), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6336));
   INVX1 U8157 (.Y(n10600), 
	.A(\ram[46][3] ));
   OAI22X1 U8158 (.Y(n1320), 
	.B1(n10601), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6338));
   INVX1 U8159 (.Y(n10601), 
	.A(\ram[46][2] ));
   OAI22X1 U8160 (.Y(n1319), 
	.B1(n10602), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6306));
   INVX1 U8161 (.Y(n10602), 
	.A(\ram[46][1] ));
   OAI22X1 U8162 (.Y(n1318), 
	.B1(n10603), 
	.B0(n10587), 
	.A1(n10586), 
	.A0(n6309));
   INVX1 U8163 (.Y(n10603), 
	.A(\ram[46][0] ));
   NOR2BX1 U8164 (.Y(n10587), 
	.B(n10586), 
	.AN(mem_write_en));
   NAND2X1 U8165 (.Y(n10586), 
	.B(n6553), 
	.A(n10585));
   OAI22X1 U8166 (.Y(n1317), 
	.B1(n10606), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6311));
   INVX1 U8167 (.Y(n10606), 
	.A(\ram[45][15] ));
   OAI22X1 U8168 (.Y(n1316), 
	.B1(n10607), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6314));
   INVX1 U8169 (.Y(n10607), 
	.A(\ram[45][14] ));
   OAI22X1 U8170 (.Y(n1315), 
	.B1(n10608), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6316));
   INVX1 U8171 (.Y(n10608), 
	.A(\ram[45][13] ));
   OAI22X1 U8172 (.Y(n1314), 
	.B1(n10609), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6318));
   INVX1 U8173 (.Y(n10609), 
	.A(\ram[45][12] ));
   OAI22X1 U8174 (.Y(n1313), 
	.B1(n10610), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6320));
   INVX1 U8175 (.Y(n10610), 
	.A(\ram[45][11] ));
   OAI22X1 U8176 (.Y(n1312), 
	.B1(n10611), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6322));
   INVX1 U8177 (.Y(n10611), 
	.A(\ram[45][10] ));
   OAI22X1 U8178 (.Y(n1311), 
	.B1(n10612), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6324));
   INVX1 U8179 (.Y(n10612), 
	.A(\ram[45][9] ));
   OAI22X1 U8180 (.Y(n1310), 
	.B1(n10613), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6326));
   INVX1 U8181 (.Y(n10613), 
	.A(\ram[45][8] ));
   OAI22X1 U8182 (.Y(n1309), 
	.B1(n10614), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6328));
   INVX1 U8183 (.Y(n10614), 
	.A(\ram[45][7] ));
   OAI22X1 U8184 (.Y(n1308), 
	.B1(n10615), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6330));
   INVX1 U8185 (.Y(n10615), 
	.A(\ram[45][6] ));
   OAI22X1 U8186 (.Y(n1307), 
	.B1(n10616), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6332));
   INVX1 U8187 (.Y(n10616), 
	.A(\ram[45][5] ));
   OAI22X1 U8188 (.Y(n1306), 
	.B1(n10617), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6334));
   INVX1 U8189 (.Y(n10617), 
	.A(\ram[45][4] ));
   OAI22X1 U8190 (.Y(n1305), 
	.B1(n10618), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6336));
   INVX1 U8191 (.Y(n10618), 
	.A(\ram[45][3] ));
   OAI22X1 U8192 (.Y(n1304), 
	.B1(n10619), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6338));
   INVX1 U8193 (.Y(n10619), 
	.A(\ram[45][2] ));
   OAI22X1 U8194 (.Y(n1303), 
	.B1(n10620), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6306));
   INVX1 U8195 (.Y(n10620), 
	.A(\ram[45][1] ));
   OAI22X1 U8196 (.Y(n1302), 
	.B1(n10621), 
	.B0(n10605), 
	.A1(n10604), 
	.A0(n6309));
   INVX1 U8197 (.Y(n10621), 
	.A(\ram[45][0] ));
   NOR2BX1 U8198 (.Y(n10605), 
	.B(n10604), 
	.AN(mem_write_en));
   NAND2X1 U8199 (.Y(n10604), 
	.B(n6572), 
	.A(n10585));
   OAI22X1 U8200 (.Y(n1301), 
	.B1(n10624), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6311));
   INVX1 U8201 (.Y(n10624), 
	.A(\ram[44][15] ));
   OAI22X1 U8202 (.Y(n1300), 
	.B1(n10625), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6314));
   INVX1 U8203 (.Y(n10625), 
	.A(\ram[44][14] ));
   OAI22X1 U8204 (.Y(n1299), 
	.B1(n10626), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6316));
   INVX1 U8205 (.Y(n10626), 
	.A(\ram[44][13] ));
   OAI22X1 U8206 (.Y(n1298), 
	.B1(n10627), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6318));
   INVX1 U8207 (.Y(n10627), 
	.A(\ram[44][12] ));
   OAI22X1 U8208 (.Y(n1297), 
	.B1(n10628), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6320));
   INVX1 U8209 (.Y(n10628), 
	.A(\ram[44][11] ));
   OAI22X1 U8210 (.Y(n1296), 
	.B1(n10629), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6322));
   INVX1 U8211 (.Y(n10629), 
	.A(\ram[44][10] ));
   OAI22X1 U8212 (.Y(n1295), 
	.B1(n10630), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6324));
   INVX1 U8213 (.Y(n10630), 
	.A(\ram[44][9] ));
   OAI22X1 U8214 (.Y(n1294), 
	.B1(n10631), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6326));
   INVX1 U8215 (.Y(n10631), 
	.A(\ram[44][8] ));
   OAI22X1 U8216 (.Y(n1293), 
	.B1(n10632), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6328));
   INVX1 U8217 (.Y(n10632), 
	.A(\ram[44][7] ));
   OAI22X1 U8218 (.Y(n1292), 
	.B1(n10633), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6330));
   INVX1 U8219 (.Y(n10633), 
	.A(\ram[44][6] ));
   OAI22X1 U8220 (.Y(n1291), 
	.B1(n10634), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6332));
   INVX1 U8221 (.Y(n10634), 
	.A(\ram[44][5] ));
   OAI22X1 U8222 (.Y(n1290), 
	.B1(n10635), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6334));
   INVX1 U8223 (.Y(n10635), 
	.A(\ram[44][4] ));
   OAI22X1 U8224 (.Y(n1289), 
	.B1(n10636), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6336));
   INVX1 U8225 (.Y(n10636), 
	.A(\ram[44][3] ));
   OAI22X1 U8226 (.Y(n1288), 
	.B1(n10637), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6338));
   INVX1 U8227 (.Y(n10637), 
	.A(\ram[44][2] ));
   OAI22X1 U8228 (.Y(n1287), 
	.B1(n10638), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6306));
   INVX1 U8229 (.Y(n10638), 
	.A(\ram[44][1] ));
   OAI22X1 U8230 (.Y(n1286), 
	.B1(n10639), 
	.B0(n10623), 
	.A1(n10622), 
	.A0(n6309));
   INVX1 U8231 (.Y(n10639), 
	.A(\ram[44][0] ));
   NOR2BX1 U8232 (.Y(n10623), 
	.B(n10622), 
	.AN(mem_write_en));
   NAND2X1 U8233 (.Y(n10622), 
	.B(n6591), 
	.A(n10585));
   OAI22X1 U8234 (.Y(n1285), 
	.B1(n10642), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6311));
   INVX1 U8235 (.Y(n10642), 
	.A(\ram[43][15] ));
   OAI22X1 U8236 (.Y(n1284), 
	.B1(n10643), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6314));
   INVX1 U8237 (.Y(n10643), 
	.A(\ram[43][14] ));
   OAI22X1 U8238 (.Y(n1283), 
	.B1(n10644), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6316));
   INVX1 U8239 (.Y(n10644), 
	.A(\ram[43][13] ));
   OAI22X1 U8240 (.Y(n1282), 
	.B1(n10645), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6318));
   INVX1 U8241 (.Y(n10645), 
	.A(\ram[43][12] ));
   OAI22X1 U8242 (.Y(n1281), 
	.B1(n10646), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6320));
   INVX1 U8243 (.Y(n10646), 
	.A(\ram[43][11] ));
   OAI22X1 U8244 (.Y(n1280), 
	.B1(n10647), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6322));
   INVX1 U8245 (.Y(n10647), 
	.A(\ram[43][10] ));
   OAI22X1 U8246 (.Y(n1279), 
	.B1(n10648), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6324));
   INVX1 U8247 (.Y(n10648), 
	.A(\ram[43][9] ));
   OAI22X1 U8248 (.Y(n1278), 
	.B1(n10649), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6326));
   INVX1 U8249 (.Y(n10649), 
	.A(\ram[43][8] ));
   OAI22X1 U8250 (.Y(n1277), 
	.B1(n10650), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6328));
   INVX1 U8251 (.Y(n10650), 
	.A(\ram[43][7] ));
   OAI22X1 U8252 (.Y(n1276), 
	.B1(n10651), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6330));
   INVX1 U8253 (.Y(n10651), 
	.A(\ram[43][6] ));
   OAI22X1 U8254 (.Y(n1275), 
	.B1(n10652), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6332));
   INVX1 U8255 (.Y(n10652), 
	.A(\ram[43][5] ));
   OAI22X1 U8256 (.Y(n1274), 
	.B1(n10653), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6334));
   INVX1 U8257 (.Y(n10653), 
	.A(\ram[43][4] ));
   OAI22X1 U8258 (.Y(n1273), 
	.B1(n10654), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6336));
   INVX1 U8259 (.Y(n10654), 
	.A(\ram[43][3] ));
   OAI22X1 U8260 (.Y(n1272), 
	.B1(n10655), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6338));
   INVX1 U8261 (.Y(n10655), 
	.A(\ram[43][2] ));
   OAI22X1 U8262 (.Y(n1271), 
	.B1(n10656), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6306));
   INVX1 U8263 (.Y(n10656), 
	.A(\ram[43][1] ));
   OAI22X1 U8264 (.Y(n1270), 
	.B1(n10657), 
	.B0(n10641), 
	.A1(n10640), 
	.A0(n6309));
   INVX1 U8265 (.Y(n10657), 
	.A(\ram[43][0] ));
   NOR2BX1 U8266 (.Y(n10641), 
	.B(n10640), 
	.AN(mem_write_en));
   NAND2X1 U8267 (.Y(n10640), 
	.B(n6610), 
	.A(n10585));
   OAI22X1 U8268 (.Y(n1269), 
	.B1(n10660), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6311));
   INVX1 U8269 (.Y(n10660), 
	.A(\ram[42][15] ));
   OAI22X1 U8270 (.Y(n1268), 
	.B1(n10661), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6314));
   INVX1 U8271 (.Y(n10661), 
	.A(\ram[42][14] ));
   OAI22X1 U8272 (.Y(n1267), 
	.B1(n10662), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6316));
   INVX1 U8273 (.Y(n10662), 
	.A(\ram[42][13] ));
   OAI22X1 U8274 (.Y(n1266), 
	.B1(n10663), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6318));
   INVX1 U8275 (.Y(n10663), 
	.A(\ram[42][12] ));
   OAI22X1 U8276 (.Y(n1265), 
	.B1(n10664), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6320));
   INVX1 U8277 (.Y(n10664), 
	.A(\ram[42][11] ));
   OAI22X1 U8278 (.Y(n1264), 
	.B1(n10665), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6322));
   INVX1 U8279 (.Y(n10665), 
	.A(\ram[42][10] ));
   OAI22X1 U8280 (.Y(n1263), 
	.B1(n10666), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6324));
   INVX1 U8281 (.Y(n10666), 
	.A(\ram[42][9] ));
   OAI22X1 U8282 (.Y(n1262), 
	.B1(n10667), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6326));
   INVX1 U8283 (.Y(n10667), 
	.A(\ram[42][8] ));
   OAI22X1 U8284 (.Y(n1261), 
	.B1(n10668), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6328));
   INVX1 U8285 (.Y(n10668), 
	.A(\ram[42][7] ));
   OAI22X1 U8286 (.Y(n1260), 
	.B1(n10669), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6330));
   INVX1 U8287 (.Y(n10669), 
	.A(\ram[42][6] ));
   OAI22X1 U8288 (.Y(n1259), 
	.B1(n10670), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6332));
   INVX1 U8289 (.Y(n10670), 
	.A(\ram[42][5] ));
   OAI22X1 U8290 (.Y(n1258), 
	.B1(n10671), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6334));
   INVX1 U8291 (.Y(n10671), 
	.A(\ram[42][4] ));
   OAI22X1 U8292 (.Y(n1257), 
	.B1(n10672), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6336));
   INVX1 U8293 (.Y(n10672), 
	.A(\ram[42][3] ));
   OAI22X1 U8294 (.Y(n1256), 
	.B1(n10673), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6338));
   INVX1 U8295 (.Y(n10673), 
	.A(\ram[42][2] ));
   OAI22X1 U8296 (.Y(n1255), 
	.B1(n10674), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6306));
   INVX1 U8297 (.Y(n10674), 
	.A(\ram[42][1] ));
   OAI22X1 U8298 (.Y(n1254), 
	.B1(n10675), 
	.B0(n10659), 
	.A1(n10658), 
	.A0(n6309));
   INVX1 U8299 (.Y(n10675), 
	.A(\ram[42][0] ));
   NOR2BX1 U8300 (.Y(n10659), 
	.B(n10658), 
	.AN(mem_write_en));
   NAND2X1 U8301 (.Y(n10658), 
	.B(n6629), 
	.A(n10585));
   OAI22X1 U8302 (.Y(n1253), 
	.B1(n10678), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6311));
   INVX1 U8303 (.Y(n10678), 
	.A(\ram[41][15] ));
   OAI22X1 U8304 (.Y(n1252), 
	.B1(n10679), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6314));
   INVX1 U8305 (.Y(n10679), 
	.A(\ram[41][14] ));
   OAI22X1 U8306 (.Y(n1251), 
	.B1(n10680), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6316));
   INVX1 U8307 (.Y(n10680), 
	.A(\ram[41][13] ));
   OAI22X1 U8308 (.Y(n1250), 
	.B1(n10681), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6318));
   INVX1 U8309 (.Y(n10681), 
	.A(\ram[41][12] ));
   OAI22X1 U8310 (.Y(n1249), 
	.B1(n10682), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6320));
   INVX1 U8311 (.Y(n10682), 
	.A(\ram[41][11] ));
   OAI22X1 U8312 (.Y(n1248), 
	.B1(n10683), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6322));
   INVX1 U8313 (.Y(n10683), 
	.A(\ram[41][10] ));
   OAI22X1 U8314 (.Y(n1247), 
	.B1(n10684), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6324));
   INVX1 U8315 (.Y(n10684), 
	.A(\ram[41][9] ));
   OAI22X1 U8316 (.Y(n1246), 
	.B1(n10685), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6326));
   INVX1 U8317 (.Y(n10685), 
	.A(\ram[41][8] ));
   OAI22X1 U8318 (.Y(n1245), 
	.B1(n10686), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6328));
   INVX1 U8319 (.Y(n10686), 
	.A(\ram[41][7] ));
   OAI22X1 U8320 (.Y(n1244), 
	.B1(n10687), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6330));
   INVX1 U8321 (.Y(n10687), 
	.A(\ram[41][6] ));
   OAI22X1 U8322 (.Y(n1243), 
	.B1(n10688), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6332));
   INVX1 U8323 (.Y(n10688), 
	.A(\ram[41][5] ));
   OAI22X1 U8324 (.Y(n1242), 
	.B1(n10689), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6334));
   INVX1 U8325 (.Y(n10689), 
	.A(\ram[41][4] ));
   OAI22X1 U8326 (.Y(n1241), 
	.B1(n10690), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6336));
   INVX1 U8327 (.Y(n10690), 
	.A(\ram[41][3] ));
   OAI22X1 U8328 (.Y(n1240), 
	.B1(n10691), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6338));
   INVX1 U8329 (.Y(n10691), 
	.A(\ram[41][2] ));
   OAI22X1 U8330 (.Y(n1239), 
	.B1(n10692), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6306));
   INVX1 U8331 (.Y(n10692), 
	.A(\ram[41][1] ));
   OAI22X1 U8332 (.Y(n1238), 
	.B1(n10693), 
	.B0(n10677), 
	.A1(n10676), 
	.A0(n6309));
   INVX1 U8333 (.Y(n10693), 
	.A(\ram[41][0] ));
   NOR2BX1 U8334 (.Y(n10677), 
	.B(n10676), 
	.AN(mem_write_en));
   NAND2X1 U8335 (.Y(n10676), 
	.B(n6342), 
	.A(n10585));
   OAI22X1 U8336 (.Y(n1237), 
	.B1(n10696), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6311));
   INVX1 U8337 (.Y(n10696), 
	.A(\ram[40][15] ));
   OAI22X1 U8338 (.Y(n1236), 
	.B1(n10697), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6314));
   INVX1 U8339 (.Y(n10697), 
	.A(\ram[40][14] ));
   OAI22X1 U8340 (.Y(n1235), 
	.B1(n10698), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6316));
   INVX1 U8341 (.Y(n10698), 
	.A(\ram[40][13] ));
   OAI22X1 U8342 (.Y(n1234), 
	.B1(n10699), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6318));
   INVX1 U8343 (.Y(n10699), 
	.A(\ram[40][12] ));
   OAI22X1 U8344 (.Y(n1233), 
	.B1(n10700), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6320));
   INVX1 U8345 (.Y(n10700), 
	.A(\ram[40][11] ));
   OAI22X1 U8346 (.Y(n1232), 
	.B1(n10701), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6322));
   INVX1 U8347 (.Y(n10701), 
	.A(\ram[40][10] ));
   OAI22X1 U8348 (.Y(n1231), 
	.B1(n10702), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6324));
   INVX1 U8349 (.Y(n10702), 
	.A(\ram[40][9] ));
   OAI22X1 U8350 (.Y(n1230), 
	.B1(n10703), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6326));
   INVX1 U8351 (.Y(n10703), 
	.A(\ram[40][8] ));
   OAI22X1 U8352 (.Y(n1229), 
	.B1(n10704), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6328));
   INVX1 U8353 (.Y(n10704), 
	.A(\ram[40][7] ));
   OAI22X1 U8354 (.Y(n1228), 
	.B1(n10705), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6330));
   INVX1 U8355 (.Y(n10705), 
	.A(\ram[40][6] ));
   OAI22X1 U8356 (.Y(n1227), 
	.B1(n10706), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6332));
   INVX1 U8357 (.Y(n10706), 
	.A(\ram[40][5] ));
   OAI22X1 U8358 (.Y(n1226), 
	.B1(n10707), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6334));
   INVX1 U8359 (.Y(n10707), 
	.A(\ram[40][4] ));
   OAI22X1 U8360 (.Y(n1225), 
	.B1(n10708), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6336));
   INVX1 U8361 (.Y(n10708), 
	.A(\ram[40][3] ));
   OAI22X1 U8362 (.Y(n1224), 
	.B1(n10709), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6338));
   INVX1 U8363 (.Y(n10709), 
	.A(\ram[40][2] ));
   OAI22X1 U8364 (.Y(n1223), 
	.B1(n10710), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6306));
   INVX1 U8365 (.Y(n10710), 
	.A(\ram[40][1] ));
   OAI22X1 U8366 (.Y(n1222), 
	.B1(n10711), 
	.B0(n10695), 
	.A1(n10694), 
	.A0(n6309));
   INVX1 U8367 (.Y(n10711), 
	.A(\ram[40][0] ));
   NOR2BX1 U8368 (.Y(n10695), 
	.B(n10694), 
	.AN(mem_write_en));
   NAND2X1 U8369 (.Y(n10694), 
	.B(n6362), 
	.A(n10585));
   OAI22X1 U8370 (.Y(n1221), 
	.B1(n10714), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6311));
   INVX1 U8371 (.Y(n10714), 
	.A(\ram[39][15] ));
   OAI22X1 U8372 (.Y(n1220), 
	.B1(n10715), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6314));
   INVX1 U8373 (.Y(n10715), 
	.A(\ram[39][14] ));
   OAI22X1 U8374 (.Y(n1219), 
	.B1(n10716), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6316));
   INVX1 U8375 (.Y(n10716), 
	.A(\ram[39][13] ));
   OAI22X1 U8376 (.Y(n1218), 
	.B1(n10717), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6318));
   INVX1 U8377 (.Y(n10717), 
	.A(\ram[39][12] ));
   OAI22X1 U8378 (.Y(n1217), 
	.B1(n10718), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6320));
   INVX1 U8379 (.Y(n10718), 
	.A(\ram[39][11] ));
   OAI22X1 U8380 (.Y(n1216), 
	.B1(n10719), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6322));
   INVX1 U8381 (.Y(n10719), 
	.A(\ram[39][10] ));
   OAI22X1 U8382 (.Y(n1215), 
	.B1(n10720), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6324));
   INVX1 U8383 (.Y(n10720), 
	.A(\ram[39][9] ));
   OAI22X1 U8384 (.Y(n1214), 
	.B1(n10721), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6326));
   INVX1 U8385 (.Y(n10721), 
	.A(\ram[39][8] ));
   OAI22X1 U8386 (.Y(n1213), 
	.B1(n10722), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6328));
   INVX1 U8387 (.Y(n10722), 
	.A(\ram[39][7] ));
   OAI22X1 U8388 (.Y(n1212), 
	.B1(n10723), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6330));
   INVX1 U8389 (.Y(n10723), 
	.A(\ram[39][6] ));
   OAI22X1 U8390 (.Y(n1211), 
	.B1(n10724), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6332));
   INVX1 U8391 (.Y(n10724), 
	.A(\ram[39][5] ));
   OAI22X1 U8392 (.Y(n1210), 
	.B1(n10725), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6334));
   INVX1 U8393 (.Y(n10725), 
	.A(\ram[39][4] ));
   OAI22X1 U8394 (.Y(n1209), 
	.B1(n10726), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6336));
   INVX1 U8395 (.Y(n10726), 
	.A(\ram[39][3] ));
   OAI22X1 U8396 (.Y(n1208), 
	.B1(n10727), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6338));
   INVX1 U8397 (.Y(n10727), 
	.A(\ram[39][2] ));
   OAI22X1 U8398 (.Y(n1207), 
	.B1(n10728), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6306));
   INVX1 U8399 (.Y(n10728), 
	.A(\ram[39][1] ));
   OAI22X1 U8400 (.Y(n1206), 
	.B1(n10729), 
	.B0(n10713), 
	.A1(n10712), 
	.A0(n6309));
   INVX1 U8401 (.Y(n10729), 
	.A(\ram[39][0] ));
   NOR2BX1 U8402 (.Y(n10713), 
	.B(n10712), 
	.AN(mem_write_en));
   NAND2X1 U8403 (.Y(n10712), 
	.B(n6381), 
	.A(n10585));
   OAI22X1 U8404 (.Y(n1205), 
	.B1(n10732), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6311));
   INVX1 U8405 (.Y(n10732), 
	.A(\ram[38][15] ));
   OAI22X1 U8406 (.Y(n1204), 
	.B1(n10733), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6314));
   INVX1 U8407 (.Y(n10733), 
	.A(\ram[38][14] ));
   OAI22X1 U8408 (.Y(n1203), 
	.B1(n10734), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6316));
   INVX1 U8409 (.Y(n10734), 
	.A(\ram[38][13] ));
   OAI22X1 U8410 (.Y(n1202), 
	.B1(n10735), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6318));
   INVX1 U8411 (.Y(n10735), 
	.A(\ram[38][12] ));
   OAI22X1 U8412 (.Y(n1201), 
	.B1(n10736), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6320));
   INVX1 U8413 (.Y(n10736), 
	.A(\ram[38][11] ));
   OAI22X1 U8414 (.Y(n1200), 
	.B1(n10737), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6322));
   INVX1 U8415 (.Y(n10737), 
	.A(\ram[38][10] ));
   OAI22X1 U8416 (.Y(n1199), 
	.B1(n10738), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6324));
   INVX1 U8417 (.Y(n10738), 
	.A(\ram[38][9] ));
   OAI22X1 U8418 (.Y(n1198), 
	.B1(n10739), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6326));
   INVX1 U8419 (.Y(n10739), 
	.A(\ram[38][8] ));
   OAI22X1 U8420 (.Y(n1197), 
	.B1(n10740), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6328));
   INVX1 U8421 (.Y(n10740), 
	.A(\ram[38][7] ));
   OAI22X1 U8422 (.Y(n1196), 
	.B1(n10741), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6330));
   INVX1 U8423 (.Y(n10741), 
	.A(\ram[38][6] ));
   OAI22X1 U8424 (.Y(n1195), 
	.B1(n10742), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6332));
   INVX1 U8425 (.Y(n10742), 
	.A(\ram[38][5] ));
   OAI22X1 U8426 (.Y(n1194), 
	.B1(n10743), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6334));
   INVX1 U8427 (.Y(n10743), 
	.A(\ram[38][4] ));
   OAI22X1 U8428 (.Y(n1193), 
	.B1(n10744), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6336));
   INVX1 U8429 (.Y(n10744), 
	.A(\ram[38][3] ));
   OAI22X1 U8430 (.Y(n1192), 
	.B1(n10745), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6338));
   INVX1 U8431 (.Y(n10745), 
	.A(\ram[38][2] ));
   OAI22X1 U8432 (.Y(n1191), 
	.B1(n10746), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6306));
   INVX1 U8433 (.Y(n10746), 
	.A(\ram[38][1] ));
   OAI22X1 U8434 (.Y(n1190), 
	.B1(n10747), 
	.B0(n10731), 
	.A1(n10730), 
	.A0(n6309));
   INVX1 U8435 (.Y(n10747), 
	.A(\ram[38][0] ));
   NOR2BX1 U8436 (.Y(n10731), 
	.B(n10730), 
	.AN(mem_write_en));
   NAND2X1 U8437 (.Y(n10730), 
	.B(n6400), 
	.A(n10585));
   OAI22X1 U8438 (.Y(n1189), 
	.B1(n10750), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6311));
   INVX1 U8439 (.Y(n10750), 
	.A(\ram[37][15] ));
   OAI22X1 U8440 (.Y(n1188), 
	.B1(n10751), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6314));
   INVX1 U8441 (.Y(n10751), 
	.A(\ram[37][14] ));
   OAI22X1 U8442 (.Y(n1187), 
	.B1(n10752), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6316));
   INVX1 U8443 (.Y(n10752), 
	.A(\ram[37][13] ));
   OAI22X1 U8444 (.Y(n1186), 
	.B1(n10753), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6318));
   INVX1 U8445 (.Y(n10753), 
	.A(\ram[37][12] ));
   OAI22X1 U8446 (.Y(n1185), 
	.B1(n10754), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6320));
   INVX1 U8447 (.Y(n10754), 
	.A(\ram[37][11] ));
   OAI22X1 U8448 (.Y(n1184), 
	.B1(n10755), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6322));
   INVX1 U8449 (.Y(n10755), 
	.A(\ram[37][10] ));
   OAI22X1 U8450 (.Y(n1183), 
	.B1(n10756), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6324));
   INVX1 U8451 (.Y(n10756), 
	.A(\ram[37][9] ));
   OAI22X1 U8452 (.Y(n1182), 
	.B1(n10757), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6326));
   INVX1 U8453 (.Y(n10757), 
	.A(\ram[37][8] ));
   OAI22X1 U8454 (.Y(n1181), 
	.B1(n10758), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6328));
   INVX1 U8455 (.Y(n10758), 
	.A(\ram[37][7] ));
   OAI22X1 U8456 (.Y(n1180), 
	.B1(n10759), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6330));
   INVX1 U8457 (.Y(n10759), 
	.A(\ram[37][6] ));
   OAI22X1 U8458 (.Y(n1179), 
	.B1(n10760), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6332));
   INVX1 U8459 (.Y(n10760), 
	.A(\ram[37][5] ));
   OAI22X1 U8460 (.Y(n1178), 
	.B1(n10761), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6334));
   INVX1 U8461 (.Y(n10761), 
	.A(\ram[37][4] ));
   OAI22X1 U8462 (.Y(n1177), 
	.B1(n10762), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6336));
   INVX1 U8463 (.Y(n10762), 
	.A(\ram[37][3] ));
   OAI22X1 U8464 (.Y(n1176), 
	.B1(n10763), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6338));
   INVX1 U8465 (.Y(n10763), 
	.A(\ram[37][2] ));
   OAI22X1 U8466 (.Y(n1175), 
	.B1(n10764), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6306));
   INVX1 U8467 (.Y(n10764), 
	.A(\ram[37][1] ));
   OAI22X1 U8468 (.Y(n1174), 
	.B1(n10765), 
	.B0(n10749), 
	.A1(n10748), 
	.A0(n6309));
   INVX1 U8469 (.Y(n10765), 
	.A(\ram[37][0] ));
   NOR2BX1 U8470 (.Y(n10749), 
	.B(n10748), 
	.AN(mem_write_en));
   NAND2X1 U8471 (.Y(n10748), 
	.B(n6419), 
	.A(n10585));
   OAI22X1 U8472 (.Y(n1173), 
	.B1(n10768), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6311));
   INVX1 U8473 (.Y(n10768), 
	.A(\ram[36][15] ));
   OAI22X1 U8474 (.Y(n1172), 
	.B1(n10769), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6314));
   INVX1 U8475 (.Y(n10769), 
	.A(\ram[36][14] ));
   OAI22X1 U8476 (.Y(n1171), 
	.B1(n10770), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6316));
   INVX1 U8477 (.Y(n10770), 
	.A(\ram[36][13] ));
   OAI22X1 U8478 (.Y(n1170), 
	.B1(n10771), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6318));
   INVX1 U8479 (.Y(n10771), 
	.A(\ram[36][12] ));
   OAI22X1 U8480 (.Y(n1169), 
	.B1(n10772), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6320));
   INVX1 U8481 (.Y(n10772), 
	.A(\ram[36][11] ));
   OAI22X1 U8482 (.Y(n1168), 
	.B1(n10773), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6322));
   INVX1 U8483 (.Y(n10773), 
	.A(\ram[36][10] ));
   OAI22X1 U8484 (.Y(n1167), 
	.B1(n10774), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6324));
   INVX1 U8485 (.Y(n10774), 
	.A(\ram[36][9] ));
   OAI22X1 U8486 (.Y(n1166), 
	.B1(n10775), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6326));
   INVX1 U8487 (.Y(n10775), 
	.A(\ram[36][8] ));
   OAI22X1 U8488 (.Y(n1165), 
	.B1(n10776), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6328));
   INVX1 U8489 (.Y(n10776), 
	.A(\ram[36][7] ));
   OAI22X1 U8490 (.Y(n1164), 
	.B1(n10777), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6330));
   INVX1 U8491 (.Y(n10777), 
	.A(\ram[36][6] ));
   OAI22X1 U8492 (.Y(n1163), 
	.B1(n10778), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6332));
   INVX1 U8493 (.Y(n10778), 
	.A(\ram[36][5] ));
   OAI22X1 U8494 (.Y(n1162), 
	.B1(n10779), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6334));
   INVX1 U8495 (.Y(n10779), 
	.A(\ram[36][4] ));
   OAI22X1 U8496 (.Y(n1161), 
	.B1(n10780), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6336));
   INVX1 U8497 (.Y(n10780), 
	.A(\ram[36][3] ));
   OAI22X1 U8498 (.Y(n1160), 
	.B1(n10781), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6338));
   INVX1 U8499 (.Y(n10781), 
	.A(\ram[36][2] ));
   OAI22X1 U8500 (.Y(n1159), 
	.B1(n10782), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6306));
   INVX1 U8501 (.Y(n10782), 
	.A(\ram[36][1] ));
   OAI22X1 U8502 (.Y(n1158), 
	.B1(n10783), 
	.B0(n10767), 
	.A1(n10766), 
	.A0(n6309));
   INVX1 U8503 (.Y(n10783), 
	.A(\ram[36][0] ));
   NOR2BX1 U8504 (.Y(n10767), 
	.B(n10766), 
	.AN(mem_write_en));
   NAND2X1 U8505 (.Y(n10766), 
	.B(n6438), 
	.A(n10585));
   OAI22X1 U8506 (.Y(n1157), 
	.B1(n10786), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6311));
   INVX1 U8507 (.Y(n10786), 
	.A(\ram[35][15] ));
   OAI22X1 U8508 (.Y(n1156), 
	.B1(n10787), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6314));
   INVX1 U8509 (.Y(n10787), 
	.A(\ram[35][14] ));
   OAI22X1 U8510 (.Y(n1155), 
	.B1(n10788), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6316));
   INVX1 U8511 (.Y(n10788), 
	.A(\ram[35][13] ));
   OAI22X1 U8512 (.Y(n1154), 
	.B1(n10789), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6318));
   INVX1 U8513 (.Y(n10789), 
	.A(\ram[35][12] ));
   OAI22X1 U8514 (.Y(n1153), 
	.B1(n10790), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6320));
   INVX1 U8515 (.Y(n10790), 
	.A(\ram[35][11] ));
   OAI22X1 U8516 (.Y(n1152), 
	.B1(n10791), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6322));
   INVX1 U8517 (.Y(n10791), 
	.A(\ram[35][10] ));
   OAI22X1 U8518 (.Y(n1151), 
	.B1(n10792), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6324));
   INVX1 U8519 (.Y(n10792), 
	.A(\ram[35][9] ));
   OAI22X1 U8520 (.Y(n1150), 
	.B1(n10793), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6326));
   INVX1 U8521 (.Y(n10793), 
	.A(\ram[35][8] ));
   OAI22X1 U8522 (.Y(n1149), 
	.B1(n10794), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6328));
   INVX1 U8523 (.Y(n10794), 
	.A(\ram[35][7] ));
   OAI22X1 U8524 (.Y(n1148), 
	.B1(n10795), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6330));
   INVX1 U8525 (.Y(n10795), 
	.A(\ram[35][6] ));
   OAI22X1 U8526 (.Y(n1147), 
	.B1(n10796), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6332));
   INVX1 U8527 (.Y(n10796), 
	.A(\ram[35][5] ));
   OAI22X1 U8528 (.Y(n1146), 
	.B1(n10797), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6334));
   INVX1 U8529 (.Y(n10797), 
	.A(\ram[35][4] ));
   OAI22X1 U8530 (.Y(n1145), 
	.B1(n10798), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6336));
   INVX1 U8531 (.Y(n10798), 
	.A(\ram[35][3] ));
   OAI22X1 U8532 (.Y(n1144), 
	.B1(n10799), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6338));
   INVX1 U8533 (.Y(n10799), 
	.A(\ram[35][2] ));
   OAI22X1 U8534 (.Y(n1143), 
	.B1(n10800), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6306));
   INVX1 U8535 (.Y(n10800), 
	.A(\ram[35][1] ));
   OAI22X1 U8536 (.Y(n1142), 
	.B1(n10801), 
	.B0(n10785), 
	.A1(n10784), 
	.A0(n6309));
   INVX1 U8537 (.Y(n10801), 
	.A(\ram[35][0] ));
   NOR2BX1 U8538 (.Y(n10785), 
	.B(n10784), 
	.AN(mem_write_en));
   NAND2X1 U8539 (.Y(n10784), 
	.B(n6457), 
	.A(n10585));
   OAI22X1 U8540 (.Y(n1141), 
	.B1(n10804), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6311));
   INVX1 U8541 (.Y(n10804), 
	.A(\ram[34][15] ));
   OAI22X1 U8542 (.Y(n1140), 
	.B1(n10805), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6314));
   INVX1 U8543 (.Y(n10805), 
	.A(\ram[34][14] ));
   OAI22X1 U8544 (.Y(n1139), 
	.B1(n10806), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6316));
   INVX1 U8545 (.Y(n10806), 
	.A(\ram[34][13] ));
   OAI22X1 U8546 (.Y(n1138), 
	.B1(n10807), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6318));
   INVX1 U8547 (.Y(n10807), 
	.A(\ram[34][12] ));
   OAI22X1 U8548 (.Y(n1137), 
	.B1(n10808), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6320));
   INVX1 U8549 (.Y(n10808), 
	.A(\ram[34][11] ));
   OAI22X1 U8550 (.Y(n1136), 
	.B1(n10809), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6322));
   INVX1 U8551 (.Y(n10809), 
	.A(\ram[34][10] ));
   OAI22X1 U8552 (.Y(n1135), 
	.B1(n10810), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6324));
   INVX1 U8553 (.Y(n10810), 
	.A(\ram[34][9] ));
   OAI22X1 U8554 (.Y(n1134), 
	.B1(n10811), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6326));
   INVX1 U8555 (.Y(n10811), 
	.A(\ram[34][8] ));
   OAI22X1 U8556 (.Y(n1133), 
	.B1(n10812), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6328));
   INVX1 U8557 (.Y(n10812), 
	.A(\ram[34][7] ));
   OAI22X1 U8558 (.Y(n1132), 
	.B1(n10813), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6330));
   INVX1 U8559 (.Y(n10813), 
	.A(\ram[34][6] ));
   OAI22X1 U8560 (.Y(n1131), 
	.B1(n10814), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6332));
   INVX1 U8561 (.Y(n10814), 
	.A(\ram[34][5] ));
   OAI22X1 U8562 (.Y(n1130), 
	.B1(n10815), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6334));
   INVX1 U8563 (.Y(n10815), 
	.A(\ram[34][4] ));
   OAI22X1 U8564 (.Y(n1129), 
	.B1(n10816), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6336));
   INVX1 U8565 (.Y(n10816), 
	.A(\ram[34][3] ));
   OAI22X1 U8566 (.Y(n1128), 
	.B1(n10817), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6338));
   INVX1 U8567 (.Y(n10817), 
	.A(\ram[34][2] ));
   OAI22X1 U8568 (.Y(n1127), 
	.B1(n10818), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6306));
   INVX1 U8569 (.Y(n10818), 
	.A(\ram[34][1] ));
   OAI22X1 U8570 (.Y(n1126), 
	.B1(n10819), 
	.B0(n10803), 
	.A1(n10802), 
	.A0(n6309));
   INVX1 U8571 (.Y(n10819), 
	.A(\ram[34][0] ));
   NOR2BX1 U8572 (.Y(n10803), 
	.B(n10802), 
	.AN(mem_write_en));
   NAND2X1 U8573 (.Y(n10802), 
	.B(n6476), 
	.A(n10585));
   OAI22X1 U8574 (.Y(n1125), 
	.B1(n10822), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6311));
   INVX1 U8575 (.Y(n10822), 
	.A(\ram[33][15] ));
   OAI22X1 U8576 (.Y(n1124), 
	.B1(n10823), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6314));
   INVX1 U8577 (.Y(n10823), 
	.A(\ram[33][14] ));
   OAI22X1 U8578 (.Y(n1123), 
	.B1(n10824), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6316));
   INVX1 U8579 (.Y(n10824), 
	.A(\ram[33][13] ));
   OAI22X1 U8580 (.Y(n1122), 
	.B1(n10825), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6318));
   INVX1 U8581 (.Y(n10825), 
	.A(\ram[33][12] ));
   OAI22X1 U8582 (.Y(n1121), 
	.B1(n10826), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6320));
   INVX1 U8583 (.Y(n10826), 
	.A(\ram[33][11] ));
   OAI22X1 U8584 (.Y(n1120), 
	.B1(n10827), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6322));
   INVX1 U8585 (.Y(n10827), 
	.A(\ram[33][10] ));
   OAI22X1 U8586 (.Y(n1119), 
	.B1(n10828), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6324));
   INVX1 U8587 (.Y(n10828), 
	.A(\ram[33][9] ));
   OAI22X1 U8588 (.Y(n1118), 
	.B1(n10829), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6326));
   INVX1 U8589 (.Y(n10829), 
	.A(\ram[33][8] ));
   OAI22X1 U8590 (.Y(n1117), 
	.B1(n10830), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6328));
   INVX1 U8591 (.Y(n10830), 
	.A(\ram[33][7] ));
   OAI22X1 U8592 (.Y(n1116), 
	.B1(n10831), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6330));
   INVX1 U8593 (.Y(n10831), 
	.A(\ram[33][6] ));
   OAI22X1 U8594 (.Y(n1115), 
	.B1(n10832), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6332));
   INVX1 U8595 (.Y(n10832), 
	.A(\ram[33][5] ));
   OAI22X1 U8596 (.Y(n1114), 
	.B1(n10833), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6334));
   INVX1 U8597 (.Y(n10833), 
	.A(\ram[33][4] ));
   OAI22X1 U8598 (.Y(n1113), 
	.B1(n10834), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6336));
   INVX1 U8599 (.Y(n10834), 
	.A(\ram[33][3] ));
   OAI22X1 U8600 (.Y(n1112), 
	.B1(n10835), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6338));
   INVX1 U8601 (.Y(n10835), 
	.A(\ram[33][2] ));
   OAI22X1 U8602 (.Y(n1111), 
	.B1(n10836), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6306));
   INVX1 U8603 (.Y(n10836), 
	.A(\ram[33][1] ));
   OAI22X1 U8604 (.Y(n1110), 
	.B1(n10837), 
	.B0(n10821), 
	.A1(n10820), 
	.A0(n6309));
   INVX1 U8605 (.Y(n10837), 
	.A(\ram[33][0] ));
   NOR2BX1 U8606 (.Y(n10821), 
	.B(n10820), 
	.AN(mem_write_en));
   NAND2X1 U8607 (.Y(n10820), 
	.B(n6495), 
	.A(n10585));
   OAI22X1 U8608 (.Y(n1109), 
	.B1(n10840), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6311));
   INVX1 U8609 (.Y(n10840), 
	.A(\ram[32][15] ));
   OAI22X1 U8610 (.Y(n1108), 
	.B1(n10841), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6314));
   INVX1 U8611 (.Y(n10841), 
	.A(\ram[32][14] ));
   OAI22X1 U8612 (.Y(n1107), 
	.B1(n10842), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6316));
   INVX1 U8613 (.Y(n10842), 
	.A(\ram[32][13] ));
   OAI22X1 U8614 (.Y(n1106), 
	.B1(n10843), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6318));
   INVX1 U8615 (.Y(n10843), 
	.A(\ram[32][12] ));
   OAI22X1 U8616 (.Y(n1105), 
	.B1(n10844), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6320));
   INVX1 U8617 (.Y(n10844), 
	.A(\ram[32][11] ));
   OAI22X1 U8618 (.Y(n1104), 
	.B1(n10845), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6322));
   INVX1 U8619 (.Y(n10845), 
	.A(\ram[32][10] ));
   OAI22X1 U8620 (.Y(n1103), 
	.B1(n10846), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6324));
   INVX1 U8621 (.Y(n10846), 
	.A(\ram[32][9] ));
   OAI22X1 U8622 (.Y(n1102), 
	.B1(n10847), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6326));
   INVX1 U8623 (.Y(n10847), 
	.A(\ram[32][8] ));
   OAI22X1 U8624 (.Y(n1101), 
	.B1(n10848), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6328));
   INVX1 U8625 (.Y(n10848), 
	.A(\ram[32][7] ));
   OAI22X1 U8626 (.Y(n1100), 
	.B1(n10849), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6330));
   INVX1 U8627 (.Y(n10849), 
	.A(\ram[32][6] ));
   OAI22X1 U8628 (.Y(n1099), 
	.B1(n10850), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6332));
   INVX1 U8629 (.Y(n10850), 
	.A(\ram[32][5] ));
   OAI22X1 U8630 (.Y(n1098), 
	.B1(n10851), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6334));
   INVX1 U8631 (.Y(n10851), 
	.A(\ram[32][4] ));
   OAI22X1 U8632 (.Y(n1097), 
	.B1(n10852), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6336));
   INVX1 U8633 (.Y(n10852), 
	.A(\ram[32][3] ));
   OAI22X1 U8634 (.Y(n1096), 
	.B1(n10853), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6338));
   INVX1 U8635 (.Y(n10853), 
	.A(\ram[32][2] ));
   OAI22X1 U8636 (.Y(n1095), 
	.B1(n10854), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6306));
   INVX1 U8637 (.Y(n10854), 
	.A(\ram[32][1] ));
   OAI22X1 U8638 (.Y(n1094), 
	.B1(n10855), 
	.B0(n10839), 
	.A1(n10838), 
	.A0(n6309));
   INVX1 U8639 (.Y(n10855), 
	.A(\ram[32][0] ));
   NOR2BX1 U8640 (.Y(n10839), 
	.B(n10838), 
	.AN(mem_write_en));
   NAND2X1 U8641 (.Y(n10838), 
	.B(n6514), 
	.A(n10585));
   OAI22X1 U8642 (.Y(n1093), 
	.B1(n10858), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6311));
   INVX1 U8643 (.Y(n10858), 
	.A(\ram[31][15] ));
   OAI22X1 U8644 (.Y(n1092), 
	.B1(n10859), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6314));
   INVX1 U8645 (.Y(n10859), 
	.A(\ram[31][14] ));
   OAI22X1 U8646 (.Y(n1091), 
	.B1(n10860), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6316));
   INVX1 U8647 (.Y(n10860), 
	.A(\ram[31][13] ));
   OAI22X1 U8648 (.Y(n1090), 
	.B1(n10861), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6318));
   INVX1 U8649 (.Y(n10861), 
	.A(\ram[31][12] ));
   OAI22X1 U8650 (.Y(n1089), 
	.B1(n10862), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6320));
   INVX1 U8651 (.Y(n10862), 
	.A(\ram[31][11] ));
   OAI22X1 U8652 (.Y(n1088), 
	.B1(n10863), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6322));
   INVX1 U8653 (.Y(n10863), 
	.A(\ram[31][10] ));
   OAI22X1 U8654 (.Y(n1087), 
	.B1(n10864), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6324));
   INVX1 U8655 (.Y(n10864), 
	.A(\ram[31][9] ));
   OAI22X1 U8656 (.Y(n1086), 
	.B1(n10865), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6326));
   INVX1 U8657 (.Y(n10865), 
	.A(\ram[31][8] ));
   OAI22X1 U8658 (.Y(n1085), 
	.B1(n10866), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6328));
   INVX1 U8659 (.Y(n10866), 
	.A(\ram[31][7] ));
   OAI22X1 U8660 (.Y(n1084), 
	.B1(n10867), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6330));
   INVX1 U8661 (.Y(n10867), 
	.A(\ram[31][6] ));
   OAI22X1 U8662 (.Y(n1083), 
	.B1(n10868), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6332));
   INVX1 U8663 (.Y(n10868), 
	.A(\ram[31][5] ));
   OAI22X1 U8664 (.Y(n1082), 
	.B1(n10869), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6334));
   INVX1 U8665 (.Y(n10869), 
	.A(\ram[31][4] ));
   OAI22X1 U8666 (.Y(n1081), 
	.B1(n10870), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6336));
   INVX1 U8667 (.Y(n10870), 
	.A(\ram[31][3] ));
   OAI22X1 U8668 (.Y(n1080), 
	.B1(n10871), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6338));
   INVX1 U8669 (.Y(n10871), 
	.A(\ram[31][2] ));
   OAI22X1 U8670 (.Y(n1079), 
	.B1(n10872), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6306));
   INVX1 U8671 (.Y(n10872), 
	.A(\ram[31][1] ));
   OAI22X1 U8672 (.Y(n1078), 
	.B1(n10873), 
	.B0(n10857), 
	.A1(n10856), 
	.A0(n6309));
   INVX1 U8673 (.Y(n10873), 
	.A(\ram[31][0] ));
   NOR2BX1 U8674 (.Y(n10857), 
	.B(n10856), 
	.AN(mem_write_en));
   NAND2X1 U8675 (.Y(n10856), 
	.B(n6343), 
	.A(n6533));
   OAI22X1 U8676 (.Y(n1077), 
	.B1(n10876), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6311));
   INVX1 U8677 (.Y(n10876), 
	.A(\ram[30][15] ));
   OAI22X1 U8678 (.Y(n1076), 
	.B1(n10877), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6314));
   INVX1 U8679 (.Y(n10877), 
	.A(\ram[30][14] ));
   OAI22X1 U8680 (.Y(n1075), 
	.B1(n10878), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6316));
   INVX1 U8681 (.Y(n10878), 
	.A(\ram[30][13] ));
   OAI22X1 U8682 (.Y(n1074), 
	.B1(n10879), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6318));
   INVX1 U8683 (.Y(n10879), 
	.A(\ram[30][12] ));
   OAI22X1 U8684 (.Y(n1073), 
	.B1(n10880), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6320));
   INVX1 U8685 (.Y(n10880), 
	.A(\ram[30][11] ));
   OAI22X1 U8686 (.Y(n1072), 
	.B1(n10881), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6322));
   INVX1 U8687 (.Y(n10881), 
	.A(\ram[30][10] ));
   OAI22X1 U8688 (.Y(n1071), 
	.B1(n10882), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6324));
   INVX1 U8689 (.Y(n10882), 
	.A(\ram[30][9] ));
   OAI22X1 U8690 (.Y(n1070), 
	.B1(n10883), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6326));
   INVX1 U8691 (.Y(n10883), 
	.A(\ram[30][8] ));
   OAI22X1 U8692 (.Y(n1069), 
	.B1(n10884), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6328));
   INVX1 U8693 (.Y(n10884), 
	.A(\ram[30][7] ));
   OAI22X1 U8694 (.Y(n1068), 
	.B1(n10885), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6330));
   INVX1 U8695 (.Y(n10885), 
	.A(\ram[30][6] ));
   OAI22X1 U8696 (.Y(n1067), 
	.B1(n10886), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6332));
   INVX1 U8697 (.Y(n10886), 
	.A(\ram[30][5] ));
   OAI22X1 U8698 (.Y(n1066), 
	.B1(n10887), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6334));
   INVX1 U8699 (.Y(n10887), 
	.A(\ram[30][4] ));
   OAI22X1 U8700 (.Y(n1065), 
	.B1(n10888), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6336));
   INVX1 U8701 (.Y(n10888), 
	.A(\ram[30][3] ));
   OAI22X1 U8702 (.Y(n1064), 
	.B1(n10889), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6338));
   INVX1 U8703 (.Y(n10889), 
	.A(\ram[30][2] ));
   OAI22X1 U8704 (.Y(n1063), 
	.B1(n10890), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6306));
   INVX1 U8705 (.Y(n10890), 
	.A(\ram[30][1] ));
   OAI22X1 U8706 (.Y(n1062), 
	.B1(n10891), 
	.B0(n10875), 
	.A1(n10874), 
	.A0(n6309));
   INVX1 U8707 (.Y(n10891), 
	.A(\ram[30][0] ));
   NOR2BX1 U8708 (.Y(n10875), 
	.B(n10874), 
	.AN(mem_write_en));
   NAND2X1 U8709 (.Y(n10874), 
	.B(n6343), 
	.A(n6553));
   OAI22X1 U8710 (.Y(n1061), 
	.B1(n10894), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6311));
   INVX1 U8711 (.Y(n10894), 
	.A(\ram[29][15] ));
   OAI22X1 U8712 (.Y(n1060), 
	.B1(n10895), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6314));
   INVX1 U8713 (.Y(n10895), 
	.A(\ram[29][14] ));
   OAI22X1 U8714 (.Y(n1059), 
	.B1(n10896), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6316));
   INVX1 U8715 (.Y(n10896), 
	.A(\ram[29][13] ));
   OAI22X1 U8716 (.Y(n1058), 
	.B1(n10897), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6318));
   INVX1 U8717 (.Y(n10897), 
	.A(\ram[29][12] ));
   OAI22X1 U8718 (.Y(n1057), 
	.B1(n10898), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6320));
   INVX1 U8719 (.Y(n10898), 
	.A(\ram[29][11] ));
   OAI22X1 U8720 (.Y(n1056), 
	.B1(n10899), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6322));
   INVX1 U8721 (.Y(n10899), 
	.A(\ram[29][10] ));
   OAI22X1 U8722 (.Y(n1055), 
	.B1(n10900), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6324));
   INVX1 U8723 (.Y(n10900), 
	.A(\ram[29][9] ));
   OAI22X1 U8724 (.Y(n1054), 
	.B1(n10901), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6326));
   INVX1 U8725 (.Y(n10901), 
	.A(\ram[29][8] ));
   OAI22X1 U8726 (.Y(n1053), 
	.B1(n10902), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6328));
   INVX1 U8727 (.Y(n10902), 
	.A(\ram[29][7] ));
   OAI22X1 U8728 (.Y(n1052), 
	.B1(n10903), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6330));
   INVX1 U8729 (.Y(n10903), 
	.A(\ram[29][6] ));
   OAI22X1 U8730 (.Y(n1051), 
	.B1(n10904), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6332));
   INVX1 U8731 (.Y(n10904), 
	.A(\ram[29][5] ));
   OAI22X1 U8732 (.Y(n1050), 
	.B1(n10905), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6334));
   INVX1 U8733 (.Y(n10905), 
	.A(\ram[29][4] ));
   OAI22X1 U8734 (.Y(n1049), 
	.B1(n10906), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6336));
   INVX1 U8735 (.Y(n10906), 
	.A(\ram[29][3] ));
   OAI22X1 U8736 (.Y(n1048), 
	.B1(n10907), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6338));
   INVX1 U8737 (.Y(n10907), 
	.A(\ram[29][2] ));
   OAI22X1 U8738 (.Y(n1047), 
	.B1(n10908), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6306));
   INVX1 U8739 (.Y(n10908), 
	.A(\ram[29][1] ));
   OAI22X1 U8740 (.Y(n1046), 
	.B1(n10909), 
	.B0(n10893), 
	.A1(n10892), 
	.A0(n6309));
   INVX1 U8741 (.Y(n10909), 
	.A(\ram[29][0] ));
   NOR2BX1 U8742 (.Y(n10893), 
	.B(n10892), 
	.AN(mem_write_en));
   NAND2X1 U8743 (.Y(n10892), 
	.B(n6343), 
	.A(n6572));
   OAI22X1 U8744 (.Y(n1045), 
	.B1(n10912), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6311));
   INVX1 U8745 (.Y(n10912), 
	.A(\ram[28][15] ));
   OAI22X1 U8746 (.Y(n1044), 
	.B1(n10913), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6314));
   INVX1 U8747 (.Y(n10913), 
	.A(\ram[28][14] ));
   OAI22X1 U8748 (.Y(n1043), 
	.B1(n10914), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6316));
   INVX1 U8749 (.Y(n10914), 
	.A(\ram[28][13] ));
   OAI22X1 U8750 (.Y(n1042), 
	.B1(n10915), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6318));
   INVX1 U8751 (.Y(n10915), 
	.A(\ram[28][12] ));
   OAI22X1 U8752 (.Y(n1041), 
	.B1(n10916), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6320));
   INVX1 U8753 (.Y(n10916), 
	.A(\ram[28][11] ));
   OAI22X1 U8754 (.Y(n1040), 
	.B1(n10917), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6322));
   INVX1 U8755 (.Y(n10917), 
	.A(\ram[28][10] ));
   OAI22X1 U8756 (.Y(n1039), 
	.B1(n10918), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6324));
   INVX1 U8757 (.Y(n10918), 
	.A(\ram[28][9] ));
   OAI22X1 U8758 (.Y(n1038), 
	.B1(n10919), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6326));
   INVX1 U8759 (.Y(n10919), 
	.A(\ram[28][8] ));
   OAI22X1 U8760 (.Y(n1037), 
	.B1(n10920), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6328));
   INVX1 U8761 (.Y(n10920), 
	.A(\ram[28][7] ));
   OAI22X1 U8762 (.Y(n1036), 
	.B1(n10921), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6330));
   INVX1 U8763 (.Y(n10921), 
	.A(\ram[28][6] ));
   OAI22X1 U8764 (.Y(n1035), 
	.B1(n10922), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6332));
   INVX1 U8765 (.Y(n10922), 
	.A(\ram[28][5] ));
   OAI22X1 U8766 (.Y(n1034), 
	.B1(n10923), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6334));
   INVX1 U8767 (.Y(n10923), 
	.A(\ram[28][4] ));
   OAI22X1 U8768 (.Y(n1033), 
	.B1(n10924), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6336));
   INVX1 U8769 (.Y(n10924), 
	.A(\ram[28][3] ));
   OAI22X1 U8770 (.Y(n1032), 
	.B1(n10925), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6338));
   INVX1 U8771 (.Y(n10925), 
	.A(\ram[28][2] ));
   OAI22X1 U8772 (.Y(n1031), 
	.B1(n10926), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6306));
   INVX1 U8773 (.Y(n10926), 
	.A(\ram[28][1] ));
   OAI22X1 U8774 (.Y(n1030), 
	.B1(n10927), 
	.B0(n10911), 
	.A1(n10910), 
	.A0(n6309));
   INVX1 U8775 (.Y(n10927), 
	.A(\ram[28][0] ));
   NOR2BX1 U8776 (.Y(n10911), 
	.B(n10910), 
	.AN(mem_write_en));
   NAND2X1 U8777 (.Y(n10910), 
	.B(n6343), 
	.A(n6591));
   OAI22X1 U8778 (.Y(n1029), 
	.B1(n10930), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6311));
   INVX1 U8779 (.Y(n10930), 
	.A(\ram[27][15] ));
   OAI22X1 U8780 (.Y(n1028), 
	.B1(n10931), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6314));
   INVX1 U8781 (.Y(n10931), 
	.A(\ram[27][14] ));
   OAI22X1 U8782 (.Y(n1027), 
	.B1(n10932), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6316));
   INVX1 U8783 (.Y(n10932), 
	.A(\ram[27][13] ));
   OAI22X1 U8784 (.Y(n1026), 
	.B1(n10933), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6318));
   INVX1 U8785 (.Y(n10933), 
	.A(\ram[27][12] ));
   OAI22X1 U8786 (.Y(n1025), 
	.B1(n10934), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6320));
   INVX1 U8787 (.Y(n10934), 
	.A(\ram[27][11] ));
   OAI22X1 U8788 (.Y(n1024), 
	.B1(n10935), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6322));
   INVX1 U8789 (.Y(n10935), 
	.A(\ram[27][10] ));
   OAI22X1 U8790 (.Y(n1023), 
	.B1(n10936), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6324));
   INVX1 U8791 (.Y(n10936), 
	.A(\ram[27][9] ));
   OAI22X1 U8792 (.Y(n1022), 
	.B1(n10937), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6326));
   INVX1 U8793 (.Y(n10937), 
	.A(\ram[27][8] ));
   OAI22X1 U8794 (.Y(n1021), 
	.B1(n10938), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6328));
   INVX1 U8795 (.Y(n10938), 
	.A(\ram[27][7] ));
   OAI22X1 U8796 (.Y(n1020), 
	.B1(n10939), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6330));
   INVX1 U8797 (.Y(n10939), 
	.A(\ram[27][6] ));
   OAI22X1 U8798 (.Y(n1019), 
	.B1(n10940), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6332));
   INVX1 U8799 (.Y(n10940), 
	.A(\ram[27][5] ));
   OAI22X1 U8800 (.Y(n1018), 
	.B1(n10941), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6334));
   INVX1 U8801 (.Y(n10941), 
	.A(\ram[27][4] ));
   OAI22X1 U8802 (.Y(n1017), 
	.B1(n10942), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6336));
   INVX1 U8803 (.Y(n10942), 
	.A(\ram[27][3] ));
   OAI22X1 U8804 (.Y(n1016), 
	.B1(n10943), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6338));
   INVX1 U8805 (.Y(n10943), 
	.A(\ram[27][2] ));
   OAI22X1 U8806 (.Y(n1015), 
	.B1(n10928), 
	.B0(n6306), 
	.A1(n10944), 
	.A0(n10929));
   NAND2X1 U8807 (.Y(n6306), 
	.B(mem_write_data[1]), 
	.A(mem_write_en));
   INVX1 U8808 (.Y(n10944), 
	.A(\ram[27][1] ));
   OAI22X1 U8809 (.Y(n1014), 
	.B1(n10945), 
	.B0(n10929), 
	.A1(n10928), 
	.A0(n6309));
   INVX1 U8810 (.Y(n10945), 
	.A(\ram[27][0] ));
   NOR2BX1 U8811 (.Y(n10929), 
	.B(n10928), 
	.AN(mem_write_en));
   NAND2X1 U8812 (.Y(n10928), 
	.B(n6343), 
	.A(n6610));
   NAND2X1 U8813 (.Y(n6309), 
	.B(mem_write_en), 
	.A(mem_write_data[0]));
   OAI22X1 U8814 (.Y(n1013), 
	.B1(n6311), 
	.B0(n6307), 
	.A1(n10946), 
	.A0(n6304));
   NAND2X1 U8815 (.Y(n6311), 
	.B(mem_write_en), 
	.A(mem_write_data[15]));
   INVX1 U8816 (.Y(n10946), 
	.A(\ram[26][15] ));
   OAI22X1 U8817 (.Y(n1012), 
	.B1(n6314), 
	.B0(n6307), 
	.A1(n10947), 
	.A0(n6304));
   NAND2X1 U8818 (.Y(n6314), 
	.B(mem_write_en), 
	.A(mem_write_data[14]));
   INVX1 U8819 (.Y(n10947), 
	.A(\ram[26][14] ));
   OAI22X1 U8820 (.Y(n1011), 
	.B1(n6316), 
	.B0(n6307), 
	.A1(n10948), 
	.A0(n6304));
   NAND2X1 U8821 (.Y(n6316), 
	.B(mem_write_en), 
	.A(mem_write_data[13]));
   INVX1 U8822 (.Y(n10948), 
	.A(\ram[26][13] ));
   OAI22X1 U8823 (.Y(n1010), 
	.B1(n6318), 
	.B0(n6307), 
	.A1(n10949), 
	.A0(n6304));
   NAND2X1 U8824 (.Y(n6318), 
	.B(mem_write_en), 
	.A(mem_write_data[12]));
   INVX1 U8825 (.Y(n10949), 
	.A(\ram[26][12] ));
   OAI22X1 U8826 (.Y(n1009), 
	.B1(n6320), 
	.B0(n6307), 
	.A1(n10950), 
	.A0(n6304));
   NAND2X1 U8827 (.Y(n6320), 
	.B(mem_write_en), 
	.A(mem_write_data[11]));
   INVX1 U8828 (.Y(n10950), 
	.A(\ram[26][11] ));
   OAI22X1 U8829 (.Y(n1008), 
	.B1(n6322), 
	.B0(n6307), 
	.A1(n10951), 
	.A0(n6304));
   NAND2X1 U8830 (.Y(n6322), 
	.B(mem_write_en), 
	.A(mem_write_data[10]));
   INVX1 U8831 (.Y(n10951), 
	.A(\ram[26][10] ));
   OAI22X1 U8832 (.Y(n1007), 
	.B1(n6324), 
	.B0(n6307), 
	.A1(n10952), 
	.A0(n6304));
   NAND2X1 U8833 (.Y(n6324), 
	.B(mem_write_en), 
	.A(mem_write_data[9]));
   INVX1 U8834 (.Y(n10952), 
	.A(\ram[26][9] ));
   OAI22X1 U8835 (.Y(n1006), 
	.B1(n6326), 
	.B0(n6307), 
	.A1(n10953), 
	.A0(n6304));
   NAND2X1 U8836 (.Y(n6326), 
	.B(mem_write_en), 
	.A(mem_write_data[8]));
   INVX1 U8837 (.Y(n10953), 
	.A(\ram[26][8] ));
   OAI22X1 U8838 (.Y(n1005), 
	.B1(n6328), 
	.B0(n6307), 
	.A1(n10954), 
	.A0(n6304));
   NAND2X1 U8839 (.Y(n6328), 
	.B(mem_write_en), 
	.A(mem_write_data[7]));
   INVX1 U8840 (.Y(n10954), 
	.A(\ram[26][7] ));
   OAI22X1 U8841 (.Y(n1004), 
	.B1(n6330), 
	.B0(n6307), 
	.A1(n10955), 
	.A0(n6304));
   NAND2X1 U8842 (.Y(n6330), 
	.B(mem_write_en), 
	.A(mem_write_data[6]));
   INVX1 U8843 (.Y(n10955), 
	.A(\ram[26][6] ));
   OAI22X1 U8844 (.Y(n1003), 
	.B1(n6332), 
	.B0(n6307), 
	.A1(n10956), 
	.A0(n6304));
   NAND2X1 U8845 (.Y(n6332), 
	.B(mem_write_en), 
	.A(mem_write_data[5]));
   INVX1 U8846 (.Y(n10956), 
	.A(\ram[26][5] ));
   OAI22X1 U8847 (.Y(n1002), 
	.B1(n6334), 
	.B0(n6307), 
	.A1(n10957), 
	.A0(n6304));
   NAND2X1 U8848 (.Y(n6334), 
	.B(mem_write_en), 
	.A(mem_write_data[4]));
   INVX1 U8849 (.Y(n10957), 
	.A(\ram[26][4] ));
   OAI22X1 U8850 (.Y(n1001), 
	.B1(n6336), 
	.B0(n6307), 
	.A1(n10958), 
	.A0(n6304));
   NAND2X1 U8851 (.Y(n6336), 
	.B(mem_write_en), 
	.A(mem_write_data[3]));
   INVX1 U8852 (.Y(n10958), 
	.A(\ram[26][3] ));
   OAI22X1 U8853 (.Y(n1000), 
	.B1(n10959), 
	.B0(n6304), 
	.A1(n6338), 
	.A0(n6307));
   INVX1 U8854 (.Y(n10959), 
	.A(\ram[26][2] ));
   NOR2BX1 U8855 (.Y(n6304), 
	.B(n6307), 
	.AN(mem_write_en));
   NAND2X1 U8856 (.Y(n6338), 
	.B(mem_write_en), 
	.A(mem_write_data[2]));
   NAND2X1 U8857 (.Y(n6307), 
	.B(n6343), 
	.A(n6629));
   OR4X1 U8858 (.Y(mem_read_data[9]), 
	.D(n10963), 
	.C(n10962), 
	.B(n10961), 
	.A(n10960));
   NAND4X1 U8859 (.Y(n10963), 
	.D(n10967), 
	.C(n10966), 
	.B(n10965), 
	.A(n10964));
   OAI21XL U8860 (.Y(n10967), 
	.B0(n6534), 
	.A1(n10969), 
	.A0(n10968));
   NAND4X1 U8861 (.Y(n10969), 
	.D(n10973), 
	.C(n10972), 
	.B(n10971), 
	.A(n10970));
   AOI22X1 U8862 (.Y(n10973), 
	.B1(n6342), 
	.B0(\ram[9][9] ), 
	.A1(n6362), 
	.A0(\ram[8][9] ));
   AOI22X1 U8863 (.Y(n10972), 
	.B1(n6381), 
	.B0(\ram[7][9] ), 
	.A1(n6400), 
	.A0(\ram[6][9] ));
   AOI22X1 U8864 (.Y(n10971), 
	.B1(n6419), 
	.B0(\ram[5][9] ), 
	.A1(n6438), 
	.A0(\ram[4][9] ));
   AOI22X1 U8865 (.Y(n10970), 
	.B1(n6457), 
	.B0(\ram[3][9] ), 
	.A1(n6476), 
	.A0(\ram[2][9] ));
   NAND4X1 U8866 (.Y(n10968), 
	.D(n10977), 
	.C(n10976), 
	.B(n10975), 
	.A(n10974));
   AOI22X1 U8867 (.Y(n10977), 
	.B1(n6495), 
	.B0(\ram[1][9] ), 
	.A1(n6514), 
	.A0(\ram[0][9] ));
   AOI22X1 U8868 (.Y(n10976), 
	.B1(n6533), 
	.B0(\ram[15][9] ), 
	.A1(n6553), 
	.A0(\ram[14][9] ));
   AOI22X1 U8869 (.Y(n10975), 
	.B1(n6572), 
	.B0(\ram[13][9] ), 
	.A1(n6591), 
	.A0(\ram[12][9] ));
   AOI22X1 U8870 (.Y(n10974), 
	.B1(n6610), 
	.B0(\ram[11][9] ), 
	.A1(n6629), 
	.A0(\ram[10][9] ));
   OAI21XL U8871 (.Y(n10966), 
	.B0(n6828), 
	.A1(n10979), 
	.A0(n10978));
   NAND4X1 U8872 (.Y(n10979), 
	.D(n10983), 
	.C(n10982), 
	.B(n10981), 
	.A(n10980));
   AOI22X1 U8873 (.Y(n10983), 
	.B1(n6342), 
	.B0(\ram[249][9] ), 
	.A1(n6362), 
	.A0(\ram[248][9] ));
   AOI22X1 U8874 (.Y(n10982), 
	.B1(n6381), 
	.B0(\ram[247][9] ), 
	.A1(n6400), 
	.A0(\ram[246][9] ));
   AOI22X1 U8875 (.Y(n10981), 
	.B1(n6419), 
	.B0(\ram[245][9] ), 
	.A1(n6438), 
	.A0(\ram[244][9] ));
   AOI22X1 U8876 (.Y(n10980), 
	.B1(n6457), 
	.B0(\ram[243][9] ), 
	.A1(n6476), 
	.A0(\ram[242][9] ));
   NAND4X1 U8877 (.Y(n10978), 
	.D(n10987), 
	.C(n10986), 
	.B(n10985), 
	.A(n10984));
   AOI22X1 U8878 (.Y(n10987), 
	.B1(n6495), 
	.B0(\ram[241][9] ), 
	.A1(n6514), 
	.A0(\ram[240][9] ));
   AOI22X1 U8879 (.Y(n10986), 
	.B1(n6533), 
	.B0(\ram[255][9] ), 
	.A1(n6553), 
	.A0(\ram[254][9] ));
   AOI22X1 U8880 (.Y(n10985), 
	.B1(n6572), 
	.B0(\ram[253][9] ), 
	.A1(n6591), 
	.A0(\ram[252][9] ));
   AOI22X1 U8881 (.Y(n10984), 
	.B1(n6610), 
	.B0(\ram[251][9] ), 
	.A1(n6629), 
	.A0(\ram[250][9] ));
   OAI21XL U8882 (.Y(n10965), 
	.B0(n7117), 
	.A1(n10989), 
	.A0(n10988));
   NAND4X1 U8883 (.Y(n10989), 
	.D(n10993), 
	.C(n10992), 
	.B(n10991), 
	.A(n10990));
   AOI22X1 U8884 (.Y(n10993), 
	.B1(n6342), 
	.B0(\ram[233][9] ), 
	.A1(n6362), 
	.A0(\ram[232][9] ));
   AOI22X1 U8885 (.Y(n10992), 
	.B1(n6381), 
	.B0(\ram[231][9] ), 
	.A1(n6400), 
	.A0(\ram[230][9] ));
   AOI22X1 U8886 (.Y(n10991), 
	.B1(n6419), 
	.B0(\ram[229][9] ), 
	.A1(n6438), 
	.A0(\ram[228][9] ));
   AOI22X1 U8887 (.Y(n10990), 
	.B1(n6457), 
	.B0(\ram[227][9] ), 
	.A1(n6476), 
	.A0(\ram[226][9] ));
   NAND4X1 U8888 (.Y(n10988), 
	.D(n10997), 
	.C(n10996), 
	.B(n10995), 
	.A(n10994));
   AOI22X1 U8889 (.Y(n10997), 
	.B1(n6495), 
	.B0(\ram[225][9] ), 
	.A1(n6514), 
	.A0(\ram[224][9] ));
   AOI22X1 U8890 (.Y(n10996), 
	.B1(n6533), 
	.B0(\ram[239][9] ), 
	.A1(n6553), 
	.A0(\ram[238][9] ));
   AOI22X1 U8891 (.Y(n10995), 
	.B1(n6572), 
	.B0(\ram[237][9] ), 
	.A1(n6591), 
	.A0(\ram[236][9] ));
   AOI22X1 U8892 (.Y(n10994), 
	.B1(n6610), 
	.B0(\ram[235][9] ), 
	.A1(n6629), 
	.A0(\ram[234][9] ));
   OAI21XL U8893 (.Y(n10964), 
	.B0(n7406), 
	.A1(n10999), 
	.A0(n10998));
   NAND4X1 U8894 (.Y(n10999), 
	.D(n11003), 
	.C(n11002), 
	.B(n11001), 
	.A(n11000));
   AOI22X1 U8895 (.Y(n11003), 
	.B1(n6342), 
	.B0(\ram[217][9] ), 
	.A1(n6362), 
	.A0(\ram[216][9] ));
   AOI22X1 U8896 (.Y(n11002), 
	.B1(n6381), 
	.B0(\ram[215][9] ), 
	.A1(n6400), 
	.A0(\ram[214][9] ));
   AOI22X1 U8897 (.Y(n11001), 
	.B1(n6419), 
	.B0(\ram[213][9] ), 
	.A1(n6438), 
	.A0(\ram[212][9] ));
   AOI22X1 U8898 (.Y(n11000), 
	.B1(n6457), 
	.B0(\ram[211][9] ), 
	.A1(n6476), 
	.A0(\ram[210][9] ));
   NAND4X1 U8899 (.Y(n10998), 
	.D(n11007), 
	.C(n11006), 
	.B(n11005), 
	.A(n11004));
   AOI22X1 U8900 (.Y(n11007), 
	.B1(n6495), 
	.B0(\ram[209][9] ), 
	.A1(n6514), 
	.A0(\ram[208][9] ));
   AOI22X1 U8901 (.Y(n11006), 
	.B1(n6533), 
	.B0(\ram[223][9] ), 
	.A1(n6553), 
	.A0(\ram[222][9] ));
   AOI22X1 U8902 (.Y(n11005), 
	.B1(n6572), 
	.B0(\ram[221][9] ), 
	.A1(n6591), 
	.A0(\ram[220][9] ));
   AOI22X1 U8903 (.Y(n11004), 
	.B1(n6610), 
	.B0(\ram[219][9] ), 
	.A1(n6629), 
	.A0(\ram[218][9] ));
   NAND4X1 U8904 (.Y(n10962), 
	.D(n11011), 
	.C(n11010), 
	.B(n11009), 
	.A(n11008));
   OAI21XL U8905 (.Y(n11011), 
	.B0(n7695), 
	.A1(n11013), 
	.A0(n11012));
   NAND4X1 U8906 (.Y(n11013), 
	.D(n11017), 
	.C(n11016), 
	.B(n11015), 
	.A(n11014));
   AOI22X1 U8907 (.Y(n11017), 
	.B1(n6342), 
	.B0(\ram[201][9] ), 
	.A1(n6362), 
	.A0(\ram[200][9] ));
   AOI22X1 U8908 (.Y(n11016), 
	.B1(n6381), 
	.B0(\ram[199][9] ), 
	.A1(n6400), 
	.A0(\ram[198][9] ));
   AOI22X1 U8909 (.Y(n11015), 
	.B1(n6419), 
	.B0(\ram[197][9] ), 
	.A1(n6438), 
	.A0(\ram[196][9] ));
   AOI22X1 U8910 (.Y(n11014), 
	.B1(n6457), 
	.B0(\ram[195][9] ), 
	.A1(n6476), 
	.A0(\ram[194][9] ));
   NAND4X1 U8911 (.Y(n11012), 
	.D(n11021), 
	.C(n11020), 
	.B(n11019), 
	.A(n11018));
   AOI22X1 U8912 (.Y(n11021), 
	.B1(n6495), 
	.B0(\ram[193][9] ), 
	.A1(n6514), 
	.A0(\ram[192][9] ));
   AOI22X1 U8913 (.Y(n11020), 
	.B1(n6533), 
	.B0(\ram[207][9] ), 
	.A1(n6553), 
	.A0(\ram[206][9] ));
   AOI22X1 U8914 (.Y(n11019), 
	.B1(n6572), 
	.B0(\ram[205][9] ), 
	.A1(n6591), 
	.A0(\ram[204][9] ));
   AOI22X1 U8915 (.Y(n11018), 
	.B1(n6610), 
	.B0(\ram[203][9] ), 
	.A1(n6629), 
	.A0(\ram[202][9] ));
   OAI21XL U8916 (.Y(n11010), 
	.B0(n7984), 
	.A1(n11023), 
	.A0(n11022));
   NAND4X1 U8917 (.Y(n11023), 
	.D(n11027), 
	.C(n11026), 
	.B(n11025), 
	.A(n11024));
   AOI22X1 U8918 (.Y(n11027), 
	.B1(n6342), 
	.B0(\ram[185][9] ), 
	.A1(n6362), 
	.A0(\ram[184][9] ));
   AOI22X1 U8919 (.Y(n11026), 
	.B1(n6381), 
	.B0(\ram[183][9] ), 
	.A1(n6400), 
	.A0(\ram[182][9] ));
   AOI22X1 U8920 (.Y(n11025), 
	.B1(n6419), 
	.B0(\ram[181][9] ), 
	.A1(n6438), 
	.A0(\ram[180][9] ));
   AOI22X1 U8921 (.Y(n11024), 
	.B1(n6457), 
	.B0(\ram[179][9] ), 
	.A1(n6476), 
	.A0(\ram[178][9] ));
   NAND4X1 U8922 (.Y(n11022), 
	.D(n11031), 
	.C(n11030), 
	.B(n11029), 
	.A(n11028));
   AOI22X1 U8923 (.Y(n11031), 
	.B1(n6495), 
	.B0(\ram[177][9] ), 
	.A1(n6514), 
	.A0(\ram[176][9] ));
   AOI22X1 U8924 (.Y(n11030), 
	.B1(n6533), 
	.B0(\ram[191][9] ), 
	.A1(n6553), 
	.A0(\ram[190][9] ));
   AOI22X1 U8925 (.Y(n11029), 
	.B1(n6572), 
	.B0(\ram[189][9] ), 
	.A1(n6591), 
	.A0(\ram[188][9] ));
   AOI22X1 U8926 (.Y(n11028), 
	.B1(n6610), 
	.B0(\ram[187][9] ), 
	.A1(n6629), 
	.A0(\ram[186][9] ));
   OAI21XL U8927 (.Y(n11009), 
	.B0(n8273), 
	.A1(n11033), 
	.A0(n11032));
   NAND4X1 U8928 (.Y(n11033), 
	.D(n11037), 
	.C(n11036), 
	.B(n11035), 
	.A(n11034));
   AOI22X1 U8929 (.Y(n11037), 
	.B1(n6342), 
	.B0(\ram[169][9] ), 
	.A1(n6362), 
	.A0(\ram[168][9] ));
   AOI22X1 U8930 (.Y(n11036), 
	.B1(n6381), 
	.B0(\ram[167][9] ), 
	.A1(n6400), 
	.A0(\ram[166][9] ));
   AOI22X1 U8931 (.Y(n11035), 
	.B1(n6419), 
	.B0(\ram[165][9] ), 
	.A1(n6438), 
	.A0(\ram[164][9] ));
   AOI22X1 U8932 (.Y(n11034), 
	.B1(n6457), 
	.B0(\ram[163][9] ), 
	.A1(n6476), 
	.A0(\ram[162][9] ));
   NAND4X1 U8933 (.Y(n11032), 
	.D(n11041), 
	.C(n11040), 
	.B(n11039), 
	.A(n11038));
   AOI22X1 U8934 (.Y(n11041), 
	.B1(n6495), 
	.B0(\ram[161][9] ), 
	.A1(n6514), 
	.A0(\ram[160][9] ));
   AOI22X1 U8935 (.Y(n11040), 
	.B1(n6533), 
	.B0(\ram[175][9] ), 
	.A1(n6553), 
	.A0(\ram[174][9] ));
   AOI22X1 U8936 (.Y(n11039), 
	.B1(n6572), 
	.B0(\ram[173][9] ), 
	.A1(n6591), 
	.A0(\ram[172][9] ));
   AOI22X1 U8937 (.Y(n11038), 
	.B1(n6610), 
	.B0(\ram[171][9] ), 
	.A1(n6629), 
	.A0(\ram[170][9] ));
   OAI21XL U8938 (.Y(n11008), 
	.B0(n8562), 
	.A1(n11043), 
	.A0(n11042));
   NAND4X1 U8939 (.Y(n11043), 
	.D(n11047), 
	.C(n11046), 
	.B(n11045), 
	.A(n11044));
   AOI22X1 U8940 (.Y(n11047), 
	.B1(n6342), 
	.B0(\ram[153][9] ), 
	.A1(n6362), 
	.A0(\ram[152][9] ));
   AOI22X1 U8941 (.Y(n11046), 
	.B1(n6381), 
	.B0(\ram[151][9] ), 
	.A1(n6400), 
	.A0(\ram[150][9] ));
   AOI22X1 U8942 (.Y(n11045), 
	.B1(n6419), 
	.B0(\ram[149][9] ), 
	.A1(n6438), 
	.A0(\ram[148][9] ));
   AOI22X1 U8943 (.Y(n11044), 
	.B1(n6457), 
	.B0(\ram[147][9] ), 
	.A1(n6476), 
	.A0(\ram[146][9] ));
   NAND4X1 U8944 (.Y(n11042), 
	.D(n11051), 
	.C(n11050), 
	.B(n11049), 
	.A(n11048));
   AOI22X1 U8945 (.Y(n11051), 
	.B1(n6495), 
	.B0(\ram[145][9] ), 
	.A1(n6514), 
	.A0(\ram[144][9] ));
   AOI22X1 U8946 (.Y(n11050), 
	.B1(n6533), 
	.B0(\ram[159][9] ), 
	.A1(n6553), 
	.A0(\ram[158][9] ));
   AOI22X1 U8947 (.Y(n11049), 
	.B1(n6572), 
	.B0(\ram[157][9] ), 
	.A1(n6591), 
	.A0(\ram[156][9] ));
   AOI22X1 U8948 (.Y(n11048), 
	.B1(n6610), 
	.B0(\ram[155][9] ), 
	.A1(n6629), 
	.A0(\ram[154][9] ));
   NAND4X1 U8949 (.Y(n10961), 
	.D(n11055), 
	.C(n11054), 
	.B(n11053), 
	.A(n11052));
   OAI21XL U8950 (.Y(n11055), 
	.B0(n8851), 
	.A1(n11057), 
	.A0(n11056));
   NAND4X1 U8951 (.Y(n11057), 
	.D(n11061), 
	.C(n11060), 
	.B(n11059), 
	.A(n11058));
   AOI22X1 U8952 (.Y(n11061), 
	.B1(n6342), 
	.B0(\ram[137][9] ), 
	.A1(n6362), 
	.A0(\ram[136][9] ));
   AOI22X1 U8953 (.Y(n11060), 
	.B1(n6381), 
	.B0(\ram[135][9] ), 
	.A1(n6400), 
	.A0(\ram[134][9] ));
   AOI22X1 U8954 (.Y(n11059), 
	.B1(n6419), 
	.B0(\ram[133][9] ), 
	.A1(n6438), 
	.A0(\ram[132][9] ));
   AOI22X1 U8955 (.Y(n11058), 
	.B1(n6457), 
	.B0(\ram[131][9] ), 
	.A1(n6476), 
	.A0(\ram[130][9] ));
   NAND4X1 U8956 (.Y(n11056), 
	.D(n11065), 
	.C(n11064), 
	.B(n11063), 
	.A(n11062));
   AOI22X1 U8957 (.Y(n11065), 
	.B1(n6495), 
	.B0(\ram[129][9] ), 
	.A1(n6514), 
	.A0(\ram[128][9] ));
   AOI22X1 U8958 (.Y(n11064), 
	.B1(n6533), 
	.B0(\ram[143][9] ), 
	.A1(n6553), 
	.A0(\ram[142][9] ));
   AOI22X1 U8959 (.Y(n11063), 
	.B1(n6572), 
	.B0(\ram[141][9] ), 
	.A1(n6591), 
	.A0(\ram[140][9] ));
   AOI22X1 U8960 (.Y(n11062), 
	.B1(n6610), 
	.B0(\ram[139][9] ), 
	.A1(n6629), 
	.A0(\ram[138][9] ));
   OAI21XL U8961 (.Y(n11054), 
	.B0(n9140), 
	.A1(n11067), 
	.A0(n11066));
   NAND4X1 U8962 (.Y(n11067), 
	.D(n11071), 
	.C(n11070), 
	.B(n11069), 
	.A(n11068));
   AOI22X1 U8963 (.Y(n11071), 
	.B1(n6342), 
	.B0(\ram[121][9] ), 
	.A1(n6362), 
	.A0(\ram[120][9] ));
   AOI22X1 U8964 (.Y(n11070), 
	.B1(n6381), 
	.B0(\ram[119][9] ), 
	.A1(n6400), 
	.A0(\ram[118][9] ));
   AOI22X1 U8965 (.Y(n11069), 
	.B1(n6419), 
	.B0(\ram[117][9] ), 
	.A1(n6438), 
	.A0(\ram[116][9] ));
   AOI22X1 U8966 (.Y(n11068), 
	.B1(n6457), 
	.B0(\ram[115][9] ), 
	.A1(n6476), 
	.A0(\ram[114][9] ));
   NAND4X1 U8967 (.Y(n11066), 
	.D(n11075), 
	.C(n11074), 
	.B(n11073), 
	.A(n11072));
   AOI22X1 U8968 (.Y(n11075), 
	.B1(n6495), 
	.B0(\ram[113][9] ), 
	.A1(n6514), 
	.A0(\ram[112][9] ));
   AOI22X1 U8969 (.Y(n11074), 
	.B1(n6533), 
	.B0(\ram[127][9] ), 
	.A1(n6553), 
	.A0(\ram[126][9] ));
   AOI22X1 U8970 (.Y(n11073), 
	.B1(n6572), 
	.B0(\ram[125][9] ), 
	.A1(n6591), 
	.A0(\ram[124][9] ));
   AOI22X1 U8971 (.Y(n11072), 
	.B1(n6610), 
	.B0(\ram[123][9] ), 
	.A1(n6629), 
	.A0(\ram[122][9] ));
   OAI21XL U8972 (.Y(n11053), 
	.B0(n9429), 
	.A1(n11077), 
	.A0(n11076));
   NAND4X1 U8973 (.Y(n11077), 
	.D(n11081), 
	.C(n11080), 
	.B(n11079), 
	.A(n11078));
   AOI22X1 U8974 (.Y(n11081), 
	.B1(n6342), 
	.B0(\ram[105][9] ), 
	.A1(n6362), 
	.A0(\ram[104][9] ));
   AOI22X1 U8975 (.Y(n11080), 
	.B1(n6381), 
	.B0(\ram[103][9] ), 
	.A1(n6400), 
	.A0(\ram[102][9] ));
   AOI22X1 U8976 (.Y(n11079), 
	.B1(n6419), 
	.B0(\ram[101][9] ), 
	.A1(n6438), 
	.A0(\ram[100][9] ));
   AOI22X1 U8977 (.Y(n11078), 
	.B1(n6457), 
	.B0(\ram[99][9] ), 
	.A1(n6476), 
	.A0(\ram[98][9] ));
   NAND4X1 U8978 (.Y(n11076), 
	.D(n11085), 
	.C(n11084), 
	.B(n11083), 
	.A(n11082));
   AOI22X1 U8979 (.Y(n11085), 
	.B1(n6495), 
	.B0(\ram[97][9] ), 
	.A1(n6514), 
	.A0(\ram[96][9] ));
   AOI22X1 U8980 (.Y(n11084), 
	.B1(n6533), 
	.B0(\ram[111][9] ), 
	.A1(n6553), 
	.A0(\ram[110][9] ));
   AOI22X1 U8981 (.Y(n11083), 
	.B1(n6572), 
	.B0(\ram[109][9] ), 
	.A1(n6591), 
	.A0(\ram[108][9] ));
   AOI22X1 U8982 (.Y(n11082), 
	.B1(n6610), 
	.B0(\ram[107][9] ), 
	.A1(n6629), 
	.A0(\ram[106][9] ));
   OAI21XL U8983 (.Y(n11052), 
	.B0(n9718), 
	.A1(n11087), 
	.A0(n11086));
   NAND4X1 U8984 (.Y(n11087), 
	.D(n11091), 
	.C(n11090), 
	.B(n11089), 
	.A(n11088));
   AOI22X1 U8985 (.Y(n11091), 
	.B1(n6342), 
	.B0(\ram[89][9] ), 
	.A1(n6362), 
	.A0(\ram[88][9] ));
   AOI22X1 U8986 (.Y(n11090), 
	.B1(n6381), 
	.B0(\ram[87][9] ), 
	.A1(n6400), 
	.A0(\ram[86][9] ));
   AOI22X1 U8987 (.Y(n11089), 
	.B1(n6419), 
	.B0(\ram[85][9] ), 
	.A1(n6438), 
	.A0(\ram[84][9] ));
   AOI22X1 U8988 (.Y(n11088), 
	.B1(n6457), 
	.B0(\ram[83][9] ), 
	.A1(n6476), 
	.A0(\ram[82][9] ));
   NAND4X1 U8989 (.Y(n11086), 
	.D(n11095), 
	.C(n11094), 
	.B(n11093), 
	.A(n11092));
   AOI22X1 U8990 (.Y(n11095), 
	.B1(n6495), 
	.B0(\ram[81][9] ), 
	.A1(n6514), 
	.A0(\ram[80][9] ));
   AOI22X1 U8991 (.Y(n11094), 
	.B1(n6533), 
	.B0(\ram[95][9] ), 
	.A1(n6553), 
	.A0(\ram[94][9] ));
   AOI22X1 U8992 (.Y(n11093), 
	.B1(n6572), 
	.B0(\ram[93][9] ), 
	.A1(n6591), 
	.A0(\ram[92][9] ));
   AOI22X1 U8993 (.Y(n11092), 
	.B1(n6610), 
	.B0(\ram[91][9] ), 
	.A1(n6629), 
	.A0(\ram[90][9] ));
   NAND4X1 U8994 (.Y(n10960), 
	.D(n11099), 
	.C(n11098), 
	.B(n11097), 
	.A(n11096));
   OAI21XL U8995 (.Y(n11099), 
	.B0(n10007), 
	.A1(n11101), 
	.A0(n11100));
   NAND4X1 U8996 (.Y(n11101), 
	.D(n11105), 
	.C(n11104), 
	.B(n11103), 
	.A(n11102));
   AOI22X1 U8997 (.Y(n11105), 
	.B1(n6342), 
	.B0(\ram[73][9] ), 
	.A1(n6362), 
	.A0(\ram[72][9] ));
   AOI22X1 U8998 (.Y(n11104), 
	.B1(n6381), 
	.B0(\ram[71][9] ), 
	.A1(n6400), 
	.A0(\ram[70][9] ));
   AOI22X1 U8999 (.Y(n11103), 
	.B1(n6419), 
	.B0(\ram[69][9] ), 
	.A1(n6438), 
	.A0(\ram[68][9] ));
   AOI22X1 U9000 (.Y(n11102), 
	.B1(n6457), 
	.B0(\ram[67][9] ), 
	.A1(n6476), 
	.A0(\ram[66][9] ));
   NAND4X1 U9001 (.Y(n11100), 
	.D(n11109), 
	.C(n11108), 
	.B(n11107), 
	.A(n11106));
   AOI22X1 U9002 (.Y(n11109), 
	.B1(n6495), 
	.B0(\ram[65][9] ), 
	.A1(n6514), 
	.A0(\ram[64][9] ));
   AOI22X1 U9003 (.Y(n11108), 
	.B1(n6533), 
	.B0(\ram[79][9] ), 
	.A1(n6553), 
	.A0(\ram[78][9] ));
   AOI22X1 U9004 (.Y(n11107), 
	.B1(n6572), 
	.B0(\ram[77][9] ), 
	.A1(n6591), 
	.A0(\ram[76][9] ));
   AOI22X1 U9005 (.Y(n11106), 
	.B1(n6610), 
	.B0(\ram[75][9] ), 
	.A1(n6629), 
	.A0(\ram[74][9] ));
   OAI21XL U9006 (.Y(n11098), 
	.B0(n10296), 
	.A1(n11111), 
	.A0(n11110));
   NAND4X1 U9007 (.Y(n11111), 
	.D(n11115), 
	.C(n11114), 
	.B(n11113), 
	.A(n11112));
   AOI22X1 U9008 (.Y(n11115), 
	.B1(n6342), 
	.B0(\ram[57][9] ), 
	.A1(n6362), 
	.A0(\ram[56][9] ));
   AOI22X1 U9009 (.Y(n11114), 
	.B1(n6381), 
	.B0(\ram[55][9] ), 
	.A1(n6400), 
	.A0(\ram[54][9] ));
   AOI22X1 U9010 (.Y(n11113), 
	.B1(n6419), 
	.B0(\ram[53][9] ), 
	.A1(n6438), 
	.A0(\ram[52][9] ));
   AOI22X1 U9011 (.Y(n11112), 
	.B1(n6457), 
	.B0(\ram[51][9] ), 
	.A1(n6476), 
	.A0(\ram[50][9] ));
   NAND4X1 U9012 (.Y(n11110), 
	.D(n11119), 
	.C(n11118), 
	.B(n11117), 
	.A(n11116));
   AOI22X1 U9013 (.Y(n11119), 
	.B1(n6495), 
	.B0(\ram[49][9] ), 
	.A1(n6514), 
	.A0(\ram[48][9] ));
   AOI22X1 U9014 (.Y(n11118), 
	.B1(n6533), 
	.B0(\ram[63][9] ), 
	.A1(n6553), 
	.A0(\ram[62][9] ));
   AOI22X1 U9015 (.Y(n11117), 
	.B1(n6572), 
	.B0(\ram[61][9] ), 
	.A1(n6591), 
	.A0(\ram[60][9] ));
   AOI22X1 U9016 (.Y(n11116), 
	.B1(n6610), 
	.B0(\ram[59][9] ), 
	.A1(n6629), 
	.A0(\ram[58][9] ));
   OAI21XL U9017 (.Y(n11097), 
	.B0(n10585), 
	.A1(n11121), 
	.A0(n11120));
   NAND4X1 U9018 (.Y(n11121), 
	.D(n11125), 
	.C(n11124), 
	.B(n11123), 
	.A(n11122));
   AOI22X1 U9019 (.Y(n11125), 
	.B1(n6342), 
	.B0(\ram[41][9] ), 
	.A1(n6362), 
	.A0(\ram[40][9] ));
   AOI22X1 U9020 (.Y(n11124), 
	.B1(n6381), 
	.B0(\ram[39][9] ), 
	.A1(n6400), 
	.A0(\ram[38][9] ));
   AOI22X1 U9021 (.Y(n11123), 
	.B1(n6419), 
	.B0(\ram[37][9] ), 
	.A1(n6438), 
	.A0(\ram[36][9] ));
   AOI22X1 U9022 (.Y(n11122), 
	.B1(n6457), 
	.B0(\ram[35][9] ), 
	.A1(n6476), 
	.A0(\ram[34][9] ));
   NAND4X1 U9023 (.Y(n11120), 
	.D(n11129), 
	.C(n11128), 
	.B(n11127), 
	.A(n11126));
   AOI22X1 U9024 (.Y(n11129), 
	.B1(n6495), 
	.B0(\ram[33][9] ), 
	.A1(n6514), 
	.A0(\ram[32][9] ));
   AOI22X1 U9025 (.Y(n11128), 
	.B1(n6533), 
	.B0(\ram[47][9] ), 
	.A1(n6553), 
	.A0(\ram[46][9] ));
   AOI22X1 U9026 (.Y(n11127), 
	.B1(n6572), 
	.B0(\ram[45][9] ), 
	.A1(n6591), 
	.A0(\ram[44][9] ));
   AOI22X1 U9027 (.Y(n11126), 
	.B1(n6610), 
	.B0(\ram[43][9] ), 
	.A1(n6629), 
	.A0(\ram[42][9] ));
   OAI21XL U9028 (.Y(n11096), 
	.B0(n6343), 
	.A1(n11131), 
	.A0(n11130));
   NAND4X1 U9029 (.Y(n11131), 
	.D(n11135), 
	.C(n11134), 
	.B(n11133), 
	.A(n11132));
   AOI22X1 U9030 (.Y(n11135), 
	.B1(n6342), 
	.B0(\ram[25][9] ), 
	.A1(n6362), 
	.A0(\ram[24][9] ));
   AOI22X1 U9031 (.Y(n11134), 
	.B1(n6381), 
	.B0(\ram[23][9] ), 
	.A1(n6400), 
	.A0(\ram[22][9] ));
   AOI22X1 U9032 (.Y(n11133), 
	.B1(n6419), 
	.B0(\ram[21][9] ), 
	.A1(n6438), 
	.A0(\ram[20][9] ));
   AOI22X1 U9033 (.Y(n11132), 
	.B1(n6457), 
	.B0(\ram[19][9] ), 
	.A1(n6476), 
	.A0(\ram[18][9] ));
   NAND4X1 U9034 (.Y(n11130), 
	.D(n11139), 
	.C(n11138), 
	.B(n11137), 
	.A(n11136));
   AOI22X1 U9035 (.Y(n11139), 
	.B1(n6495), 
	.B0(\ram[17][9] ), 
	.A1(n6514), 
	.A0(\ram[16][9] ));
   AOI22X1 U9036 (.Y(n11138), 
	.B1(n6533), 
	.B0(\ram[31][9] ), 
	.A1(n6553), 
	.A0(\ram[30][9] ));
   AOI22X1 U9037 (.Y(n11137), 
	.B1(n6572), 
	.B0(\ram[29][9] ), 
	.A1(n6591), 
	.A0(\ram[28][9] ));
   AOI22X1 U9038 (.Y(n11136), 
	.B1(n6610), 
	.B0(\ram[27][9] ), 
	.A1(n6629), 
	.A0(\ram[26][9] ));
   OR4X1 U9039 (.Y(mem_read_data[8]), 
	.D(n11143), 
	.C(n11142), 
	.B(n11141), 
	.A(n11140));
   NAND4X1 U9040 (.Y(n11143), 
	.D(n11147), 
	.C(n11146), 
	.B(n11145), 
	.A(n11144));
   OAI21XL U9041 (.Y(n11147), 
	.B0(n6534), 
	.A1(n11149), 
	.A0(n11148));
   NAND4X1 U9042 (.Y(n11149), 
	.D(n11153), 
	.C(n11152), 
	.B(n11151), 
	.A(n11150));
   AOI22X1 U9043 (.Y(n11153), 
	.B1(n6342), 
	.B0(\ram[9][8] ), 
	.A1(n6362), 
	.A0(\ram[8][8] ));
   AOI22X1 U9044 (.Y(n11152), 
	.B1(n6381), 
	.B0(\ram[7][8] ), 
	.A1(n6400), 
	.A0(\ram[6][8] ));
   AOI22X1 U9045 (.Y(n11151), 
	.B1(n6419), 
	.B0(\ram[5][8] ), 
	.A1(n6438), 
	.A0(\ram[4][8] ));
   AOI22X1 U9046 (.Y(n11150), 
	.B1(n6457), 
	.B0(\ram[3][8] ), 
	.A1(n6476), 
	.A0(\ram[2][8] ));
   NAND4X1 U9047 (.Y(n11148), 
	.D(n11157), 
	.C(n11156), 
	.B(n11155), 
	.A(n11154));
   AOI22X1 U9048 (.Y(n11157), 
	.B1(n6495), 
	.B0(\ram[1][8] ), 
	.A1(n6514), 
	.A0(\ram[0][8] ));
   AOI22X1 U9049 (.Y(n11156), 
	.B1(n6533), 
	.B0(\ram[15][8] ), 
	.A1(n6553), 
	.A0(\ram[14][8] ));
   AOI22X1 U9050 (.Y(n11155), 
	.B1(n6572), 
	.B0(\ram[13][8] ), 
	.A1(n6591), 
	.A0(\ram[12][8] ));
   AOI22X1 U9051 (.Y(n11154), 
	.B1(n6610), 
	.B0(\ram[11][8] ), 
	.A1(n6629), 
	.A0(\ram[10][8] ));
   OAI21XL U9052 (.Y(n11146), 
	.B0(n6828), 
	.A1(n11159), 
	.A0(n11158));
   NAND4X1 U9053 (.Y(n11159), 
	.D(n11163), 
	.C(n11162), 
	.B(n11161), 
	.A(n11160));
   AOI22X1 U9054 (.Y(n11163), 
	.B1(n6342), 
	.B0(\ram[249][8] ), 
	.A1(n6362), 
	.A0(\ram[248][8] ));
   AOI22X1 U9055 (.Y(n11162), 
	.B1(n6381), 
	.B0(\ram[247][8] ), 
	.A1(n6400), 
	.A0(\ram[246][8] ));
   AOI22X1 U9056 (.Y(n11161), 
	.B1(n6419), 
	.B0(\ram[245][8] ), 
	.A1(n6438), 
	.A0(\ram[244][8] ));
   AOI22X1 U9057 (.Y(n11160), 
	.B1(n6457), 
	.B0(\ram[243][8] ), 
	.A1(n6476), 
	.A0(\ram[242][8] ));
   NAND4X1 U9058 (.Y(n11158), 
	.D(n11167), 
	.C(n11166), 
	.B(n11165), 
	.A(n11164));
   AOI22X1 U9059 (.Y(n11167), 
	.B1(n6495), 
	.B0(\ram[241][8] ), 
	.A1(n6514), 
	.A0(\ram[240][8] ));
   AOI22X1 U9060 (.Y(n11166), 
	.B1(n6533), 
	.B0(\ram[255][8] ), 
	.A1(n6553), 
	.A0(\ram[254][8] ));
   AOI22X1 U9061 (.Y(n11165), 
	.B1(n6572), 
	.B0(\ram[253][8] ), 
	.A1(n6591), 
	.A0(\ram[252][8] ));
   AOI22X1 U9062 (.Y(n11164), 
	.B1(n6610), 
	.B0(\ram[251][8] ), 
	.A1(n6629), 
	.A0(\ram[250][8] ));
   OAI21XL U9063 (.Y(n11145), 
	.B0(n7117), 
	.A1(n11169), 
	.A0(n11168));
   NAND4X1 U9064 (.Y(n11169), 
	.D(n11173), 
	.C(n11172), 
	.B(n11171), 
	.A(n11170));
   AOI22X1 U9065 (.Y(n11173), 
	.B1(n6342), 
	.B0(\ram[233][8] ), 
	.A1(n6362), 
	.A0(\ram[232][8] ));
   AOI22X1 U9066 (.Y(n11172), 
	.B1(n6381), 
	.B0(\ram[231][8] ), 
	.A1(n6400), 
	.A0(\ram[230][8] ));
   AOI22X1 U9067 (.Y(n11171), 
	.B1(n6419), 
	.B0(\ram[229][8] ), 
	.A1(n6438), 
	.A0(\ram[228][8] ));
   AOI22X1 U9068 (.Y(n11170), 
	.B1(n6457), 
	.B0(\ram[227][8] ), 
	.A1(n6476), 
	.A0(\ram[226][8] ));
   NAND4X1 U9069 (.Y(n11168), 
	.D(n11177), 
	.C(n11176), 
	.B(n11175), 
	.A(n11174));
   AOI22X1 U9070 (.Y(n11177), 
	.B1(n6495), 
	.B0(\ram[225][8] ), 
	.A1(n6514), 
	.A0(\ram[224][8] ));
   AOI22X1 U9071 (.Y(n11176), 
	.B1(n6533), 
	.B0(\ram[239][8] ), 
	.A1(n6553), 
	.A0(\ram[238][8] ));
   AOI22X1 U9072 (.Y(n11175), 
	.B1(n6572), 
	.B0(\ram[237][8] ), 
	.A1(n6591), 
	.A0(\ram[236][8] ));
   AOI22X1 U9073 (.Y(n11174), 
	.B1(n6610), 
	.B0(\ram[235][8] ), 
	.A1(n6629), 
	.A0(\ram[234][8] ));
   OAI21XL U9074 (.Y(n11144), 
	.B0(n7406), 
	.A1(n11179), 
	.A0(n11178));
   NAND4X1 U9075 (.Y(n11179), 
	.D(n11183), 
	.C(n11182), 
	.B(n11181), 
	.A(n11180));
   AOI22X1 U9076 (.Y(n11183), 
	.B1(n6342), 
	.B0(\ram[217][8] ), 
	.A1(n6362), 
	.A0(\ram[216][8] ));
   AOI22X1 U9077 (.Y(n11182), 
	.B1(n6381), 
	.B0(\ram[215][8] ), 
	.A1(n6400), 
	.A0(\ram[214][8] ));
   AOI22X1 U9078 (.Y(n11181), 
	.B1(n6419), 
	.B0(\ram[213][8] ), 
	.A1(n6438), 
	.A0(\ram[212][8] ));
   AOI22X1 U9079 (.Y(n11180), 
	.B1(n6457), 
	.B0(\ram[211][8] ), 
	.A1(n6476), 
	.A0(\ram[210][8] ));
   NAND4X1 U9080 (.Y(n11178), 
	.D(n11187), 
	.C(n11186), 
	.B(n11185), 
	.A(n11184));
   AOI22X1 U9081 (.Y(n11187), 
	.B1(n6495), 
	.B0(\ram[209][8] ), 
	.A1(n6514), 
	.A0(\ram[208][8] ));
   AOI22X1 U9082 (.Y(n11186), 
	.B1(n6533), 
	.B0(\ram[223][8] ), 
	.A1(n6553), 
	.A0(\ram[222][8] ));
   AOI22X1 U9083 (.Y(n11185), 
	.B1(n6572), 
	.B0(\ram[221][8] ), 
	.A1(n6591), 
	.A0(\ram[220][8] ));
   AOI22X1 U9084 (.Y(n11184), 
	.B1(n6610), 
	.B0(\ram[219][8] ), 
	.A1(n6629), 
	.A0(\ram[218][8] ));
   NAND4X1 U9085 (.Y(n11142), 
	.D(n11191), 
	.C(n11190), 
	.B(n11189), 
	.A(n11188));
   OAI21XL U9086 (.Y(n11191), 
	.B0(n7695), 
	.A1(n11193), 
	.A0(n11192));
   NAND4X1 U9087 (.Y(n11193), 
	.D(n11197), 
	.C(n11196), 
	.B(n11195), 
	.A(n11194));
   AOI22X1 U9088 (.Y(n11197), 
	.B1(n6342), 
	.B0(\ram[201][8] ), 
	.A1(n6362), 
	.A0(\ram[200][8] ));
   AOI22X1 U9089 (.Y(n11196), 
	.B1(n6381), 
	.B0(\ram[199][8] ), 
	.A1(n6400), 
	.A0(\ram[198][8] ));
   AOI22X1 U9090 (.Y(n11195), 
	.B1(n6419), 
	.B0(\ram[197][8] ), 
	.A1(n6438), 
	.A0(\ram[196][8] ));
   AOI22X1 U9091 (.Y(n11194), 
	.B1(n6457), 
	.B0(\ram[195][8] ), 
	.A1(n6476), 
	.A0(\ram[194][8] ));
   NAND4X1 U9092 (.Y(n11192), 
	.D(n11201), 
	.C(n11200), 
	.B(n11199), 
	.A(n11198));
   AOI22X1 U9093 (.Y(n11201), 
	.B1(n6495), 
	.B0(\ram[193][8] ), 
	.A1(n6514), 
	.A0(\ram[192][8] ));
   AOI22X1 U9094 (.Y(n11200), 
	.B1(n6533), 
	.B0(\ram[207][8] ), 
	.A1(n6553), 
	.A0(\ram[206][8] ));
   AOI22X1 U9095 (.Y(n11199), 
	.B1(n6572), 
	.B0(\ram[205][8] ), 
	.A1(n6591), 
	.A0(\ram[204][8] ));
   AOI22X1 U9096 (.Y(n11198), 
	.B1(n6610), 
	.B0(\ram[203][8] ), 
	.A1(n6629), 
	.A0(\ram[202][8] ));
   OAI21XL U9097 (.Y(n11190), 
	.B0(n7984), 
	.A1(n11203), 
	.A0(n11202));
   NAND4X1 U9098 (.Y(n11203), 
	.D(n11207), 
	.C(n11206), 
	.B(n11205), 
	.A(n11204));
   AOI22X1 U9099 (.Y(n11207), 
	.B1(n6342), 
	.B0(\ram[185][8] ), 
	.A1(n6362), 
	.A0(\ram[184][8] ));
   AOI22X1 U9100 (.Y(n11206), 
	.B1(n6381), 
	.B0(\ram[183][8] ), 
	.A1(n6400), 
	.A0(\ram[182][8] ));
   AOI22X1 U9101 (.Y(n11205), 
	.B1(n6419), 
	.B0(\ram[181][8] ), 
	.A1(n6438), 
	.A0(\ram[180][8] ));
   AOI22X1 U9102 (.Y(n11204), 
	.B1(n6457), 
	.B0(\ram[179][8] ), 
	.A1(n6476), 
	.A0(\ram[178][8] ));
   NAND4X1 U9103 (.Y(n11202), 
	.D(n11211), 
	.C(n11210), 
	.B(n11209), 
	.A(n11208));
   AOI22X1 U9104 (.Y(n11211), 
	.B1(n6495), 
	.B0(\ram[177][8] ), 
	.A1(n6514), 
	.A0(\ram[176][8] ));
   AOI22X1 U9105 (.Y(n11210), 
	.B1(n6533), 
	.B0(\ram[191][8] ), 
	.A1(n6553), 
	.A0(\ram[190][8] ));
   AOI22X1 U9106 (.Y(n11209), 
	.B1(n6572), 
	.B0(\ram[189][8] ), 
	.A1(n6591), 
	.A0(\ram[188][8] ));
   AOI22X1 U9107 (.Y(n11208), 
	.B1(n6610), 
	.B0(\ram[187][8] ), 
	.A1(n6629), 
	.A0(\ram[186][8] ));
   OAI21XL U9108 (.Y(n11189), 
	.B0(n8273), 
	.A1(n11213), 
	.A0(n11212));
   NAND4X1 U9109 (.Y(n11213), 
	.D(n11217), 
	.C(n11216), 
	.B(n11215), 
	.A(n11214));
   AOI22X1 U9110 (.Y(n11217), 
	.B1(n6342), 
	.B0(\ram[169][8] ), 
	.A1(n6362), 
	.A0(\ram[168][8] ));
   AOI22X1 U9111 (.Y(n11216), 
	.B1(n6381), 
	.B0(\ram[167][8] ), 
	.A1(n6400), 
	.A0(\ram[166][8] ));
   AOI22X1 U9112 (.Y(n11215), 
	.B1(n6419), 
	.B0(\ram[165][8] ), 
	.A1(n6438), 
	.A0(\ram[164][8] ));
   AOI22X1 U9113 (.Y(n11214), 
	.B1(n6457), 
	.B0(\ram[163][8] ), 
	.A1(n6476), 
	.A0(\ram[162][8] ));
   NAND4X1 U9114 (.Y(n11212), 
	.D(n11221), 
	.C(n11220), 
	.B(n11219), 
	.A(n11218));
   AOI22X1 U9115 (.Y(n11221), 
	.B1(n6495), 
	.B0(\ram[161][8] ), 
	.A1(n6514), 
	.A0(\ram[160][8] ));
   AOI22X1 U9116 (.Y(n11220), 
	.B1(n6533), 
	.B0(\ram[175][8] ), 
	.A1(n6553), 
	.A0(\ram[174][8] ));
   AOI22X1 U9117 (.Y(n11219), 
	.B1(n6572), 
	.B0(\ram[173][8] ), 
	.A1(n6591), 
	.A0(\ram[172][8] ));
   AOI22X1 U9118 (.Y(n11218), 
	.B1(n6610), 
	.B0(\ram[171][8] ), 
	.A1(n6629), 
	.A0(\ram[170][8] ));
   OAI21XL U9119 (.Y(n11188), 
	.B0(n8562), 
	.A1(n11223), 
	.A0(n11222));
   NAND4X1 U9120 (.Y(n11223), 
	.D(n11227), 
	.C(n11226), 
	.B(n11225), 
	.A(n11224));
   AOI22X1 U9121 (.Y(n11227), 
	.B1(n6342), 
	.B0(\ram[153][8] ), 
	.A1(n6362), 
	.A0(\ram[152][8] ));
   AOI22X1 U9122 (.Y(n11226), 
	.B1(n6381), 
	.B0(\ram[151][8] ), 
	.A1(n6400), 
	.A0(\ram[150][8] ));
   AOI22X1 U9123 (.Y(n11225), 
	.B1(n6419), 
	.B0(\ram[149][8] ), 
	.A1(n6438), 
	.A0(\ram[148][8] ));
   AOI22X1 U9124 (.Y(n11224), 
	.B1(n6457), 
	.B0(\ram[147][8] ), 
	.A1(n6476), 
	.A0(\ram[146][8] ));
   NAND4X1 U9125 (.Y(n11222), 
	.D(n11231), 
	.C(n11230), 
	.B(n11229), 
	.A(n11228));
   AOI22X1 U9126 (.Y(n11231), 
	.B1(n6495), 
	.B0(\ram[145][8] ), 
	.A1(n6514), 
	.A0(\ram[144][8] ));
   AOI22X1 U9127 (.Y(n11230), 
	.B1(n6533), 
	.B0(\ram[159][8] ), 
	.A1(n6553), 
	.A0(\ram[158][8] ));
   AOI22X1 U9128 (.Y(n11229), 
	.B1(n6572), 
	.B0(\ram[157][8] ), 
	.A1(n6591), 
	.A0(\ram[156][8] ));
   AOI22X1 U9129 (.Y(n11228), 
	.B1(n6610), 
	.B0(\ram[155][8] ), 
	.A1(n6629), 
	.A0(\ram[154][8] ));
   NAND4X1 U9130 (.Y(n11141), 
	.D(n11235), 
	.C(n11234), 
	.B(n11233), 
	.A(n11232));
   OAI21XL U9131 (.Y(n11235), 
	.B0(n8851), 
	.A1(n11237), 
	.A0(n11236));
   NAND4X1 U9132 (.Y(n11237), 
	.D(n11241), 
	.C(n11240), 
	.B(n11239), 
	.A(n11238));
   AOI22X1 U9133 (.Y(n11241), 
	.B1(n6342), 
	.B0(\ram[137][8] ), 
	.A1(n6362), 
	.A0(\ram[136][8] ));
   AOI22X1 U9134 (.Y(n11240), 
	.B1(n6381), 
	.B0(\ram[135][8] ), 
	.A1(n6400), 
	.A0(\ram[134][8] ));
   AOI22X1 U9135 (.Y(n11239), 
	.B1(n6419), 
	.B0(\ram[133][8] ), 
	.A1(n6438), 
	.A0(\ram[132][8] ));
   AOI22X1 U9136 (.Y(n11238), 
	.B1(n6457), 
	.B0(\ram[131][8] ), 
	.A1(n6476), 
	.A0(\ram[130][8] ));
   NAND4X1 U9137 (.Y(n11236), 
	.D(n11245), 
	.C(n11244), 
	.B(n11243), 
	.A(n11242));
   AOI22X1 U9138 (.Y(n11245), 
	.B1(n6495), 
	.B0(\ram[129][8] ), 
	.A1(n6514), 
	.A0(\ram[128][8] ));
   AOI22X1 U9139 (.Y(n11244), 
	.B1(n6533), 
	.B0(\ram[143][8] ), 
	.A1(n6553), 
	.A0(\ram[142][8] ));
   AOI22X1 U9140 (.Y(n11243), 
	.B1(n6572), 
	.B0(\ram[141][8] ), 
	.A1(n6591), 
	.A0(\ram[140][8] ));
   AOI22X1 U9141 (.Y(n11242), 
	.B1(n6610), 
	.B0(\ram[139][8] ), 
	.A1(n6629), 
	.A0(\ram[138][8] ));
   OAI21XL U9142 (.Y(n11234), 
	.B0(n9140), 
	.A1(n11247), 
	.A0(n11246));
   NAND4X1 U9143 (.Y(n11247), 
	.D(n11251), 
	.C(n11250), 
	.B(n11249), 
	.A(n11248));
   AOI22X1 U9144 (.Y(n11251), 
	.B1(n6342), 
	.B0(\ram[121][8] ), 
	.A1(n6362), 
	.A0(\ram[120][8] ));
   AOI22X1 U9145 (.Y(n11250), 
	.B1(n6381), 
	.B0(\ram[119][8] ), 
	.A1(n6400), 
	.A0(\ram[118][8] ));
   AOI22X1 U9146 (.Y(n11249), 
	.B1(n6419), 
	.B0(\ram[117][8] ), 
	.A1(n6438), 
	.A0(\ram[116][8] ));
   AOI22X1 U9147 (.Y(n11248), 
	.B1(n6457), 
	.B0(\ram[115][8] ), 
	.A1(n6476), 
	.A0(\ram[114][8] ));
   NAND4X1 U9148 (.Y(n11246), 
	.D(n11255), 
	.C(n11254), 
	.B(n11253), 
	.A(n11252));
   AOI22X1 U9149 (.Y(n11255), 
	.B1(n6495), 
	.B0(\ram[113][8] ), 
	.A1(n6514), 
	.A0(\ram[112][8] ));
   AOI22X1 U9150 (.Y(n11254), 
	.B1(n6533), 
	.B0(\ram[127][8] ), 
	.A1(n6553), 
	.A0(\ram[126][8] ));
   AOI22X1 U9151 (.Y(n11253), 
	.B1(n6572), 
	.B0(\ram[125][8] ), 
	.A1(n6591), 
	.A0(\ram[124][8] ));
   AOI22X1 U9152 (.Y(n11252), 
	.B1(n6610), 
	.B0(\ram[123][8] ), 
	.A1(n6629), 
	.A0(\ram[122][8] ));
   OAI21XL U9153 (.Y(n11233), 
	.B0(n9429), 
	.A1(n11257), 
	.A0(n11256));
   NAND4X1 U9154 (.Y(n11257), 
	.D(n11261), 
	.C(n11260), 
	.B(n11259), 
	.A(n11258));
   AOI22X1 U9155 (.Y(n11261), 
	.B1(n6342), 
	.B0(\ram[105][8] ), 
	.A1(n6362), 
	.A0(\ram[104][8] ));
   AOI22X1 U9156 (.Y(n11260), 
	.B1(n6381), 
	.B0(\ram[103][8] ), 
	.A1(n6400), 
	.A0(\ram[102][8] ));
   AOI22X1 U9157 (.Y(n11259), 
	.B1(n6419), 
	.B0(\ram[101][8] ), 
	.A1(n6438), 
	.A0(\ram[100][8] ));
   AOI22X1 U9158 (.Y(n11258), 
	.B1(n6457), 
	.B0(\ram[99][8] ), 
	.A1(n6476), 
	.A0(\ram[98][8] ));
   NAND4X1 U9159 (.Y(n11256), 
	.D(n11265), 
	.C(n11264), 
	.B(n11263), 
	.A(n11262));
   AOI22X1 U9160 (.Y(n11265), 
	.B1(n6495), 
	.B0(\ram[97][8] ), 
	.A1(n6514), 
	.A0(\ram[96][8] ));
   AOI22X1 U9161 (.Y(n11264), 
	.B1(n6533), 
	.B0(\ram[111][8] ), 
	.A1(n6553), 
	.A0(\ram[110][8] ));
   AOI22X1 U9162 (.Y(n11263), 
	.B1(n6572), 
	.B0(\ram[109][8] ), 
	.A1(n6591), 
	.A0(\ram[108][8] ));
   AOI22X1 U9163 (.Y(n11262), 
	.B1(n6610), 
	.B0(\ram[107][8] ), 
	.A1(n6629), 
	.A0(\ram[106][8] ));
   OAI21XL U9164 (.Y(n11232), 
	.B0(n9718), 
	.A1(n11267), 
	.A0(n11266));
   NAND4X1 U9165 (.Y(n11267), 
	.D(n11271), 
	.C(n11270), 
	.B(n11269), 
	.A(n11268));
   AOI22X1 U9166 (.Y(n11271), 
	.B1(n6342), 
	.B0(\ram[89][8] ), 
	.A1(n6362), 
	.A0(\ram[88][8] ));
   AOI22X1 U9167 (.Y(n11270), 
	.B1(n6381), 
	.B0(\ram[87][8] ), 
	.A1(n6400), 
	.A0(\ram[86][8] ));
   AOI22X1 U9168 (.Y(n11269), 
	.B1(n6419), 
	.B0(\ram[85][8] ), 
	.A1(n6438), 
	.A0(\ram[84][8] ));
   AOI22X1 U9169 (.Y(n11268), 
	.B1(n6457), 
	.B0(\ram[83][8] ), 
	.A1(n6476), 
	.A0(\ram[82][8] ));
   NAND4X1 U9170 (.Y(n11266), 
	.D(n11275), 
	.C(n11274), 
	.B(n11273), 
	.A(n11272));
   AOI22X1 U9171 (.Y(n11275), 
	.B1(n6495), 
	.B0(\ram[81][8] ), 
	.A1(n6514), 
	.A0(\ram[80][8] ));
   AOI22X1 U9172 (.Y(n11274), 
	.B1(n6533), 
	.B0(\ram[95][8] ), 
	.A1(n6553), 
	.A0(\ram[94][8] ));
   AOI22X1 U9173 (.Y(n11273), 
	.B1(n6572), 
	.B0(\ram[93][8] ), 
	.A1(n6591), 
	.A0(\ram[92][8] ));
   AOI22X1 U9174 (.Y(n11272), 
	.B1(n6610), 
	.B0(\ram[91][8] ), 
	.A1(n6629), 
	.A0(\ram[90][8] ));
   NAND4X1 U9175 (.Y(n11140), 
	.D(n11279), 
	.C(n11278), 
	.B(n11277), 
	.A(n11276));
   OAI21XL U9176 (.Y(n11279), 
	.B0(n10007), 
	.A1(n11281), 
	.A0(n11280));
   NAND4X1 U9177 (.Y(n11281), 
	.D(n11285), 
	.C(n11284), 
	.B(n11283), 
	.A(n11282));
   AOI22X1 U9178 (.Y(n11285), 
	.B1(n6342), 
	.B0(\ram[73][8] ), 
	.A1(n6362), 
	.A0(\ram[72][8] ));
   AOI22X1 U9179 (.Y(n11284), 
	.B1(n6381), 
	.B0(\ram[71][8] ), 
	.A1(n6400), 
	.A0(\ram[70][8] ));
   AOI22X1 U9180 (.Y(n11283), 
	.B1(n6419), 
	.B0(\ram[69][8] ), 
	.A1(n6438), 
	.A0(\ram[68][8] ));
   AOI22X1 U9181 (.Y(n11282), 
	.B1(n6457), 
	.B0(\ram[67][8] ), 
	.A1(n6476), 
	.A0(\ram[66][8] ));
   NAND4X1 U9182 (.Y(n11280), 
	.D(n11289), 
	.C(n11288), 
	.B(n11287), 
	.A(n11286));
   AOI22X1 U9183 (.Y(n11289), 
	.B1(n6495), 
	.B0(\ram[65][8] ), 
	.A1(n6514), 
	.A0(\ram[64][8] ));
   AOI22X1 U9184 (.Y(n11288), 
	.B1(n6533), 
	.B0(\ram[79][8] ), 
	.A1(n6553), 
	.A0(\ram[78][8] ));
   AOI22X1 U9185 (.Y(n11287), 
	.B1(n6572), 
	.B0(\ram[77][8] ), 
	.A1(n6591), 
	.A0(\ram[76][8] ));
   AOI22X1 U9186 (.Y(n11286), 
	.B1(n6610), 
	.B0(\ram[75][8] ), 
	.A1(n6629), 
	.A0(\ram[74][8] ));
   OAI21XL U9187 (.Y(n11278), 
	.B0(n10296), 
	.A1(n11291), 
	.A0(n11290));
   NAND4X1 U9188 (.Y(n11291), 
	.D(n11295), 
	.C(n11294), 
	.B(n11293), 
	.A(n11292));
   AOI22X1 U9189 (.Y(n11295), 
	.B1(n6342), 
	.B0(\ram[57][8] ), 
	.A1(n6362), 
	.A0(\ram[56][8] ));
   AOI22X1 U9190 (.Y(n11294), 
	.B1(n6381), 
	.B0(\ram[55][8] ), 
	.A1(n6400), 
	.A0(\ram[54][8] ));
   AOI22X1 U9191 (.Y(n11293), 
	.B1(n6419), 
	.B0(\ram[53][8] ), 
	.A1(n6438), 
	.A0(\ram[52][8] ));
   AOI22X1 U9192 (.Y(n11292), 
	.B1(n6457), 
	.B0(\ram[51][8] ), 
	.A1(n6476), 
	.A0(\ram[50][8] ));
   NAND4X1 U9193 (.Y(n11290), 
	.D(n11299), 
	.C(n11298), 
	.B(n11297), 
	.A(n11296));
   AOI22X1 U9194 (.Y(n11299), 
	.B1(n6495), 
	.B0(\ram[49][8] ), 
	.A1(n6514), 
	.A0(\ram[48][8] ));
   AOI22X1 U9195 (.Y(n11298), 
	.B1(n6533), 
	.B0(\ram[63][8] ), 
	.A1(n6553), 
	.A0(\ram[62][8] ));
   AOI22X1 U9196 (.Y(n11297), 
	.B1(n6572), 
	.B0(\ram[61][8] ), 
	.A1(n6591), 
	.A0(\ram[60][8] ));
   AOI22X1 U9197 (.Y(n11296), 
	.B1(n6610), 
	.B0(\ram[59][8] ), 
	.A1(n6629), 
	.A0(\ram[58][8] ));
   OAI21XL U9198 (.Y(n11277), 
	.B0(n10585), 
	.A1(n11301), 
	.A0(n11300));
   NAND4X1 U9199 (.Y(n11301), 
	.D(n11305), 
	.C(n11304), 
	.B(n11303), 
	.A(n11302));
   AOI22X1 U9200 (.Y(n11305), 
	.B1(n6342), 
	.B0(\ram[41][8] ), 
	.A1(n6362), 
	.A0(\ram[40][8] ));
   AOI22X1 U9201 (.Y(n11304), 
	.B1(n6381), 
	.B0(\ram[39][8] ), 
	.A1(n6400), 
	.A0(\ram[38][8] ));
   AOI22X1 U9202 (.Y(n11303), 
	.B1(n6419), 
	.B0(\ram[37][8] ), 
	.A1(n6438), 
	.A0(\ram[36][8] ));
   AOI22X1 U9203 (.Y(n11302), 
	.B1(n6457), 
	.B0(\ram[35][8] ), 
	.A1(n6476), 
	.A0(\ram[34][8] ));
   NAND4X1 U9204 (.Y(n11300), 
	.D(n11309), 
	.C(n11308), 
	.B(n11307), 
	.A(n11306));
   AOI22X1 U9205 (.Y(n11309), 
	.B1(n6495), 
	.B0(\ram[33][8] ), 
	.A1(n6514), 
	.A0(\ram[32][8] ));
   AOI22X1 U9206 (.Y(n11308), 
	.B1(n6533), 
	.B0(\ram[47][8] ), 
	.A1(n6553), 
	.A0(\ram[46][8] ));
   AOI22X1 U9207 (.Y(n11307), 
	.B1(n6572), 
	.B0(\ram[45][8] ), 
	.A1(n6591), 
	.A0(\ram[44][8] ));
   AOI22X1 U9208 (.Y(n11306), 
	.B1(n6610), 
	.B0(\ram[43][8] ), 
	.A1(n6629), 
	.A0(\ram[42][8] ));
   OAI21XL U9209 (.Y(n11276), 
	.B0(n6343), 
	.A1(n11311), 
	.A0(n11310));
   NAND4X1 U9210 (.Y(n11311), 
	.D(n11315), 
	.C(n11314), 
	.B(n11313), 
	.A(n11312));
   AOI22X1 U9211 (.Y(n11315), 
	.B1(n6342), 
	.B0(\ram[25][8] ), 
	.A1(n6362), 
	.A0(\ram[24][8] ));
   AOI22X1 U9212 (.Y(n11314), 
	.B1(n6381), 
	.B0(\ram[23][8] ), 
	.A1(n6400), 
	.A0(\ram[22][8] ));
   AOI22X1 U9213 (.Y(n11313), 
	.B1(n6419), 
	.B0(\ram[21][8] ), 
	.A1(n6438), 
	.A0(\ram[20][8] ));
   AOI22X1 U9214 (.Y(n11312), 
	.B1(n6457), 
	.B0(\ram[19][8] ), 
	.A1(n6476), 
	.A0(\ram[18][8] ));
   NAND4X1 U9215 (.Y(n11310), 
	.D(n11319), 
	.C(n11318), 
	.B(n11317), 
	.A(n11316));
   AOI22X1 U9216 (.Y(n11319), 
	.B1(n6495), 
	.B0(\ram[17][8] ), 
	.A1(n6514), 
	.A0(\ram[16][8] ));
   AOI22X1 U9217 (.Y(n11318), 
	.B1(n6533), 
	.B0(\ram[31][8] ), 
	.A1(n6553), 
	.A0(\ram[30][8] ));
   AOI22X1 U9218 (.Y(n11317), 
	.B1(n6572), 
	.B0(\ram[29][8] ), 
	.A1(n6591), 
	.A0(\ram[28][8] ));
   AOI22X1 U9219 (.Y(n11316), 
	.B1(n6610), 
	.B0(\ram[27][8] ), 
	.A1(n6629), 
	.A0(\ram[26][8] ));
   OR4X1 U9220 (.Y(mem_read_data[7]), 
	.D(n11323), 
	.C(n11322), 
	.B(n11321), 
	.A(n11320));
   NAND4X1 U9221 (.Y(n11323), 
	.D(n11327), 
	.C(n11326), 
	.B(n11325), 
	.A(n11324));
   OAI21XL U9222 (.Y(n11327), 
	.B0(n6534), 
	.A1(n11329), 
	.A0(n11328));
   NAND4X1 U9223 (.Y(n11329), 
	.D(n11333), 
	.C(n11332), 
	.B(n11331), 
	.A(n11330));
   AOI22X1 U9224 (.Y(n11333), 
	.B1(n6342), 
	.B0(\ram[9][7] ), 
	.A1(n6362), 
	.A0(\ram[8][7] ));
   AOI22X1 U9225 (.Y(n11332), 
	.B1(n6381), 
	.B0(\ram[7][7] ), 
	.A1(n6400), 
	.A0(\ram[6][7] ));
   AOI22X1 U9226 (.Y(n11331), 
	.B1(n6419), 
	.B0(\ram[5][7] ), 
	.A1(n6438), 
	.A0(\ram[4][7] ));
   AOI22X1 U9227 (.Y(n11330), 
	.B1(n6457), 
	.B0(\ram[3][7] ), 
	.A1(n6476), 
	.A0(\ram[2][7] ));
   NAND4X1 U9228 (.Y(n11328), 
	.D(n11337), 
	.C(n11336), 
	.B(n11335), 
	.A(n11334));
   AOI22X1 U9229 (.Y(n11337), 
	.B1(n6495), 
	.B0(\ram[1][7] ), 
	.A1(n6514), 
	.A0(\ram[0][7] ));
   AOI22X1 U9230 (.Y(n11336), 
	.B1(n6533), 
	.B0(\ram[15][7] ), 
	.A1(n6553), 
	.A0(\ram[14][7] ));
   AOI22X1 U9231 (.Y(n11335), 
	.B1(n6572), 
	.B0(\ram[13][7] ), 
	.A1(n6591), 
	.A0(\ram[12][7] ));
   AOI22X1 U9232 (.Y(n11334), 
	.B1(n6610), 
	.B0(\ram[11][7] ), 
	.A1(n6629), 
	.A0(\ram[10][7] ));
   OAI21XL U9233 (.Y(n11326), 
	.B0(n6828), 
	.A1(n11339), 
	.A0(n11338));
   NAND4X1 U9234 (.Y(n11339), 
	.D(n11343), 
	.C(n11342), 
	.B(n11341), 
	.A(n11340));
   AOI22X1 U9235 (.Y(n11343), 
	.B1(n6342), 
	.B0(\ram[249][7] ), 
	.A1(n6362), 
	.A0(\ram[248][7] ));
   AOI22X1 U9236 (.Y(n11342), 
	.B1(n6381), 
	.B0(\ram[247][7] ), 
	.A1(n6400), 
	.A0(\ram[246][7] ));
   AOI22X1 U9237 (.Y(n11341), 
	.B1(n6419), 
	.B0(\ram[245][7] ), 
	.A1(n6438), 
	.A0(\ram[244][7] ));
   AOI22X1 U9238 (.Y(n11340), 
	.B1(n6457), 
	.B0(\ram[243][7] ), 
	.A1(n6476), 
	.A0(\ram[242][7] ));
   NAND4X1 U9239 (.Y(n11338), 
	.D(n11347), 
	.C(n11346), 
	.B(n11345), 
	.A(n11344));
   AOI22X1 U9240 (.Y(n11347), 
	.B1(n6495), 
	.B0(\ram[241][7] ), 
	.A1(n6514), 
	.A0(\ram[240][7] ));
   AOI22X1 U9241 (.Y(n11346), 
	.B1(n6533), 
	.B0(\ram[255][7] ), 
	.A1(n6553), 
	.A0(\ram[254][7] ));
   AOI22X1 U9242 (.Y(n11345), 
	.B1(n6572), 
	.B0(\ram[253][7] ), 
	.A1(n6591), 
	.A0(\ram[252][7] ));
   AOI22X1 U9243 (.Y(n11344), 
	.B1(n6610), 
	.B0(\ram[251][7] ), 
	.A1(n6629), 
	.A0(\ram[250][7] ));
   OAI21XL U9244 (.Y(n11325), 
	.B0(n7117), 
	.A1(n11349), 
	.A0(n11348));
   NAND4X1 U9245 (.Y(n11349), 
	.D(n11353), 
	.C(n11352), 
	.B(n11351), 
	.A(n11350));
   AOI22X1 U9246 (.Y(n11353), 
	.B1(n6342), 
	.B0(\ram[233][7] ), 
	.A1(n6362), 
	.A0(\ram[232][7] ));
   AOI22X1 U9247 (.Y(n11352), 
	.B1(n6381), 
	.B0(\ram[231][7] ), 
	.A1(n6400), 
	.A0(\ram[230][7] ));
   AOI22X1 U9248 (.Y(n11351), 
	.B1(n6419), 
	.B0(\ram[229][7] ), 
	.A1(n6438), 
	.A0(\ram[228][7] ));
   AOI22X1 U9249 (.Y(n11350), 
	.B1(n6457), 
	.B0(\ram[227][7] ), 
	.A1(n6476), 
	.A0(\ram[226][7] ));
   NAND4X1 U9250 (.Y(n11348), 
	.D(n11357), 
	.C(n11356), 
	.B(n11355), 
	.A(n11354));
   AOI22X1 U9251 (.Y(n11357), 
	.B1(n6495), 
	.B0(\ram[225][7] ), 
	.A1(n6514), 
	.A0(\ram[224][7] ));
   AOI22X1 U9252 (.Y(n11356), 
	.B1(n6533), 
	.B0(\ram[239][7] ), 
	.A1(n6553), 
	.A0(\ram[238][7] ));
   AOI22X1 U9253 (.Y(n11355), 
	.B1(n6572), 
	.B0(\ram[237][7] ), 
	.A1(n6591), 
	.A0(\ram[236][7] ));
   AOI22X1 U9254 (.Y(n11354), 
	.B1(n6610), 
	.B0(\ram[235][7] ), 
	.A1(n6629), 
	.A0(\ram[234][7] ));
   OAI21XL U9255 (.Y(n11324), 
	.B0(n7406), 
	.A1(n11359), 
	.A0(n11358));
   NAND4X1 U9256 (.Y(n11359), 
	.D(n11363), 
	.C(n11362), 
	.B(n11361), 
	.A(n11360));
   AOI22X1 U9257 (.Y(n11363), 
	.B1(n6342), 
	.B0(\ram[217][7] ), 
	.A1(n6362), 
	.A0(\ram[216][7] ));
   AOI22X1 U9258 (.Y(n11362), 
	.B1(n6381), 
	.B0(\ram[215][7] ), 
	.A1(n6400), 
	.A0(\ram[214][7] ));
   AOI22X1 U9259 (.Y(n11361), 
	.B1(n6419), 
	.B0(\ram[213][7] ), 
	.A1(n6438), 
	.A0(\ram[212][7] ));
   AOI22X1 U9260 (.Y(n11360), 
	.B1(n6457), 
	.B0(\ram[211][7] ), 
	.A1(n6476), 
	.A0(\ram[210][7] ));
   NAND4X1 U9261 (.Y(n11358), 
	.D(n11367), 
	.C(n11366), 
	.B(n11365), 
	.A(n11364));
   AOI22X1 U9262 (.Y(n11367), 
	.B1(n6495), 
	.B0(\ram[209][7] ), 
	.A1(n6514), 
	.A0(\ram[208][7] ));
   AOI22X1 U9263 (.Y(n11366), 
	.B1(n6533), 
	.B0(\ram[223][7] ), 
	.A1(n6553), 
	.A0(\ram[222][7] ));
   AOI22X1 U9264 (.Y(n11365), 
	.B1(n6572), 
	.B0(\ram[221][7] ), 
	.A1(n6591), 
	.A0(\ram[220][7] ));
   AOI22X1 U9265 (.Y(n11364), 
	.B1(n6610), 
	.B0(\ram[219][7] ), 
	.A1(n6629), 
	.A0(\ram[218][7] ));
   NAND4X1 U9266 (.Y(n11322), 
	.D(n11371), 
	.C(n11370), 
	.B(n11369), 
	.A(n11368));
   OAI21XL U9267 (.Y(n11371), 
	.B0(n7695), 
	.A1(n11373), 
	.A0(n11372));
   NAND4X1 U9268 (.Y(n11373), 
	.D(n11377), 
	.C(n11376), 
	.B(n11375), 
	.A(n11374));
   AOI22X1 U9269 (.Y(n11377), 
	.B1(n6342), 
	.B0(\ram[201][7] ), 
	.A1(n6362), 
	.A0(\ram[200][7] ));
   AOI22X1 U9270 (.Y(n11376), 
	.B1(n6381), 
	.B0(\ram[199][7] ), 
	.A1(n6400), 
	.A0(\ram[198][7] ));
   AOI22X1 U9271 (.Y(n11375), 
	.B1(n6419), 
	.B0(\ram[197][7] ), 
	.A1(n6438), 
	.A0(\ram[196][7] ));
   AOI22X1 U9272 (.Y(n11374), 
	.B1(n6457), 
	.B0(\ram[195][7] ), 
	.A1(n6476), 
	.A0(\ram[194][7] ));
   NAND4X1 U9273 (.Y(n11372), 
	.D(n11381), 
	.C(n11380), 
	.B(n11379), 
	.A(n11378));
   AOI22X1 U9274 (.Y(n11381), 
	.B1(n6495), 
	.B0(\ram[193][7] ), 
	.A1(n6514), 
	.A0(\ram[192][7] ));
   AOI22X1 U9275 (.Y(n11380), 
	.B1(n6533), 
	.B0(\ram[207][7] ), 
	.A1(n6553), 
	.A0(\ram[206][7] ));
   AOI22X1 U9276 (.Y(n11379), 
	.B1(n6572), 
	.B0(\ram[205][7] ), 
	.A1(n6591), 
	.A0(\ram[204][7] ));
   AOI22X1 U9277 (.Y(n11378), 
	.B1(n6610), 
	.B0(\ram[203][7] ), 
	.A1(n6629), 
	.A0(\ram[202][7] ));
   OAI21XL U9278 (.Y(n11370), 
	.B0(n7984), 
	.A1(n11383), 
	.A0(n11382));
   NAND4X1 U9279 (.Y(n11383), 
	.D(n11387), 
	.C(n11386), 
	.B(n11385), 
	.A(n11384));
   AOI22X1 U9280 (.Y(n11387), 
	.B1(n6342), 
	.B0(\ram[185][7] ), 
	.A1(n6362), 
	.A0(\ram[184][7] ));
   AOI22X1 U9281 (.Y(n11386), 
	.B1(n6381), 
	.B0(\ram[183][7] ), 
	.A1(n6400), 
	.A0(\ram[182][7] ));
   AOI22X1 U9282 (.Y(n11385), 
	.B1(n6419), 
	.B0(\ram[181][7] ), 
	.A1(n6438), 
	.A0(\ram[180][7] ));
   AOI22X1 U9283 (.Y(n11384), 
	.B1(n6457), 
	.B0(\ram[179][7] ), 
	.A1(n6476), 
	.A0(\ram[178][7] ));
   NAND4X1 U9284 (.Y(n11382), 
	.D(n11391), 
	.C(n11390), 
	.B(n11389), 
	.A(n11388));
   AOI22X1 U9285 (.Y(n11391), 
	.B1(n6495), 
	.B0(\ram[177][7] ), 
	.A1(n6514), 
	.A0(\ram[176][7] ));
   AOI22X1 U9286 (.Y(n11390), 
	.B1(n6533), 
	.B0(\ram[191][7] ), 
	.A1(n6553), 
	.A0(\ram[190][7] ));
   AOI22X1 U9287 (.Y(n11389), 
	.B1(n6572), 
	.B0(\ram[189][7] ), 
	.A1(n6591), 
	.A0(\ram[188][7] ));
   AOI22X1 U9288 (.Y(n11388), 
	.B1(n6610), 
	.B0(\ram[187][7] ), 
	.A1(n6629), 
	.A0(\ram[186][7] ));
   OAI21XL U9289 (.Y(n11369), 
	.B0(n8273), 
	.A1(n11393), 
	.A0(n11392));
   NAND4X1 U9290 (.Y(n11393), 
	.D(n11397), 
	.C(n11396), 
	.B(n11395), 
	.A(n11394));
   AOI22X1 U9291 (.Y(n11397), 
	.B1(n6342), 
	.B0(\ram[169][7] ), 
	.A1(n6362), 
	.A0(\ram[168][7] ));
   AOI22X1 U9292 (.Y(n11396), 
	.B1(n6381), 
	.B0(\ram[167][7] ), 
	.A1(n6400), 
	.A0(\ram[166][7] ));
   AOI22X1 U9293 (.Y(n11395), 
	.B1(n6419), 
	.B0(\ram[165][7] ), 
	.A1(n6438), 
	.A0(\ram[164][7] ));
   AOI22X1 U9294 (.Y(n11394), 
	.B1(n6457), 
	.B0(\ram[163][7] ), 
	.A1(n6476), 
	.A0(\ram[162][7] ));
   NAND4X1 U9295 (.Y(n11392), 
	.D(n11401), 
	.C(n11400), 
	.B(n11399), 
	.A(n11398));
   AOI22X1 U9296 (.Y(n11401), 
	.B1(n6495), 
	.B0(\ram[161][7] ), 
	.A1(n6514), 
	.A0(\ram[160][7] ));
   AOI22X1 U9297 (.Y(n11400), 
	.B1(n6533), 
	.B0(\ram[175][7] ), 
	.A1(n6553), 
	.A0(\ram[174][7] ));
   AOI22X1 U9298 (.Y(n11399), 
	.B1(n6572), 
	.B0(\ram[173][7] ), 
	.A1(n6591), 
	.A0(\ram[172][7] ));
   AOI22X1 U9299 (.Y(n11398), 
	.B1(n6610), 
	.B0(\ram[171][7] ), 
	.A1(n6629), 
	.A0(\ram[170][7] ));
   OAI21XL U9300 (.Y(n11368), 
	.B0(n8562), 
	.A1(n11403), 
	.A0(n11402));
   NAND4X1 U9301 (.Y(n11403), 
	.D(n11407), 
	.C(n11406), 
	.B(n11405), 
	.A(n11404));
   AOI22X1 U9302 (.Y(n11407), 
	.B1(n6342), 
	.B0(\ram[153][7] ), 
	.A1(n6362), 
	.A0(\ram[152][7] ));
   AOI22X1 U9303 (.Y(n11406), 
	.B1(n6381), 
	.B0(\ram[151][7] ), 
	.A1(n6400), 
	.A0(\ram[150][7] ));
   AOI22X1 U9304 (.Y(n11405), 
	.B1(n6419), 
	.B0(\ram[149][7] ), 
	.A1(n6438), 
	.A0(\ram[148][7] ));
   AOI22X1 U9305 (.Y(n11404), 
	.B1(n6457), 
	.B0(\ram[147][7] ), 
	.A1(n6476), 
	.A0(\ram[146][7] ));
   NAND4X1 U9306 (.Y(n11402), 
	.D(n11411), 
	.C(n11410), 
	.B(n11409), 
	.A(n11408));
   AOI22X1 U9307 (.Y(n11411), 
	.B1(n6495), 
	.B0(\ram[145][7] ), 
	.A1(n6514), 
	.A0(\ram[144][7] ));
   AOI22X1 U9308 (.Y(n11410), 
	.B1(n6533), 
	.B0(\ram[159][7] ), 
	.A1(n6553), 
	.A0(\ram[158][7] ));
   AOI22X1 U9309 (.Y(n11409), 
	.B1(n6572), 
	.B0(\ram[157][7] ), 
	.A1(n6591), 
	.A0(\ram[156][7] ));
   AOI22X1 U9310 (.Y(n11408), 
	.B1(n6610), 
	.B0(\ram[155][7] ), 
	.A1(n6629), 
	.A0(\ram[154][7] ));
   NAND4X1 U9311 (.Y(n11321), 
	.D(n11415), 
	.C(n11414), 
	.B(n11413), 
	.A(n11412));
   OAI21XL U9312 (.Y(n11415), 
	.B0(n8851), 
	.A1(n11417), 
	.A0(n11416));
   NAND4X1 U9313 (.Y(n11417), 
	.D(n11421), 
	.C(n11420), 
	.B(n11419), 
	.A(n11418));
   AOI22X1 U9314 (.Y(n11421), 
	.B1(n6342), 
	.B0(\ram[137][7] ), 
	.A1(n6362), 
	.A0(\ram[136][7] ));
   AOI22X1 U9315 (.Y(n11420), 
	.B1(n6381), 
	.B0(\ram[135][7] ), 
	.A1(n6400), 
	.A0(\ram[134][7] ));
   AOI22X1 U9316 (.Y(n11419), 
	.B1(n6419), 
	.B0(\ram[133][7] ), 
	.A1(n6438), 
	.A0(\ram[132][7] ));
   AOI22X1 U9317 (.Y(n11418), 
	.B1(n6457), 
	.B0(\ram[131][7] ), 
	.A1(n6476), 
	.A0(\ram[130][7] ));
   NAND4X1 U9318 (.Y(n11416), 
	.D(n11425), 
	.C(n11424), 
	.B(n11423), 
	.A(n11422));
   AOI22X1 U9319 (.Y(n11425), 
	.B1(n6495), 
	.B0(\ram[129][7] ), 
	.A1(n6514), 
	.A0(\ram[128][7] ));
   AOI22X1 U9320 (.Y(n11424), 
	.B1(n6533), 
	.B0(\ram[143][7] ), 
	.A1(n6553), 
	.A0(\ram[142][7] ));
   AOI22X1 U9321 (.Y(n11423), 
	.B1(n6572), 
	.B0(\ram[141][7] ), 
	.A1(n6591), 
	.A0(\ram[140][7] ));
   AOI22X1 U9322 (.Y(n11422), 
	.B1(n6610), 
	.B0(\ram[139][7] ), 
	.A1(n6629), 
	.A0(\ram[138][7] ));
   OAI21XL U9323 (.Y(n11414), 
	.B0(n9140), 
	.A1(n11427), 
	.A0(n11426));
   NAND4X1 U9324 (.Y(n11427), 
	.D(n11431), 
	.C(n11430), 
	.B(n11429), 
	.A(n11428));
   AOI22X1 U9325 (.Y(n11431), 
	.B1(n6342), 
	.B0(\ram[121][7] ), 
	.A1(n6362), 
	.A0(\ram[120][7] ));
   AOI22X1 U9326 (.Y(n11430), 
	.B1(n6381), 
	.B0(\ram[119][7] ), 
	.A1(n6400), 
	.A0(\ram[118][7] ));
   AOI22X1 U9327 (.Y(n11429), 
	.B1(n6419), 
	.B0(\ram[117][7] ), 
	.A1(n6438), 
	.A0(\ram[116][7] ));
   AOI22X1 U9328 (.Y(n11428), 
	.B1(n6457), 
	.B0(\ram[115][7] ), 
	.A1(n6476), 
	.A0(\ram[114][7] ));
   NAND4X1 U9329 (.Y(n11426), 
	.D(n11435), 
	.C(n11434), 
	.B(n11433), 
	.A(n11432));
   AOI22X1 U9330 (.Y(n11435), 
	.B1(n6495), 
	.B0(\ram[113][7] ), 
	.A1(n6514), 
	.A0(\ram[112][7] ));
   AOI22X1 U9331 (.Y(n11434), 
	.B1(n6533), 
	.B0(\ram[127][7] ), 
	.A1(n6553), 
	.A0(\ram[126][7] ));
   AOI22X1 U9332 (.Y(n11433), 
	.B1(n6572), 
	.B0(\ram[125][7] ), 
	.A1(n6591), 
	.A0(\ram[124][7] ));
   AOI22X1 U9333 (.Y(n11432), 
	.B1(n6610), 
	.B0(\ram[123][7] ), 
	.A1(n6629), 
	.A0(\ram[122][7] ));
   OAI21XL U9334 (.Y(n11413), 
	.B0(n9429), 
	.A1(n11437), 
	.A0(n11436));
   NAND4X1 U9335 (.Y(n11437), 
	.D(n11441), 
	.C(n11440), 
	.B(n11439), 
	.A(n11438));
   AOI22X1 U9336 (.Y(n11441), 
	.B1(n6342), 
	.B0(\ram[105][7] ), 
	.A1(n6362), 
	.A0(\ram[104][7] ));
   AOI22X1 U9337 (.Y(n11440), 
	.B1(n6381), 
	.B0(\ram[103][7] ), 
	.A1(n6400), 
	.A0(\ram[102][7] ));
   AOI22X1 U9338 (.Y(n11439), 
	.B1(n6419), 
	.B0(\ram[101][7] ), 
	.A1(n6438), 
	.A0(\ram[100][7] ));
   AOI22X1 U9339 (.Y(n11438), 
	.B1(n6457), 
	.B0(\ram[99][7] ), 
	.A1(n6476), 
	.A0(\ram[98][7] ));
   NAND4X1 U9340 (.Y(n11436), 
	.D(n11445), 
	.C(n11444), 
	.B(n11443), 
	.A(n11442));
   AOI22X1 U9341 (.Y(n11445), 
	.B1(n6495), 
	.B0(\ram[97][7] ), 
	.A1(n6514), 
	.A0(\ram[96][7] ));
   AOI22X1 U9342 (.Y(n11444), 
	.B1(n6533), 
	.B0(\ram[111][7] ), 
	.A1(n6553), 
	.A0(\ram[110][7] ));
   AOI22X1 U9343 (.Y(n11443), 
	.B1(n6572), 
	.B0(\ram[109][7] ), 
	.A1(n6591), 
	.A0(\ram[108][7] ));
   AOI22X1 U9344 (.Y(n11442), 
	.B1(n6610), 
	.B0(\ram[107][7] ), 
	.A1(n6629), 
	.A0(\ram[106][7] ));
   OAI21XL U9345 (.Y(n11412), 
	.B0(n9718), 
	.A1(n11447), 
	.A0(n11446));
   NAND4X1 U9346 (.Y(n11447), 
	.D(n11451), 
	.C(n11450), 
	.B(n11449), 
	.A(n11448));
   AOI22X1 U9347 (.Y(n11451), 
	.B1(n6342), 
	.B0(\ram[89][7] ), 
	.A1(n6362), 
	.A0(\ram[88][7] ));
   AOI22X1 U9348 (.Y(n11450), 
	.B1(n6381), 
	.B0(\ram[87][7] ), 
	.A1(n6400), 
	.A0(\ram[86][7] ));
   AOI22X1 U9349 (.Y(n11449), 
	.B1(n6419), 
	.B0(\ram[85][7] ), 
	.A1(n6438), 
	.A0(\ram[84][7] ));
   AOI22X1 U9350 (.Y(n11448), 
	.B1(n6457), 
	.B0(\ram[83][7] ), 
	.A1(n6476), 
	.A0(\ram[82][7] ));
   NAND4X1 U9351 (.Y(n11446), 
	.D(n11455), 
	.C(n11454), 
	.B(n11453), 
	.A(n11452));
   AOI22X1 U9352 (.Y(n11455), 
	.B1(n6495), 
	.B0(\ram[81][7] ), 
	.A1(n6514), 
	.A0(\ram[80][7] ));
   AOI22X1 U9353 (.Y(n11454), 
	.B1(n6533), 
	.B0(\ram[95][7] ), 
	.A1(n6553), 
	.A0(\ram[94][7] ));
   AOI22X1 U9354 (.Y(n11453), 
	.B1(n6572), 
	.B0(\ram[93][7] ), 
	.A1(n6591), 
	.A0(\ram[92][7] ));
   AOI22X1 U9355 (.Y(n11452), 
	.B1(n6610), 
	.B0(\ram[91][7] ), 
	.A1(n6629), 
	.A0(\ram[90][7] ));
   NAND4X1 U9356 (.Y(n11320), 
	.D(n11459), 
	.C(n11458), 
	.B(n11457), 
	.A(n11456));
   OAI21XL U9357 (.Y(n11459), 
	.B0(n10007), 
	.A1(n11461), 
	.A0(n11460));
   NAND4X1 U9358 (.Y(n11461), 
	.D(n11465), 
	.C(n11464), 
	.B(n11463), 
	.A(n11462));
   AOI22X1 U9359 (.Y(n11465), 
	.B1(n6342), 
	.B0(\ram[73][7] ), 
	.A1(n6362), 
	.A0(\ram[72][7] ));
   AOI22X1 U9360 (.Y(n11464), 
	.B1(n6381), 
	.B0(\ram[71][7] ), 
	.A1(n6400), 
	.A0(\ram[70][7] ));
   AOI22X1 U9361 (.Y(n11463), 
	.B1(n6419), 
	.B0(\ram[69][7] ), 
	.A1(n6438), 
	.A0(\ram[68][7] ));
   AOI22X1 U9362 (.Y(n11462), 
	.B1(n6457), 
	.B0(\ram[67][7] ), 
	.A1(n6476), 
	.A0(\ram[66][7] ));
   NAND4X1 U9363 (.Y(n11460), 
	.D(n11469), 
	.C(n11468), 
	.B(n11467), 
	.A(n11466));
   AOI22X1 U9364 (.Y(n11469), 
	.B1(n6495), 
	.B0(\ram[65][7] ), 
	.A1(n6514), 
	.A0(\ram[64][7] ));
   AOI22X1 U9365 (.Y(n11468), 
	.B1(n6533), 
	.B0(\ram[79][7] ), 
	.A1(n6553), 
	.A0(\ram[78][7] ));
   AOI22X1 U9366 (.Y(n11467), 
	.B1(n6572), 
	.B0(\ram[77][7] ), 
	.A1(n6591), 
	.A0(\ram[76][7] ));
   AOI22X1 U9367 (.Y(n11466), 
	.B1(n6610), 
	.B0(\ram[75][7] ), 
	.A1(n6629), 
	.A0(\ram[74][7] ));
   OAI21XL U9368 (.Y(n11458), 
	.B0(n10296), 
	.A1(n11471), 
	.A0(n11470));
   NAND4X1 U9369 (.Y(n11471), 
	.D(n11475), 
	.C(n11474), 
	.B(n11473), 
	.A(n11472));
   AOI22X1 U9370 (.Y(n11475), 
	.B1(n6342), 
	.B0(\ram[57][7] ), 
	.A1(n6362), 
	.A0(\ram[56][7] ));
   AOI22X1 U9371 (.Y(n11474), 
	.B1(n6381), 
	.B0(\ram[55][7] ), 
	.A1(n6400), 
	.A0(\ram[54][7] ));
   AOI22X1 U9372 (.Y(n11473), 
	.B1(n6419), 
	.B0(\ram[53][7] ), 
	.A1(n6438), 
	.A0(\ram[52][7] ));
   AOI22X1 U9373 (.Y(n11472), 
	.B1(n6457), 
	.B0(\ram[51][7] ), 
	.A1(n6476), 
	.A0(\ram[50][7] ));
   NAND4X1 U9374 (.Y(n11470), 
	.D(n11479), 
	.C(n11478), 
	.B(n11477), 
	.A(n11476));
   AOI22X1 U9375 (.Y(n11479), 
	.B1(n6495), 
	.B0(\ram[49][7] ), 
	.A1(n6514), 
	.A0(\ram[48][7] ));
   AOI22X1 U9376 (.Y(n11478), 
	.B1(n6533), 
	.B0(\ram[63][7] ), 
	.A1(n6553), 
	.A0(\ram[62][7] ));
   AOI22X1 U9377 (.Y(n11477), 
	.B1(n6572), 
	.B0(\ram[61][7] ), 
	.A1(n6591), 
	.A0(\ram[60][7] ));
   AOI22X1 U9378 (.Y(n11476), 
	.B1(n6610), 
	.B0(\ram[59][7] ), 
	.A1(n6629), 
	.A0(\ram[58][7] ));
   OAI21XL U9379 (.Y(n11457), 
	.B0(n10585), 
	.A1(n11481), 
	.A0(n11480));
   NAND4X1 U9380 (.Y(n11481), 
	.D(n11485), 
	.C(n11484), 
	.B(n11483), 
	.A(n11482));
   AOI22X1 U9381 (.Y(n11485), 
	.B1(n6342), 
	.B0(\ram[41][7] ), 
	.A1(n6362), 
	.A0(\ram[40][7] ));
   AOI22X1 U9382 (.Y(n11484), 
	.B1(n6381), 
	.B0(\ram[39][7] ), 
	.A1(n6400), 
	.A0(\ram[38][7] ));
   AOI22X1 U9383 (.Y(n11483), 
	.B1(n6419), 
	.B0(\ram[37][7] ), 
	.A1(n6438), 
	.A0(\ram[36][7] ));
   AOI22X1 U9384 (.Y(n11482), 
	.B1(n6457), 
	.B0(\ram[35][7] ), 
	.A1(n6476), 
	.A0(\ram[34][7] ));
   NAND4X1 U9385 (.Y(n11480), 
	.D(n11489), 
	.C(n11488), 
	.B(n11487), 
	.A(n11486));
   AOI22X1 U9386 (.Y(n11489), 
	.B1(n6495), 
	.B0(\ram[33][7] ), 
	.A1(n6514), 
	.A0(\ram[32][7] ));
   AOI22X1 U9387 (.Y(n11488), 
	.B1(n6533), 
	.B0(\ram[47][7] ), 
	.A1(n6553), 
	.A0(\ram[46][7] ));
   AOI22X1 U9388 (.Y(n11487), 
	.B1(n6572), 
	.B0(\ram[45][7] ), 
	.A1(n6591), 
	.A0(\ram[44][7] ));
   AOI22X1 U9389 (.Y(n11486), 
	.B1(n6610), 
	.B0(\ram[43][7] ), 
	.A1(n6629), 
	.A0(\ram[42][7] ));
   OAI21XL U9390 (.Y(n11456), 
	.B0(n6343), 
	.A1(n11491), 
	.A0(n11490));
   NAND4X1 U9391 (.Y(n11491), 
	.D(n11495), 
	.C(n11494), 
	.B(n11493), 
	.A(n11492));
   AOI22X1 U9392 (.Y(n11495), 
	.B1(n6342), 
	.B0(\ram[25][7] ), 
	.A1(n6362), 
	.A0(\ram[24][7] ));
   AOI22X1 U9393 (.Y(n11494), 
	.B1(n6381), 
	.B0(\ram[23][7] ), 
	.A1(n6400), 
	.A0(\ram[22][7] ));
   AOI22X1 U9394 (.Y(n11493), 
	.B1(n6419), 
	.B0(\ram[21][7] ), 
	.A1(n6438), 
	.A0(\ram[20][7] ));
   AOI22X1 U9395 (.Y(n11492), 
	.B1(n6457), 
	.B0(\ram[19][7] ), 
	.A1(n6476), 
	.A0(\ram[18][7] ));
   NAND4X1 U9396 (.Y(n11490), 
	.D(n11499), 
	.C(n11498), 
	.B(n11497), 
	.A(n11496));
   AOI22X1 U9397 (.Y(n11499), 
	.B1(n6495), 
	.B0(\ram[17][7] ), 
	.A1(n6514), 
	.A0(\ram[16][7] ));
   AOI22X1 U9398 (.Y(n11498), 
	.B1(n6533), 
	.B0(\ram[31][7] ), 
	.A1(n6553), 
	.A0(\ram[30][7] ));
   AOI22X1 U9399 (.Y(n11497), 
	.B1(n6572), 
	.B0(\ram[29][7] ), 
	.A1(n6591), 
	.A0(\ram[28][7] ));
   AOI22X1 U9400 (.Y(n11496), 
	.B1(n6610), 
	.B0(\ram[27][7] ), 
	.A1(n6629), 
	.A0(\ram[26][7] ));
   OR4X1 U9401 (.Y(mem_read_data[6]), 
	.D(n11503), 
	.C(n11502), 
	.B(n11501), 
	.A(n11500));
   NAND4X1 U9402 (.Y(n11503), 
	.D(n11507), 
	.C(n11506), 
	.B(n11505), 
	.A(n11504));
   OAI21XL U9403 (.Y(n11507), 
	.B0(n6534), 
	.A1(n11509), 
	.A0(n11508));
   NAND4X1 U9404 (.Y(n11509), 
	.D(n11513), 
	.C(n11512), 
	.B(n11511), 
	.A(n11510));
   AOI22X1 U9405 (.Y(n11513), 
	.B1(n6342), 
	.B0(\ram[9][6] ), 
	.A1(n6362), 
	.A0(\ram[8][6] ));
   AOI22X1 U9406 (.Y(n11512), 
	.B1(n6381), 
	.B0(\ram[7][6] ), 
	.A1(n6400), 
	.A0(\ram[6][6] ));
   AOI22X1 U9407 (.Y(n11511), 
	.B1(n6419), 
	.B0(\ram[5][6] ), 
	.A1(n6438), 
	.A0(\ram[4][6] ));
   AOI22X1 U9408 (.Y(n11510), 
	.B1(n6457), 
	.B0(\ram[3][6] ), 
	.A1(n6476), 
	.A0(\ram[2][6] ));
   NAND4X1 U9409 (.Y(n11508), 
	.D(n11517), 
	.C(n11516), 
	.B(n11515), 
	.A(n11514));
   AOI22X1 U9410 (.Y(n11517), 
	.B1(n6495), 
	.B0(\ram[1][6] ), 
	.A1(n6514), 
	.A0(\ram[0][6] ));
   AOI22X1 U9411 (.Y(n11516), 
	.B1(n6533), 
	.B0(\ram[15][6] ), 
	.A1(n6553), 
	.A0(\ram[14][6] ));
   AOI22X1 U9412 (.Y(n11515), 
	.B1(n6572), 
	.B0(\ram[13][6] ), 
	.A1(n6591), 
	.A0(\ram[12][6] ));
   AOI22X1 U9413 (.Y(n11514), 
	.B1(n6610), 
	.B0(\ram[11][6] ), 
	.A1(n6629), 
	.A0(\ram[10][6] ));
   OAI21XL U9414 (.Y(n11506), 
	.B0(n6828), 
	.A1(n11519), 
	.A0(n11518));
   NAND4X1 U9415 (.Y(n11519), 
	.D(n11523), 
	.C(n11522), 
	.B(n11521), 
	.A(n11520));
   AOI22X1 U9416 (.Y(n11523), 
	.B1(n6342), 
	.B0(\ram[249][6] ), 
	.A1(n6362), 
	.A0(\ram[248][6] ));
   AOI22X1 U9417 (.Y(n11522), 
	.B1(n6381), 
	.B0(\ram[247][6] ), 
	.A1(n6400), 
	.A0(\ram[246][6] ));
   AOI22X1 U9418 (.Y(n11521), 
	.B1(n6419), 
	.B0(\ram[245][6] ), 
	.A1(n6438), 
	.A0(\ram[244][6] ));
   AOI22X1 U9419 (.Y(n11520), 
	.B1(n6457), 
	.B0(\ram[243][6] ), 
	.A1(n6476), 
	.A0(\ram[242][6] ));
   NAND4X1 U9420 (.Y(n11518), 
	.D(n11527), 
	.C(n11526), 
	.B(n11525), 
	.A(n11524));
   AOI22X1 U9421 (.Y(n11527), 
	.B1(n6495), 
	.B0(\ram[241][6] ), 
	.A1(n6514), 
	.A0(\ram[240][6] ));
   AOI22X1 U9422 (.Y(n11526), 
	.B1(n6533), 
	.B0(\ram[255][6] ), 
	.A1(n6553), 
	.A0(\ram[254][6] ));
   AOI22X1 U9423 (.Y(n11525), 
	.B1(n6572), 
	.B0(\ram[253][6] ), 
	.A1(n6591), 
	.A0(\ram[252][6] ));
   AOI22X1 U9424 (.Y(n11524), 
	.B1(n6610), 
	.B0(\ram[251][6] ), 
	.A1(n6629), 
	.A0(\ram[250][6] ));
   OAI21XL U9425 (.Y(n11505), 
	.B0(n7117), 
	.A1(n11529), 
	.A0(n11528));
   NAND4X1 U9426 (.Y(n11529), 
	.D(n11533), 
	.C(n11532), 
	.B(n11531), 
	.A(n11530));
   AOI22X1 U9427 (.Y(n11533), 
	.B1(n6342), 
	.B0(\ram[233][6] ), 
	.A1(n6362), 
	.A0(\ram[232][6] ));
   AOI22X1 U9428 (.Y(n11532), 
	.B1(n6381), 
	.B0(\ram[231][6] ), 
	.A1(n6400), 
	.A0(\ram[230][6] ));
   AOI22X1 U9429 (.Y(n11531), 
	.B1(n6419), 
	.B0(\ram[229][6] ), 
	.A1(n6438), 
	.A0(\ram[228][6] ));
   AOI22X1 U9430 (.Y(n11530), 
	.B1(n6457), 
	.B0(\ram[227][6] ), 
	.A1(n6476), 
	.A0(\ram[226][6] ));
   NAND4X1 U9431 (.Y(n11528), 
	.D(n11537), 
	.C(n11536), 
	.B(n11535), 
	.A(n11534));
   AOI22X1 U9432 (.Y(n11537), 
	.B1(n6495), 
	.B0(\ram[225][6] ), 
	.A1(n6514), 
	.A0(\ram[224][6] ));
   AOI22X1 U9433 (.Y(n11536), 
	.B1(n6533), 
	.B0(\ram[239][6] ), 
	.A1(n6553), 
	.A0(\ram[238][6] ));
   AOI22X1 U9434 (.Y(n11535), 
	.B1(n6572), 
	.B0(\ram[237][6] ), 
	.A1(n6591), 
	.A0(\ram[236][6] ));
   AOI22X1 U9435 (.Y(n11534), 
	.B1(n6610), 
	.B0(\ram[235][6] ), 
	.A1(n6629), 
	.A0(\ram[234][6] ));
   OAI21XL U9436 (.Y(n11504), 
	.B0(n7406), 
	.A1(n11539), 
	.A0(n11538));
   NAND4X1 U9437 (.Y(n11539), 
	.D(n11543), 
	.C(n11542), 
	.B(n11541), 
	.A(n11540));
   AOI22X1 U9438 (.Y(n11543), 
	.B1(n6342), 
	.B0(\ram[217][6] ), 
	.A1(n6362), 
	.A0(\ram[216][6] ));
   AOI22X1 U9439 (.Y(n11542), 
	.B1(n6381), 
	.B0(\ram[215][6] ), 
	.A1(n6400), 
	.A0(\ram[214][6] ));
   AOI22X1 U9440 (.Y(n11541), 
	.B1(n6419), 
	.B0(\ram[213][6] ), 
	.A1(n6438), 
	.A0(\ram[212][6] ));
   AOI22X1 U9441 (.Y(n11540), 
	.B1(n6457), 
	.B0(\ram[211][6] ), 
	.A1(n6476), 
	.A0(\ram[210][6] ));
   NAND4X1 U9442 (.Y(n11538), 
	.D(n11547), 
	.C(n11546), 
	.B(n11545), 
	.A(n11544));
   AOI22X1 U9443 (.Y(n11547), 
	.B1(n6495), 
	.B0(\ram[209][6] ), 
	.A1(n6514), 
	.A0(\ram[208][6] ));
   AOI22X1 U9444 (.Y(n11546), 
	.B1(n6533), 
	.B0(\ram[223][6] ), 
	.A1(n6553), 
	.A0(\ram[222][6] ));
   AOI22X1 U9445 (.Y(n11545), 
	.B1(n6572), 
	.B0(\ram[221][6] ), 
	.A1(n6591), 
	.A0(\ram[220][6] ));
   AOI22X1 U9446 (.Y(n11544), 
	.B1(n6610), 
	.B0(\ram[219][6] ), 
	.A1(n6629), 
	.A0(\ram[218][6] ));
   NAND4X1 U9447 (.Y(n11502), 
	.D(n11551), 
	.C(n11550), 
	.B(n11549), 
	.A(n11548));
   OAI21XL U9448 (.Y(n11551), 
	.B0(n7695), 
	.A1(n11553), 
	.A0(n11552));
   NAND4X1 U9449 (.Y(n11553), 
	.D(n11557), 
	.C(n11556), 
	.B(n11555), 
	.A(n11554));
   AOI22X1 U9450 (.Y(n11557), 
	.B1(n6342), 
	.B0(\ram[201][6] ), 
	.A1(n6362), 
	.A0(\ram[200][6] ));
   AOI22X1 U9451 (.Y(n11556), 
	.B1(n6381), 
	.B0(\ram[199][6] ), 
	.A1(n6400), 
	.A0(\ram[198][6] ));
   AOI22X1 U9452 (.Y(n11555), 
	.B1(n6419), 
	.B0(\ram[197][6] ), 
	.A1(n6438), 
	.A0(\ram[196][6] ));
   AOI22X1 U9453 (.Y(n11554), 
	.B1(n6457), 
	.B0(\ram[195][6] ), 
	.A1(n6476), 
	.A0(\ram[194][6] ));
   NAND4X1 U9454 (.Y(n11552), 
	.D(n11561), 
	.C(n11560), 
	.B(n11559), 
	.A(n11558));
   AOI22X1 U9455 (.Y(n11561), 
	.B1(n6495), 
	.B0(\ram[193][6] ), 
	.A1(n6514), 
	.A0(\ram[192][6] ));
   AOI22X1 U9456 (.Y(n11560), 
	.B1(n6533), 
	.B0(\ram[207][6] ), 
	.A1(n6553), 
	.A0(\ram[206][6] ));
   AOI22X1 U9457 (.Y(n11559), 
	.B1(n6572), 
	.B0(\ram[205][6] ), 
	.A1(n6591), 
	.A0(\ram[204][6] ));
   AOI22X1 U9458 (.Y(n11558), 
	.B1(n6610), 
	.B0(\ram[203][6] ), 
	.A1(n6629), 
	.A0(\ram[202][6] ));
   OAI21XL U9459 (.Y(n11550), 
	.B0(n7984), 
	.A1(n11563), 
	.A0(n11562));
   NAND4X1 U9460 (.Y(n11563), 
	.D(n11567), 
	.C(n11566), 
	.B(n11565), 
	.A(n11564));
   AOI22X1 U9461 (.Y(n11567), 
	.B1(n6342), 
	.B0(\ram[185][6] ), 
	.A1(n6362), 
	.A0(\ram[184][6] ));
   AOI22X1 U9462 (.Y(n11566), 
	.B1(n6381), 
	.B0(\ram[183][6] ), 
	.A1(n6400), 
	.A0(\ram[182][6] ));
   AOI22X1 U9463 (.Y(n11565), 
	.B1(n6419), 
	.B0(\ram[181][6] ), 
	.A1(n6438), 
	.A0(\ram[180][6] ));
   AOI22X1 U9464 (.Y(n11564), 
	.B1(n6457), 
	.B0(\ram[179][6] ), 
	.A1(n6476), 
	.A0(\ram[178][6] ));
   NAND4X1 U9465 (.Y(n11562), 
	.D(n11571), 
	.C(n11570), 
	.B(n11569), 
	.A(n11568));
   AOI22X1 U9466 (.Y(n11571), 
	.B1(n6495), 
	.B0(\ram[177][6] ), 
	.A1(n6514), 
	.A0(\ram[176][6] ));
   AOI22X1 U9467 (.Y(n11570), 
	.B1(n6533), 
	.B0(\ram[191][6] ), 
	.A1(n6553), 
	.A0(\ram[190][6] ));
   AOI22X1 U9468 (.Y(n11569), 
	.B1(n6572), 
	.B0(\ram[189][6] ), 
	.A1(n6591), 
	.A0(\ram[188][6] ));
   AOI22X1 U9469 (.Y(n11568), 
	.B1(n6610), 
	.B0(\ram[187][6] ), 
	.A1(n6629), 
	.A0(\ram[186][6] ));
   OAI21XL U9470 (.Y(n11549), 
	.B0(n8273), 
	.A1(n11573), 
	.A0(n11572));
   NAND4X1 U9471 (.Y(n11573), 
	.D(n11577), 
	.C(n11576), 
	.B(n11575), 
	.A(n11574));
   AOI22X1 U9472 (.Y(n11577), 
	.B1(n6342), 
	.B0(\ram[169][6] ), 
	.A1(n6362), 
	.A0(\ram[168][6] ));
   AOI22X1 U9473 (.Y(n11576), 
	.B1(n6381), 
	.B0(\ram[167][6] ), 
	.A1(n6400), 
	.A0(\ram[166][6] ));
   AOI22X1 U9474 (.Y(n11575), 
	.B1(n6419), 
	.B0(\ram[165][6] ), 
	.A1(n6438), 
	.A0(\ram[164][6] ));
   AOI22X1 U9475 (.Y(n11574), 
	.B1(n6457), 
	.B0(\ram[163][6] ), 
	.A1(n6476), 
	.A0(\ram[162][6] ));
   NAND4X1 U9476 (.Y(n11572), 
	.D(n11581), 
	.C(n11580), 
	.B(n11579), 
	.A(n11578));
   AOI22X1 U9477 (.Y(n11581), 
	.B1(n6495), 
	.B0(\ram[161][6] ), 
	.A1(n6514), 
	.A0(\ram[160][6] ));
   AOI22X1 U9478 (.Y(n11580), 
	.B1(n6533), 
	.B0(\ram[175][6] ), 
	.A1(n6553), 
	.A0(\ram[174][6] ));
   AOI22X1 U9479 (.Y(n11579), 
	.B1(n6572), 
	.B0(\ram[173][6] ), 
	.A1(n6591), 
	.A0(\ram[172][6] ));
   AOI22X1 U9480 (.Y(n11578), 
	.B1(n6610), 
	.B0(\ram[171][6] ), 
	.A1(n6629), 
	.A0(\ram[170][6] ));
   OAI21XL U9481 (.Y(n11548), 
	.B0(n8562), 
	.A1(n11583), 
	.A0(n11582));
   NAND4X1 U9482 (.Y(n11583), 
	.D(n11587), 
	.C(n11586), 
	.B(n11585), 
	.A(n11584));
   AOI22X1 U9483 (.Y(n11587), 
	.B1(n6342), 
	.B0(\ram[153][6] ), 
	.A1(n6362), 
	.A0(\ram[152][6] ));
   AOI22X1 U9484 (.Y(n11586), 
	.B1(n6381), 
	.B0(\ram[151][6] ), 
	.A1(n6400), 
	.A0(\ram[150][6] ));
   AOI22X1 U9485 (.Y(n11585), 
	.B1(n6419), 
	.B0(\ram[149][6] ), 
	.A1(n6438), 
	.A0(\ram[148][6] ));
   AOI22X1 U9486 (.Y(n11584), 
	.B1(n6457), 
	.B0(\ram[147][6] ), 
	.A1(n6476), 
	.A0(\ram[146][6] ));
   NAND4X1 U9487 (.Y(n11582), 
	.D(n11591), 
	.C(n11590), 
	.B(n11589), 
	.A(n11588));
   AOI22X1 U9488 (.Y(n11591), 
	.B1(n6495), 
	.B0(\ram[145][6] ), 
	.A1(n6514), 
	.A0(\ram[144][6] ));
   AOI22X1 U9489 (.Y(n11590), 
	.B1(n6533), 
	.B0(\ram[159][6] ), 
	.A1(n6553), 
	.A0(\ram[158][6] ));
   AOI22X1 U9490 (.Y(n11589), 
	.B1(n6572), 
	.B0(\ram[157][6] ), 
	.A1(n6591), 
	.A0(\ram[156][6] ));
   AOI22X1 U9491 (.Y(n11588), 
	.B1(n6610), 
	.B0(\ram[155][6] ), 
	.A1(n6629), 
	.A0(\ram[154][6] ));
   NAND4X1 U9492 (.Y(n11501), 
	.D(n11595), 
	.C(n11594), 
	.B(n11593), 
	.A(n11592));
   OAI21XL U9493 (.Y(n11595), 
	.B0(n8851), 
	.A1(n11597), 
	.A0(n11596));
   NAND4X1 U9494 (.Y(n11597), 
	.D(n11601), 
	.C(n11600), 
	.B(n11599), 
	.A(n11598));
   AOI22X1 U9495 (.Y(n11601), 
	.B1(n6342), 
	.B0(\ram[137][6] ), 
	.A1(n6362), 
	.A0(\ram[136][6] ));
   AOI22X1 U9496 (.Y(n11600), 
	.B1(n6381), 
	.B0(\ram[135][6] ), 
	.A1(n6400), 
	.A0(\ram[134][6] ));
   AOI22X1 U9497 (.Y(n11599), 
	.B1(n6419), 
	.B0(\ram[133][6] ), 
	.A1(n6438), 
	.A0(\ram[132][6] ));
   AOI22X1 U9498 (.Y(n11598), 
	.B1(n6457), 
	.B0(\ram[131][6] ), 
	.A1(n6476), 
	.A0(\ram[130][6] ));
   NAND4X1 U9499 (.Y(n11596), 
	.D(n11605), 
	.C(n11604), 
	.B(n11603), 
	.A(n11602));
   AOI22X1 U9500 (.Y(n11605), 
	.B1(n6495), 
	.B0(\ram[129][6] ), 
	.A1(n6514), 
	.A0(\ram[128][6] ));
   AOI22X1 U9501 (.Y(n11604), 
	.B1(n6533), 
	.B0(\ram[143][6] ), 
	.A1(n6553), 
	.A0(\ram[142][6] ));
   AOI22X1 U9502 (.Y(n11603), 
	.B1(n6572), 
	.B0(\ram[141][6] ), 
	.A1(n6591), 
	.A0(\ram[140][6] ));
   AOI22X1 U9503 (.Y(n11602), 
	.B1(n6610), 
	.B0(\ram[139][6] ), 
	.A1(n6629), 
	.A0(\ram[138][6] ));
   OAI21XL U9504 (.Y(n11594), 
	.B0(n9140), 
	.A1(n11607), 
	.A0(n11606));
   NAND4X1 U9505 (.Y(n11607), 
	.D(n11611), 
	.C(n11610), 
	.B(n11609), 
	.A(n11608));
   AOI22X1 U9506 (.Y(n11611), 
	.B1(n6342), 
	.B0(\ram[121][6] ), 
	.A1(n6362), 
	.A0(\ram[120][6] ));
   AOI22X1 U9507 (.Y(n11610), 
	.B1(n6381), 
	.B0(\ram[119][6] ), 
	.A1(n6400), 
	.A0(\ram[118][6] ));
   AOI22X1 U9508 (.Y(n11609), 
	.B1(n6419), 
	.B0(\ram[117][6] ), 
	.A1(n6438), 
	.A0(\ram[116][6] ));
   AOI22X1 U9509 (.Y(n11608), 
	.B1(n6457), 
	.B0(\ram[115][6] ), 
	.A1(n6476), 
	.A0(\ram[114][6] ));
   NAND4X1 U9510 (.Y(n11606), 
	.D(n11615), 
	.C(n11614), 
	.B(n11613), 
	.A(n11612));
   AOI22X1 U9511 (.Y(n11615), 
	.B1(n6495), 
	.B0(\ram[113][6] ), 
	.A1(n6514), 
	.A0(\ram[112][6] ));
   AOI22X1 U9512 (.Y(n11614), 
	.B1(n6533), 
	.B0(\ram[127][6] ), 
	.A1(n6553), 
	.A0(\ram[126][6] ));
   AOI22X1 U9513 (.Y(n11613), 
	.B1(n6572), 
	.B0(\ram[125][6] ), 
	.A1(n6591), 
	.A0(\ram[124][6] ));
   AOI22X1 U9514 (.Y(n11612), 
	.B1(n6610), 
	.B0(\ram[123][6] ), 
	.A1(n6629), 
	.A0(\ram[122][6] ));
   OAI21XL U9515 (.Y(n11593), 
	.B0(n9429), 
	.A1(n11617), 
	.A0(n11616));
   NAND4X1 U9516 (.Y(n11617), 
	.D(n11621), 
	.C(n11620), 
	.B(n11619), 
	.A(n11618));
   AOI22X1 U9517 (.Y(n11621), 
	.B1(n6342), 
	.B0(\ram[105][6] ), 
	.A1(n6362), 
	.A0(\ram[104][6] ));
   AOI22X1 U9518 (.Y(n11620), 
	.B1(n6381), 
	.B0(\ram[103][6] ), 
	.A1(n6400), 
	.A0(\ram[102][6] ));
   AOI22X1 U9519 (.Y(n11619), 
	.B1(n6419), 
	.B0(\ram[101][6] ), 
	.A1(n6438), 
	.A0(\ram[100][6] ));
   AOI22X1 U9520 (.Y(n11618), 
	.B1(n6457), 
	.B0(\ram[99][6] ), 
	.A1(n6476), 
	.A0(\ram[98][6] ));
   NAND4X1 U9521 (.Y(n11616), 
	.D(n11625), 
	.C(n11624), 
	.B(n11623), 
	.A(n11622));
   AOI22X1 U9522 (.Y(n11625), 
	.B1(n6495), 
	.B0(\ram[97][6] ), 
	.A1(n6514), 
	.A0(\ram[96][6] ));
   AOI22X1 U9523 (.Y(n11624), 
	.B1(n6533), 
	.B0(\ram[111][6] ), 
	.A1(n6553), 
	.A0(\ram[110][6] ));
   AOI22X1 U9524 (.Y(n11623), 
	.B1(n6572), 
	.B0(\ram[109][6] ), 
	.A1(n6591), 
	.A0(\ram[108][6] ));
   AOI22X1 U9525 (.Y(n11622), 
	.B1(n6610), 
	.B0(\ram[107][6] ), 
	.A1(n6629), 
	.A0(\ram[106][6] ));
   OAI21XL U9526 (.Y(n11592), 
	.B0(n9718), 
	.A1(n11627), 
	.A0(n11626));
   NAND4X1 U9527 (.Y(n11627), 
	.D(n11631), 
	.C(n11630), 
	.B(n11629), 
	.A(n11628));
   AOI22X1 U9528 (.Y(n11631), 
	.B1(n6342), 
	.B0(\ram[89][6] ), 
	.A1(n6362), 
	.A0(\ram[88][6] ));
   AOI22X1 U9529 (.Y(n11630), 
	.B1(n6381), 
	.B0(\ram[87][6] ), 
	.A1(n6400), 
	.A0(\ram[86][6] ));
   AOI22X1 U9530 (.Y(n11629), 
	.B1(n6419), 
	.B0(\ram[85][6] ), 
	.A1(n6438), 
	.A0(\ram[84][6] ));
   AOI22X1 U9531 (.Y(n11628), 
	.B1(n6457), 
	.B0(\ram[83][6] ), 
	.A1(n6476), 
	.A0(\ram[82][6] ));
   NAND4X1 U9532 (.Y(n11626), 
	.D(n11635), 
	.C(n11634), 
	.B(n11633), 
	.A(n11632));
   AOI22X1 U9533 (.Y(n11635), 
	.B1(n6495), 
	.B0(\ram[81][6] ), 
	.A1(n6514), 
	.A0(\ram[80][6] ));
   AOI22X1 U9534 (.Y(n11634), 
	.B1(n6533), 
	.B0(\ram[95][6] ), 
	.A1(n6553), 
	.A0(\ram[94][6] ));
   AOI22X1 U9535 (.Y(n11633), 
	.B1(n6572), 
	.B0(\ram[93][6] ), 
	.A1(n6591), 
	.A0(\ram[92][6] ));
   AOI22X1 U9536 (.Y(n11632), 
	.B1(n6610), 
	.B0(\ram[91][6] ), 
	.A1(n6629), 
	.A0(\ram[90][6] ));
   NAND4X1 U9537 (.Y(n11500), 
	.D(n11639), 
	.C(n11638), 
	.B(n11637), 
	.A(n11636));
   OAI21XL U9538 (.Y(n11639), 
	.B0(n10007), 
	.A1(n11641), 
	.A0(n11640));
   NAND4X1 U9539 (.Y(n11641), 
	.D(n11645), 
	.C(n11644), 
	.B(n11643), 
	.A(n11642));
   AOI22X1 U9540 (.Y(n11645), 
	.B1(n6342), 
	.B0(\ram[73][6] ), 
	.A1(n6362), 
	.A0(\ram[72][6] ));
   AOI22X1 U9541 (.Y(n11644), 
	.B1(n6381), 
	.B0(\ram[71][6] ), 
	.A1(n6400), 
	.A0(\ram[70][6] ));
   AOI22X1 U9542 (.Y(n11643), 
	.B1(n6419), 
	.B0(\ram[69][6] ), 
	.A1(n6438), 
	.A0(\ram[68][6] ));
   AOI22X1 U9543 (.Y(n11642), 
	.B1(n6457), 
	.B0(\ram[67][6] ), 
	.A1(n6476), 
	.A0(\ram[66][6] ));
   NAND4X1 U9544 (.Y(n11640), 
	.D(n11649), 
	.C(n11648), 
	.B(n11647), 
	.A(n11646));
   AOI22X1 U9545 (.Y(n11649), 
	.B1(n6495), 
	.B0(\ram[65][6] ), 
	.A1(n6514), 
	.A0(\ram[64][6] ));
   AOI22X1 U9546 (.Y(n11648), 
	.B1(n6533), 
	.B0(\ram[79][6] ), 
	.A1(n6553), 
	.A0(\ram[78][6] ));
   AOI22X1 U9547 (.Y(n11647), 
	.B1(n6572), 
	.B0(\ram[77][6] ), 
	.A1(n6591), 
	.A0(\ram[76][6] ));
   AOI22X1 U9548 (.Y(n11646), 
	.B1(n6610), 
	.B0(\ram[75][6] ), 
	.A1(n6629), 
	.A0(\ram[74][6] ));
   OAI21XL U9549 (.Y(n11638), 
	.B0(n10296), 
	.A1(n11651), 
	.A0(n11650));
   NAND4X1 U9550 (.Y(n11651), 
	.D(n11655), 
	.C(n11654), 
	.B(n11653), 
	.A(n11652));
   AOI22X1 U9551 (.Y(n11655), 
	.B1(n6342), 
	.B0(\ram[57][6] ), 
	.A1(n6362), 
	.A0(\ram[56][6] ));
   AOI22X1 U9552 (.Y(n11654), 
	.B1(n6381), 
	.B0(\ram[55][6] ), 
	.A1(n6400), 
	.A0(\ram[54][6] ));
   AOI22X1 U9553 (.Y(n11653), 
	.B1(n6419), 
	.B0(\ram[53][6] ), 
	.A1(n6438), 
	.A0(\ram[52][6] ));
   AOI22X1 U9554 (.Y(n11652), 
	.B1(n6457), 
	.B0(\ram[51][6] ), 
	.A1(n6476), 
	.A0(\ram[50][6] ));
   NAND4X1 U9555 (.Y(n11650), 
	.D(n11659), 
	.C(n11658), 
	.B(n11657), 
	.A(n11656));
   AOI22X1 U9556 (.Y(n11659), 
	.B1(n6495), 
	.B0(\ram[49][6] ), 
	.A1(n6514), 
	.A0(\ram[48][6] ));
   AOI22X1 U9557 (.Y(n11658), 
	.B1(n6533), 
	.B0(\ram[63][6] ), 
	.A1(n6553), 
	.A0(\ram[62][6] ));
   AOI22X1 U9558 (.Y(n11657), 
	.B1(n6572), 
	.B0(\ram[61][6] ), 
	.A1(n6591), 
	.A0(\ram[60][6] ));
   AOI22X1 U9559 (.Y(n11656), 
	.B1(n6610), 
	.B0(\ram[59][6] ), 
	.A1(n6629), 
	.A0(\ram[58][6] ));
   OAI21XL U9560 (.Y(n11637), 
	.B0(n10585), 
	.A1(n11661), 
	.A0(n11660));
   NAND4X1 U9561 (.Y(n11661), 
	.D(n11665), 
	.C(n11664), 
	.B(n11663), 
	.A(n11662));
   AOI22X1 U9562 (.Y(n11665), 
	.B1(n6342), 
	.B0(\ram[41][6] ), 
	.A1(n6362), 
	.A0(\ram[40][6] ));
   AOI22X1 U9563 (.Y(n11664), 
	.B1(n6381), 
	.B0(\ram[39][6] ), 
	.A1(n6400), 
	.A0(\ram[38][6] ));
   AOI22X1 U9564 (.Y(n11663), 
	.B1(n6419), 
	.B0(\ram[37][6] ), 
	.A1(n6438), 
	.A0(\ram[36][6] ));
   AOI22X1 U9565 (.Y(n11662), 
	.B1(n6457), 
	.B0(\ram[35][6] ), 
	.A1(n6476), 
	.A0(\ram[34][6] ));
   NAND4X1 U9566 (.Y(n11660), 
	.D(n11669), 
	.C(n11668), 
	.B(n11667), 
	.A(n11666));
   AOI22X1 U9567 (.Y(n11669), 
	.B1(n6495), 
	.B0(\ram[33][6] ), 
	.A1(n6514), 
	.A0(\ram[32][6] ));
   AOI22X1 U9568 (.Y(n11668), 
	.B1(n6533), 
	.B0(\ram[47][6] ), 
	.A1(n6553), 
	.A0(\ram[46][6] ));
   AOI22X1 U9569 (.Y(n11667), 
	.B1(n6572), 
	.B0(\ram[45][6] ), 
	.A1(n6591), 
	.A0(\ram[44][6] ));
   AOI22X1 U9570 (.Y(n11666), 
	.B1(n6610), 
	.B0(\ram[43][6] ), 
	.A1(n6629), 
	.A0(\ram[42][6] ));
   OAI21XL U9571 (.Y(n11636), 
	.B0(n6343), 
	.A1(n11671), 
	.A0(n11670));
   NAND4X1 U9572 (.Y(n11671), 
	.D(n11675), 
	.C(n11674), 
	.B(n11673), 
	.A(n11672));
   AOI22X1 U9573 (.Y(n11675), 
	.B1(n6342), 
	.B0(\ram[25][6] ), 
	.A1(n6362), 
	.A0(\ram[24][6] ));
   AOI22X1 U9574 (.Y(n11674), 
	.B1(n6381), 
	.B0(\ram[23][6] ), 
	.A1(n6400), 
	.A0(\ram[22][6] ));
   AOI22X1 U9575 (.Y(n11673), 
	.B1(n6419), 
	.B0(\ram[21][6] ), 
	.A1(n6438), 
	.A0(\ram[20][6] ));
   AOI22X1 U9576 (.Y(n11672), 
	.B1(n6457), 
	.B0(\ram[19][6] ), 
	.A1(n6476), 
	.A0(\ram[18][6] ));
   NAND4X1 U9577 (.Y(n11670), 
	.D(n11679), 
	.C(n11678), 
	.B(n11677), 
	.A(n11676));
   AOI22X1 U9578 (.Y(n11679), 
	.B1(n6495), 
	.B0(\ram[17][6] ), 
	.A1(n6514), 
	.A0(\ram[16][6] ));
   AOI22X1 U9579 (.Y(n11678), 
	.B1(n6533), 
	.B0(\ram[31][6] ), 
	.A1(n6553), 
	.A0(\ram[30][6] ));
   AOI22X1 U9580 (.Y(n11677), 
	.B1(n6572), 
	.B0(\ram[29][6] ), 
	.A1(n6591), 
	.A0(\ram[28][6] ));
   AOI22X1 U9581 (.Y(n11676), 
	.B1(n6610), 
	.B0(\ram[27][6] ), 
	.A1(n6629), 
	.A0(\ram[26][6] ));
   OR4X1 U9582 (.Y(mem_read_data[5]), 
	.D(n11683), 
	.C(n11682), 
	.B(n11681), 
	.A(n11680));
   NAND4X1 U9583 (.Y(n11683), 
	.D(n11687), 
	.C(n11686), 
	.B(n11685), 
	.A(n11684));
   OAI21XL U9584 (.Y(n11687), 
	.B0(n6534), 
	.A1(n11689), 
	.A0(n11688));
   NAND4X1 U9585 (.Y(n11689), 
	.D(n11693), 
	.C(n11692), 
	.B(n11691), 
	.A(n11690));
   AOI22X1 U9586 (.Y(n11693), 
	.B1(n6342), 
	.B0(\ram[9][5] ), 
	.A1(n6362), 
	.A0(\ram[8][5] ));
   AOI22X1 U9587 (.Y(n11692), 
	.B1(n6381), 
	.B0(\ram[7][5] ), 
	.A1(n6400), 
	.A0(\ram[6][5] ));
   AOI22X1 U9588 (.Y(n11691), 
	.B1(n6419), 
	.B0(\ram[5][5] ), 
	.A1(n6438), 
	.A0(\ram[4][5] ));
   AOI22X1 U9589 (.Y(n11690), 
	.B1(n6457), 
	.B0(\ram[3][5] ), 
	.A1(n6476), 
	.A0(\ram[2][5] ));
   NAND4X1 U9590 (.Y(n11688), 
	.D(n11697), 
	.C(n11696), 
	.B(n11695), 
	.A(n11694));
   AOI22X1 U9591 (.Y(n11697), 
	.B1(n6495), 
	.B0(\ram[1][5] ), 
	.A1(n6514), 
	.A0(\ram[0][5] ));
   AOI22X1 U9592 (.Y(n11696), 
	.B1(n6533), 
	.B0(\ram[15][5] ), 
	.A1(n6553), 
	.A0(\ram[14][5] ));
   AOI22X1 U9593 (.Y(n11695), 
	.B1(n6572), 
	.B0(\ram[13][5] ), 
	.A1(n6591), 
	.A0(\ram[12][5] ));
   AOI22X1 U9594 (.Y(n11694), 
	.B1(n6610), 
	.B0(\ram[11][5] ), 
	.A1(n6629), 
	.A0(\ram[10][5] ));
   OAI21XL U9595 (.Y(n11686), 
	.B0(n6828), 
	.A1(n11699), 
	.A0(n11698));
   NAND4X1 U9596 (.Y(n11699), 
	.D(n11703), 
	.C(n11702), 
	.B(n11701), 
	.A(n11700));
   AOI22X1 U9597 (.Y(n11703), 
	.B1(n6342), 
	.B0(\ram[249][5] ), 
	.A1(n6362), 
	.A0(\ram[248][5] ));
   AOI22X1 U9598 (.Y(n11702), 
	.B1(n6381), 
	.B0(\ram[247][5] ), 
	.A1(n6400), 
	.A0(\ram[246][5] ));
   AOI22X1 U9599 (.Y(n11701), 
	.B1(n6419), 
	.B0(\ram[245][5] ), 
	.A1(n6438), 
	.A0(\ram[244][5] ));
   AOI22X1 U9600 (.Y(n11700), 
	.B1(n6457), 
	.B0(\ram[243][5] ), 
	.A1(n6476), 
	.A0(\ram[242][5] ));
   NAND4X1 U9601 (.Y(n11698), 
	.D(n11707), 
	.C(n11706), 
	.B(n11705), 
	.A(n11704));
   AOI22X1 U9602 (.Y(n11707), 
	.B1(n6495), 
	.B0(\ram[241][5] ), 
	.A1(n6514), 
	.A0(\ram[240][5] ));
   AOI22X1 U9603 (.Y(n11706), 
	.B1(n6533), 
	.B0(\ram[255][5] ), 
	.A1(n6553), 
	.A0(\ram[254][5] ));
   AOI22X1 U9604 (.Y(n11705), 
	.B1(n6572), 
	.B0(\ram[253][5] ), 
	.A1(n6591), 
	.A0(\ram[252][5] ));
   AOI22X1 U9605 (.Y(n11704), 
	.B1(n6610), 
	.B0(\ram[251][5] ), 
	.A1(n6629), 
	.A0(\ram[250][5] ));
   OAI21XL U9606 (.Y(n11685), 
	.B0(n7117), 
	.A1(n11709), 
	.A0(n11708));
   NAND4X1 U9607 (.Y(n11709), 
	.D(n11713), 
	.C(n11712), 
	.B(n11711), 
	.A(n11710));
   AOI22X1 U9608 (.Y(n11713), 
	.B1(n6342), 
	.B0(\ram[233][5] ), 
	.A1(n6362), 
	.A0(\ram[232][5] ));
   AOI22X1 U9609 (.Y(n11712), 
	.B1(n6381), 
	.B0(\ram[231][5] ), 
	.A1(n6400), 
	.A0(\ram[230][5] ));
   AOI22X1 U9610 (.Y(n11711), 
	.B1(n6419), 
	.B0(\ram[229][5] ), 
	.A1(n6438), 
	.A0(\ram[228][5] ));
   AOI22X1 U9611 (.Y(n11710), 
	.B1(n6457), 
	.B0(\ram[227][5] ), 
	.A1(n6476), 
	.A0(\ram[226][5] ));
   NAND4X1 U9612 (.Y(n11708), 
	.D(n11717), 
	.C(n11716), 
	.B(n11715), 
	.A(n11714));
   AOI22X1 U9613 (.Y(n11717), 
	.B1(n6495), 
	.B0(\ram[225][5] ), 
	.A1(n6514), 
	.A0(\ram[224][5] ));
   AOI22X1 U9614 (.Y(n11716), 
	.B1(n6533), 
	.B0(\ram[239][5] ), 
	.A1(n6553), 
	.A0(\ram[238][5] ));
   AOI22X1 U9615 (.Y(n11715), 
	.B1(n6572), 
	.B0(\ram[237][5] ), 
	.A1(n6591), 
	.A0(\ram[236][5] ));
   AOI22X1 U9616 (.Y(n11714), 
	.B1(n6610), 
	.B0(\ram[235][5] ), 
	.A1(n6629), 
	.A0(\ram[234][5] ));
   OAI21XL U9617 (.Y(n11684), 
	.B0(n7406), 
	.A1(n11719), 
	.A0(n11718));
   NAND4X1 U9618 (.Y(n11719), 
	.D(n11723), 
	.C(n11722), 
	.B(n11721), 
	.A(n11720));
   AOI22X1 U9619 (.Y(n11723), 
	.B1(n6342), 
	.B0(\ram[217][5] ), 
	.A1(n6362), 
	.A0(\ram[216][5] ));
   AOI22X1 U9620 (.Y(n11722), 
	.B1(n6381), 
	.B0(\ram[215][5] ), 
	.A1(n6400), 
	.A0(\ram[214][5] ));
   AOI22X1 U9621 (.Y(n11721), 
	.B1(n6419), 
	.B0(\ram[213][5] ), 
	.A1(n6438), 
	.A0(\ram[212][5] ));
   AOI22X1 U9622 (.Y(n11720), 
	.B1(n6457), 
	.B0(\ram[211][5] ), 
	.A1(n6476), 
	.A0(\ram[210][5] ));
   NAND4X1 U9623 (.Y(n11718), 
	.D(n11727), 
	.C(n11726), 
	.B(n11725), 
	.A(n11724));
   AOI22X1 U9624 (.Y(n11727), 
	.B1(n6495), 
	.B0(\ram[209][5] ), 
	.A1(n6514), 
	.A0(\ram[208][5] ));
   AOI22X1 U9625 (.Y(n11726), 
	.B1(n6533), 
	.B0(\ram[223][5] ), 
	.A1(n6553), 
	.A0(\ram[222][5] ));
   AOI22X1 U9626 (.Y(n11725), 
	.B1(n6572), 
	.B0(\ram[221][5] ), 
	.A1(n6591), 
	.A0(\ram[220][5] ));
   AOI22X1 U9627 (.Y(n11724), 
	.B1(n6610), 
	.B0(\ram[219][5] ), 
	.A1(n6629), 
	.A0(\ram[218][5] ));
   NAND4X1 U9628 (.Y(n11682), 
	.D(n11731), 
	.C(n11730), 
	.B(n11729), 
	.A(n11728));
   OAI21XL U9629 (.Y(n11731), 
	.B0(n7695), 
	.A1(n11733), 
	.A0(n11732));
   NAND4X1 U9630 (.Y(n11733), 
	.D(n11737), 
	.C(n11736), 
	.B(n11735), 
	.A(n11734));
   AOI22X1 U9631 (.Y(n11737), 
	.B1(n6342), 
	.B0(\ram[201][5] ), 
	.A1(n6362), 
	.A0(\ram[200][5] ));
   AOI22X1 U9632 (.Y(n11736), 
	.B1(n6381), 
	.B0(\ram[199][5] ), 
	.A1(n6400), 
	.A0(\ram[198][5] ));
   AOI22X1 U9633 (.Y(n11735), 
	.B1(n6419), 
	.B0(\ram[197][5] ), 
	.A1(n6438), 
	.A0(\ram[196][5] ));
   AOI22X1 U9634 (.Y(n11734), 
	.B1(n6457), 
	.B0(\ram[195][5] ), 
	.A1(n6476), 
	.A0(\ram[194][5] ));
   NAND4X1 U9635 (.Y(n11732), 
	.D(n11741), 
	.C(n11740), 
	.B(n11739), 
	.A(n11738));
   AOI22X1 U9636 (.Y(n11741), 
	.B1(n6495), 
	.B0(\ram[193][5] ), 
	.A1(n6514), 
	.A0(\ram[192][5] ));
   AOI22X1 U9637 (.Y(n11740), 
	.B1(n6533), 
	.B0(\ram[207][5] ), 
	.A1(n6553), 
	.A0(\ram[206][5] ));
   AOI22X1 U9638 (.Y(n11739), 
	.B1(n6572), 
	.B0(\ram[205][5] ), 
	.A1(n6591), 
	.A0(\ram[204][5] ));
   AOI22X1 U9639 (.Y(n11738), 
	.B1(n6610), 
	.B0(\ram[203][5] ), 
	.A1(n6629), 
	.A0(\ram[202][5] ));
   OAI21XL U9640 (.Y(n11730), 
	.B0(n7984), 
	.A1(n11743), 
	.A0(n11742));
   NAND4X1 U9641 (.Y(n11743), 
	.D(n11747), 
	.C(n11746), 
	.B(n11745), 
	.A(n11744));
   AOI22X1 U9642 (.Y(n11747), 
	.B1(n6342), 
	.B0(\ram[185][5] ), 
	.A1(n6362), 
	.A0(\ram[184][5] ));
   AOI22X1 U9643 (.Y(n11746), 
	.B1(n6381), 
	.B0(\ram[183][5] ), 
	.A1(n6400), 
	.A0(\ram[182][5] ));
   AOI22X1 U9644 (.Y(n11745), 
	.B1(n6419), 
	.B0(\ram[181][5] ), 
	.A1(n6438), 
	.A0(\ram[180][5] ));
   AOI22X1 U9645 (.Y(n11744), 
	.B1(n6457), 
	.B0(\ram[179][5] ), 
	.A1(n6476), 
	.A0(\ram[178][5] ));
   NAND4X1 U9646 (.Y(n11742), 
	.D(n11751), 
	.C(n11750), 
	.B(n11749), 
	.A(n11748));
   AOI22X1 U9647 (.Y(n11751), 
	.B1(n6495), 
	.B0(\ram[177][5] ), 
	.A1(n6514), 
	.A0(\ram[176][5] ));
   AOI22X1 U9648 (.Y(n11750), 
	.B1(n6533), 
	.B0(\ram[191][5] ), 
	.A1(n6553), 
	.A0(\ram[190][5] ));
   AOI22X1 U9649 (.Y(n11749), 
	.B1(n6572), 
	.B0(\ram[189][5] ), 
	.A1(n6591), 
	.A0(\ram[188][5] ));
   AOI22X1 U9650 (.Y(n11748), 
	.B1(n6610), 
	.B0(\ram[187][5] ), 
	.A1(n6629), 
	.A0(\ram[186][5] ));
   OAI21XL U9651 (.Y(n11729), 
	.B0(n8273), 
	.A1(n11753), 
	.A0(n11752));
   NAND4X1 U9652 (.Y(n11753), 
	.D(n11757), 
	.C(n11756), 
	.B(n11755), 
	.A(n11754));
   AOI22X1 U9653 (.Y(n11757), 
	.B1(n6342), 
	.B0(\ram[169][5] ), 
	.A1(n6362), 
	.A0(\ram[168][5] ));
   AOI22X1 U9654 (.Y(n11756), 
	.B1(n6381), 
	.B0(\ram[167][5] ), 
	.A1(n6400), 
	.A0(\ram[166][5] ));
   AOI22X1 U9655 (.Y(n11755), 
	.B1(n6419), 
	.B0(\ram[165][5] ), 
	.A1(n6438), 
	.A0(\ram[164][5] ));
   AOI22X1 U9656 (.Y(n11754), 
	.B1(n6457), 
	.B0(\ram[163][5] ), 
	.A1(n6476), 
	.A0(\ram[162][5] ));
   NAND4X1 U9657 (.Y(n11752), 
	.D(n11761), 
	.C(n11760), 
	.B(n11759), 
	.A(n11758));
   AOI22X1 U9658 (.Y(n11761), 
	.B1(n6495), 
	.B0(\ram[161][5] ), 
	.A1(n6514), 
	.A0(\ram[160][5] ));
   AOI22X1 U9659 (.Y(n11760), 
	.B1(n6533), 
	.B0(\ram[175][5] ), 
	.A1(n6553), 
	.A0(\ram[174][5] ));
   AOI22X1 U9660 (.Y(n11759), 
	.B1(n6572), 
	.B0(\ram[173][5] ), 
	.A1(n6591), 
	.A0(\ram[172][5] ));
   AOI22X1 U9661 (.Y(n11758), 
	.B1(n6610), 
	.B0(\ram[171][5] ), 
	.A1(n6629), 
	.A0(\ram[170][5] ));
   OAI21XL U9662 (.Y(n11728), 
	.B0(n8562), 
	.A1(n11763), 
	.A0(n11762));
   NAND4X1 U9663 (.Y(n11763), 
	.D(n11767), 
	.C(n11766), 
	.B(n11765), 
	.A(n11764));
   AOI22X1 U9664 (.Y(n11767), 
	.B1(n6342), 
	.B0(\ram[153][5] ), 
	.A1(n6362), 
	.A0(\ram[152][5] ));
   AOI22X1 U9665 (.Y(n11766), 
	.B1(n6381), 
	.B0(\ram[151][5] ), 
	.A1(n6400), 
	.A0(\ram[150][5] ));
   AOI22X1 U9666 (.Y(n11765), 
	.B1(n6419), 
	.B0(\ram[149][5] ), 
	.A1(n6438), 
	.A0(\ram[148][5] ));
   AOI22X1 U9667 (.Y(n11764), 
	.B1(n6457), 
	.B0(\ram[147][5] ), 
	.A1(n6476), 
	.A0(\ram[146][5] ));
   NAND4X1 U9668 (.Y(n11762), 
	.D(n11771), 
	.C(n11770), 
	.B(n11769), 
	.A(n11768));
   AOI22X1 U9669 (.Y(n11771), 
	.B1(n6495), 
	.B0(\ram[145][5] ), 
	.A1(n6514), 
	.A0(\ram[144][5] ));
   AOI22X1 U9670 (.Y(n11770), 
	.B1(n6533), 
	.B0(\ram[159][5] ), 
	.A1(n6553), 
	.A0(\ram[158][5] ));
   AOI22X1 U9671 (.Y(n11769), 
	.B1(n6572), 
	.B0(\ram[157][5] ), 
	.A1(n6591), 
	.A0(\ram[156][5] ));
   AOI22X1 U9672 (.Y(n11768), 
	.B1(n6610), 
	.B0(\ram[155][5] ), 
	.A1(n6629), 
	.A0(\ram[154][5] ));
   NAND4X1 U9673 (.Y(n11681), 
	.D(n11775), 
	.C(n11774), 
	.B(n11773), 
	.A(n11772));
   OAI21XL U9674 (.Y(n11775), 
	.B0(n8851), 
	.A1(n11777), 
	.A0(n11776));
   NAND4X1 U9675 (.Y(n11777), 
	.D(n11781), 
	.C(n11780), 
	.B(n11779), 
	.A(n11778));
   AOI22X1 U9676 (.Y(n11781), 
	.B1(n6342), 
	.B0(\ram[137][5] ), 
	.A1(n6362), 
	.A0(\ram[136][5] ));
   AOI22X1 U9677 (.Y(n11780), 
	.B1(n6381), 
	.B0(\ram[135][5] ), 
	.A1(n6400), 
	.A0(\ram[134][5] ));
   AOI22X1 U9678 (.Y(n11779), 
	.B1(n6419), 
	.B0(\ram[133][5] ), 
	.A1(n6438), 
	.A0(\ram[132][5] ));
   AOI22X1 U9679 (.Y(n11778), 
	.B1(n6457), 
	.B0(\ram[131][5] ), 
	.A1(n6476), 
	.A0(\ram[130][5] ));
   NAND4X1 U9680 (.Y(n11776), 
	.D(n11785), 
	.C(n11784), 
	.B(n11783), 
	.A(n11782));
   AOI22X1 U9681 (.Y(n11785), 
	.B1(n6495), 
	.B0(\ram[129][5] ), 
	.A1(n6514), 
	.A0(\ram[128][5] ));
   AOI22X1 U9682 (.Y(n11784), 
	.B1(n6533), 
	.B0(\ram[143][5] ), 
	.A1(n6553), 
	.A0(\ram[142][5] ));
   AOI22X1 U9683 (.Y(n11783), 
	.B1(n6572), 
	.B0(\ram[141][5] ), 
	.A1(n6591), 
	.A0(\ram[140][5] ));
   AOI22X1 U9684 (.Y(n11782), 
	.B1(n6610), 
	.B0(\ram[139][5] ), 
	.A1(n6629), 
	.A0(\ram[138][5] ));
   OAI21XL U9685 (.Y(n11774), 
	.B0(n9140), 
	.A1(n11787), 
	.A0(n11786));
   NAND4X1 U9686 (.Y(n11787), 
	.D(n11791), 
	.C(n11790), 
	.B(n11789), 
	.A(n11788));
   AOI22X1 U9687 (.Y(n11791), 
	.B1(n6342), 
	.B0(\ram[121][5] ), 
	.A1(n6362), 
	.A0(\ram[120][5] ));
   AOI22X1 U9688 (.Y(n11790), 
	.B1(n6381), 
	.B0(\ram[119][5] ), 
	.A1(n6400), 
	.A0(\ram[118][5] ));
   AOI22X1 U9689 (.Y(n11789), 
	.B1(n6419), 
	.B0(\ram[117][5] ), 
	.A1(n6438), 
	.A0(\ram[116][5] ));
   AOI22X1 U9690 (.Y(n11788), 
	.B1(n6457), 
	.B0(\ram[115][5] ), 
	.A1(n6476), 
	.A0(\ram[114][5] ));
   NAND4X1 U9691 (.Y(n11786), 
	.D(n11795), 
	.C(n11794), 
	.B(n11793), 
	.A(n11792));
   AOI22X1 U9692 (.Y(n11795), 
	.B1(n6495), 
	.B0(\ram[113][5] ), 
	.A1(n6514), 
	.A0(\ram[112][5] ));
   AOI22X1 U9693 (.Y(n11794), 
	.B1(n6533), 
	.B0(\ram[127][5] ), 
	.A1(n6553), 
	.A0(\ram[126][5] ));
   AOI22X1 U9694 (.Y(n11793), 
	.B1(n6572), 
	.B0(\ram[125][5] ), 
	.A1(n6591), 
	.A0(\ram[124][5] ));
   AOI22X1 U9695 (.Y(n11792), 
	.B1(n6610), 
	.B0(\ram[123][5] ), 
	.A1(n6629), 
	.A0(\ram[122][5] ));
   OAI21XL U9696 (.Y(n11773), 
	.B0(n9429), 
	.A1(n11797), 
	.A0(n11796));
   NAND4X1 U9697 (.Y(n11797), 
	.D(n11801), 
	.C(n11800), 
	.B(n11799), 
	.A(n11798));
   AOI22X1 U9698 (.Y(n11801), 
	.B1(n6342), 
	.B0(\ram[105][5] ), 
	.A1(n6362), 
	.A0(\ram[104][5] ));
   AOI22X1 U9699 (.Y(n11800), 
	.B1(n6381), 
	.B0(\ram[103][5] ), 
	.A1(n6400), 
	.A0(\ram[102][5] ));
   AOI22X1 U9700 (.Y(n11799), 
	.B1(n6419), 
	.B0(\ram[101][5] ), 
	.A1(n6438), 
	.A0(\ram[100][5] ));
   AOI22X1 U9701 (.Y(n11798), 
	.B1(n6457), 
	.B0(\ram[99][5] ), 
	.A1(n6476), 
	.A0(\ram[98][5] ));
   NAND4X1 U9702 (.Y(n11796), 
	.D(n11805), 
	.C(n11804), 
	.B(n11803), 
	.A(n11802));
   AOI22X1 U9703 (.Y(n11805), 
	.B1(n6495), 
	.B0(\ram[97][5] ), 
	.A1(n6514), 
	.A0(\ram[96][5] ));
   AOI22X1 U9704 (.Y(n11804), 
	.B1(n6533), 
	.B0(\ram[111][5] ), 
	.A1(n6553), 
	.A0(\ram[110][5] ));
   AOI22X1 U9705 (.Y(n11803), 
	.B1(n6572), 
	.B0(\ram[109][5] ), 
	.A1(n6591), 
	.A0(\ram[108][5] ));
   AOI22X1 U9706 (.Y(n11802), 
	.B1(n6610), 
	.B0(\ram[107][5] ), 
	.A1(n6629), 
	.A0(\ram[106][5] ));
   OAI21XL U9707 (.Y(n11772), 
	.B0(n9718), 
	.A1(n11807), 
	.A0(n11806));
   NAND4X1 U9708 (.Y(n11807), 
	.D(n11811), 
	.C(n11810), 
	.B(n11809), 
	.A(n11808));
   AOI22X1 U9709 (.Y(n11811), 
	.B1(n6342), 
	.B0(\ram[89][5] ), 
	.A1(n6362), 
	.A0(\ram[88][5] ));
   AOI22X1 U9710 (.Y(n11810), 
	.B1(n6381), 
	.B0(\ram[87][5] ), 
	.A1(n6400), 
	.A0(\ram[86][5] ));
   AOI22X1 U9711 (.Y(n11809), 
	.B1(n6419), 
	.B0(\ram[85][5] ), 
	.A1(n6438), 
	.A0(\ram[84][5] ));
   AOI22X1 U9712 (.Y(n11808), 
	.B1(n6457), 
	.B0(\ram[83][5] ), 
	.A1(n6476), 
	.A0(\ram[82][5] ));
   NAND4X1 U9713 (.Y(n11806), 
	.D(n11815), 
	.C(n11814), 
	.B(n11813), 
	.A(n11812));
   AOI22X1 U9714 (.Y(n11815), 
	.B1(n6495), 
	.B0(\ram[81][5] ), 
	.A1(n6514), 
	.A0(\ram[80][5] ));
   AOI22X1 U9715 (.Y(n11814), 
	.B1(n6533), 
	.B0(\ram[95][5] ), 
	.A1(n6553), 
	.A0(\ram[94][5] ));
   AOI22X1 U9716 (.Y(n11813), 
	.B1(n6572), 
	.B0(\ram[93][5] ), 
	.A1(n6591), 
	.A0(\ram[92][5] ));
   AOI22X1 U9717 (.Y(n11812), 
	.B1(n6610), 
	.B0(\ram[91][5] ), 
	.A1(n6629), 
	.A0(\ram[90][5] ));
   NAND4X1 U9718 (.Y(n11680), 
	.D(n11819), 
	.C(n11818), 
	.B(n11817), 
	.A(n11816));
   OAI21XL U9719 (.Y(n11819), 
	.B0(n10007), 
	.A1(n11821), 
	.A0(n11820));
   NAND4X1 U9720 (.Y(n11821), 
	.D(n11825), 
	.C(n11824), 
	.B(n11823), 
	.A(n11822));
   AOI22X1 U9721 (.Y(n11825), 
	.B1(n6342), 
	.B0(\ram[73][5] ), 
	.A1(n6362), 
	.A0(\ram[72][5] ));
   AOI22X1 U9722 (.Y(n11824), 
	.B1(n6381), 
	.B0(\ram[71][5] ), 
	.A1(n6400), 
	.A0(\ram[70][5] ));
   AOI22X1 U9723 (.Y(n11823), 
	.B1(n6419), 
	.B0(\ram[69][5] ), 
	.A1(n6438), 
	.A0(\ram[68][5] ));
   AOI22X1 U9724 (.Y(n11822), 
	.B1(n6457), 
	.B0(\ram[67][5] ), 
	.A1(n6476), 
	.A0(\ram[66][5] ));
   NAND4X1 U9725 (.Y(n11820), 
	.D(n11829), 
	.C(n11828), 
	.B(n11827), 
	.A(n11826));
   AOI22X1 U9726 (.Y(n11829), 
	.B1(n6495), 
	.B0(\ram[65][5] ), 
	.A1(n6514), 
	.A0(\ram[64][5] ));
   AOI22X1 U9727 (.Y(n11828), 
	.B1(n6533), 
	.B0(\ram[79][5] ), 
	.A1(n6553), 
	.A0(\ram[78][5] ));
   AOI22X1 U9728 (.Y(n11827), 
	.B1(n6572), 
	.B0(\ram[77][5] ), 
	.A1(n6591), 
	.A0(\ram[76][5] ));
   AOI22X1 U9729 (.Y(n11826), 
	.B1(n6610), 
	.B0(\ram[75][5] ), 
	.A1(n6629), 
	.A0(\ram[74][5] ));
   OAI21XL U9730 (.Y(n11818), 
	.B0(n10296), 
	.A1(n11831), 
	.A0(n11830));
   NAND4X1 U9731 (.Y(n11831), 
	.D(n11835), 
	.C(n11834), 
	.B(n11833), 
	.A(n11832));
   AOI22X1 U9732 (.Y(n11835), 
	.B1(n6342), 
	.B0(\ram[57][5] ), 
	.A1(n6362), 
	.A0(\ram[56][5] ));
   AOI22X1 U9733 (.Y(n11834), 
	.B1(n6381), 
	.B0(\ram[55][5] ), 
	.A1(n6400), 
	.A0(\ram[54][5] ));
   AOI22X1 U9734 (.Y(n11833), 
	.B1(n6419), 
	.B0(\ram[53][5] ), 
	.A1(n6438), 
	.A0(\ram[52][5] ));
   AOI22X1 U9735 (.Y(n11832), 
	.B1(n6457), 
	.B0(\ram[51][5] ), 
	.A1(n6476), 
	.A0(\ram[50][5] ));
   NAND4X1 U9736 (.Y(n11830), 
	.D(n11839), 
	.C(n11838), 
	.B(n11837), 
	.A(n11836));
   AOI22X1 U9737 (.Y(n11839), 
	.B1(n6495), 
	.B0(\ram[49][5] ), 
	.A1(n6514), 
	.A0(\ram[48][5] ));
   AOI22X1 U9738 (.Y(n11838), 
	.B1(n6533), 
	.B0(\ram[63][5] ), 
	.A1(n6553), 
	.A0(\ram[62][5] ));
   AOI22X1 U9739 (.Y(n11837), 
	.B1(n6572), 
	.B0(\ram[61][5] ), 
	.A1(n6591), 
	.A0(\ram[60][5] ));
   AOI22X1 U9740 (.Y(n11836), 
	.B1(n6610), 
	.B0(\ram[59][5] ), 
	.A1(n6629), 
	.A0(\ram[58][5] ));
   OAI21XL U9741 (.Y(n11817), 
	.B0(n10585), 
	.A1(n11841), 
	.A0(n11840));
   NAND4X1 U9742 (.Y(n11841), 
	.D(n11845), 
	.C(n11844), 
	.B(n11843), 
	.A(n11842));
   AOI22X1 U9743 (.Y(n11845), 
	.B1(n6342), 
	.B0(\ram[41][5] ), 
	.A1(n6362), 
	.A0(\ram[40][5] ));
   AOI22X1 U9744 (.Y(n11844), 
	.B1(n6381), 
	.B0(\ram[39][5] ), 
	.A1(n6400), 
	.A0(\ram[38][5] ));
   AOI22X1 U9745 (.Y(n11843), 
	.B1(n6419), 
	.B0(\ram[37][5] ), 
	.A1(n6438), 
	.A0(\ram[36][5] ));
   AOI22X1 U9746 (.Y(n11842), 
	.B1(n6457), 
	.B0(\ram[35][5] ), 
	.A1(n6476), 
	.A0(\ram[34][5] ));
   NAND4X1 U9747 (.Y(n11840), 
	.D(n11849), 
	.C(n11848), 
	.B(n11847), 
	.A(n11846));
   AOI22X1 U9748 (.Y(n11849), 
	.B1(n6495), 
	.B0(\ram[33][5] ), 
	.A1(n6514), 
	.A0(\ram[32][5] ));
   AOI22X1 U9749 (.Y(n11848), 
	.B1(n6533), 
	.B0(\ram[47][5] ), 
	.A1(n6553), 
	.A0(\ram[46][5] ));
   AOI22X1 U9750 (.Y(n11847), 
	.B1(n6572), 
	.B0(\ram[45][5] ), 
	.A1(n6591), 
	.A0(\ram[44][5] ));
   AOI22X1 U9751 (.Y(n11846), 
	.B1(n6610), 
	.B0(\ram[43][5] ), 
	.A1(n6629), 
	.A0(\ram[42][5] ));
   OAI21XL U9752 (.Y(n11816), 
	.B0(n6343), 
	.A1(n11851), 
	.A0(n11850));
   NAND4X1 U9753 (.Y(n11851), 
	.D(n11855), 
	.C(n11854), 
	.B(n11853), 
	.A(n11852));
   AOI22X1 U9754 (.Y(n11855), 
	.B1(n6342), 
	.B0(\ram[25][5] ), 
	.A1(n6362), 
	.A0(\ram[24][5] ));
   AOI22X1 U9755 (.Y(n11854), 
	.B1(n6381), 
	.B0(\ram[23][5] ), 
	.A1(n6400), 
	.A0(\ram[22][5] ));
   AOI22X1 U9756 (.Y(n11853), 
	.B1(n6419), 
	.B0(\ram[21][5] ), 
	.A1(n6438), 
	.A0(\ram[20][5] ));
   AOI22X1 U9757 (.Y(n11852), 
	.B1(n6457), 
	.B0(\ram[19][5] ), 
	.A1(n6476), 
	.A0(\ram[18][5] ));
   NAND4X1 U9758 (.Y(n11850), 
	.D(n11859), 
	.C(n11858), 
	.B(n11857), 
	.A(n11856));
   AOI22X1 U9759 (.Y(n11859), 
	.B1(n6495), 
	.B0(\ram[17][5] ), 
	.A1(n6514), 
	.A0(\ram[16][5] ));
   AOI22X1 U9760 (.Y(n11858), 
	.B1(n6533), 
	.B0(\ram[31][5] ), 
	.A1(n6553), 
	.A0(\ram[30][5] ));
   AOI22X1 U9761 (.Y(n11857), 
	.B1(n6572), 
	.B0(\ram[29][5] ), 
	.A1(n6591), 
	.A0(\ram[28][5] ));
   AOI22X1 U9762 (.Y(n11856), 
	.B1(n6610), 
	.B0(\ram[27][5] ), 
	.A1(n6629), 
	.A0(\ram[26][5] ));
   OR4X1 U9763 (.Y(mem_read_data[4]), 
	.D(n11863), 
	.C(n11862), 
	.B(n11861), 
	.A(n11860));
   NAND4X1 U9764 (.Y(n11863), 
	.D(n11867), 
	.C(n11866), 
	.B(n11865), 
	.A(n11864));
   OAI21XL U9765 (.Y(n11867), 
	.B0(n6534), 
	.A1(n11869), 
	.A0(n11868));
   NAND4X1 U9766 (.Y(n11869), 
	.D(n11873), 
	.C(n11872), 
	.B(n11871), 
	.A(n11870));
   AOI22X1 U9767 (.Y(n11873), 
	.B1(n6342), 
	.B0(\ram[9][4] ), 
	.A1(n6362), 
	.A0(\ram[8][4] ));
   AOI22X1 U9768 (.Y(n11872), 
	.B1(n6381), 
	.B0(\ram[7][4] ), 
	.A1(n6400), 
	.A0(\ram[6][4] ));
   AOI22X1 U9769 (.Y(n11871), 
	.B1(n6419), 
	.B0(\ram[5][4] ), 
	.A1(n6438), 
	.A0(\ram[4][4] ));
   AOI22X1 U9770 (.Y(n11870), 
	.B1(n6457), 
	.B0(\ram[3][4] ), 
	.A1(n6476), 
	.A0(\ram[2][4] ));
   NAND4X1 U9771 (.Y(n11868), 
	.D(n11877), 
	.C(n11876), 
	.B(n11875), 
	.A(n11874));
   AOI22X1 U9772 (.Y(n11877), 
	.B1(n6495), 
	.B0(\ram[1][4] ), 
	.A1(n6514), 
	.A0(\ram[0][4] ));
   AOI22X1 U9773 (.Y(n11876), 
	.B1(n6533), 
	.B0(\ram[15][4] ), 
	.A1(n6553), 
	.A0(\ram[14][4] ));
   AOI22X1 U9774 (.Y(n11875), 
	.B1(n6572), 
	.B0(\ram[13][4] ), 
	.A1(n6591), 
	.A0(\ram[12][4] ));
   AOI22X1 U9775 (.Y(n11874), 
	.B1(n6610), 
	.B0(\ram[11][4] ), 
	.A1(n6629), 
	.A0(\ram[10][4] ));
   OAI21XL U9776 (.Y(n11866), 
	.B0(n6828), 
	.A1(n11879), 
	.A0(n11878));
   NAND4X1 U9777 (.Y(n11879), 
	.D(n11883), 
	.C(n11882), 
	.B(n11881), 
	.A(n11880));
   AOI22X1 U9778 (.Y(n11883), 
	.B1(n6342), 
	.B0(\ram[249][4] ), 
	.A1(n6362), 
	.A0(\ram[248][4] ));
   AOI22X1 U9779 (.Y(n11882), 
	.B1(n6381), 
	.B0(\ram[247][4] ), 
	.A1(n6400), 
	.A0(\ram[246][4] ));
   AOI22X1 U9780 (.Y(n11881), 
	.B1(n6419), 
	.B0(\ram[245][4] ), 
	.A1(n6438), 
	.A0(\ram[244][4] ));
   AOI22X1 U9781 (.Y(n11880), 
	.B1(n6457), 
	.B0(\ram[243][4] ), 
	.A1(n6476), 
	.A0(\ram[242][4] ));
   NAND4X1 U9782 (.Y(n11878), 
	.D(n11887), 
	.C(n11886), 
	.B(n11885), 
	.A(n11884));
   AOI22X1 U9783 (.Y(n11887), 
	.B1(n6495), 
	.B0(\ram[241][4] ), 
	.A1(n6514), 
	.A0(\ram[240][4] ));
   AOI22X1 U9784 (.Y(n11886), 
	.B1(n6533), 
	.B0(\ram[255][4] ), 
	.A1(n6553), 
	.A0(\ram[254][4] ));
   AOI22X1 U9785 (.Y(n11885), 
	.B1(n6572), 
	.B0(\ram[253][4] ), 
	.A1(n6591), 
	.A0(\ram[252][4] ));
   AOI22X1 U9786 (.Y(n11884), 
	.B1(n6610), 
	.B0(\ram[251][4] ), 
	.A1(n6629), 
	.A0(\ram[250][4] ));
   OAI21XL U9787 (.Y(n11865), 
	.B0(n7117), 
	.A1(n11889), 
	.A0(n11888));
   NAND4X1 U9788 (.Y(n11889), 
	.D(n11893), 
	.C(n11892), 
	.B(n11891), 
	.A(n11890));
   AOI22X1 U9789 (.Y(n11893), 
	.B1(n6342), 
	.B0(\ram[233][4] ), 
	.A1(n6362), 
	.A0(\ram[232][4] ));
   AOI22X1 U9790 (.Y(n11892), 
	.B1(n6381), 
	.B0(\ram[231][4] ), 
	.A1(n6400), 
	.A0(\ram[230][4] ));
   AOI22X1 U9791 (.Y(n11891), 
	.B1(n6419), 
	.B0(\ram[229][4] ), 
	.A1(n6438), 
	.A0(\ram[228][4] ));
   AOI22X1 U9792 (.Y(n11890), 
	.B1(n6457), 
	.B0(\ram[227][4] ), 
	.A1(n6476), 
	.A0(\ram[226][4] ));
   NAND4X1 U9793 (.Y(n11888), 
	.D(n11897), 
	.C(n11896), 
	.B(n11895), 
	.A(n11894));
   AOI22X1 U9794 (.Y(n11897), 
	.B1(n6495), 
	.B0(\ram[225][4] ), 
	.A1(n6514), 
	.A0(\ram[224][4] ));
   AOI22X1 U9795 (.Y(n11896), 
	.B1(n6533), 
	.B0(\ram[239][4] ), 
	.A1(n6553), 
	.A0(\ram[238][4] ));
   AOI22X1 U9796 (.Y(n11895), 
	.B1(n6572), 
	.B0(\ram[237][4] ), 
	.A1(n6591), 
	.A0(\ram[236][4] ));
   AOI22X1 U9797 (.Y(n11894), 
	.B1(n6610), 
	.B0(\ram[235][4] ), 
	.A1(n6629), 
	.A0(\ram[234][4] ));
   OAI21XL U9798 (.Y(n11864), 
	.B0(n7406), 
	.A1(n11899), 
	.A0(n11898));
   NAND4X1 U9799 (.Y(n11899), 
	.D(n11903), 
	.C(n11902), 
	.B(n11901), 
	.A(n11900));
   AOI22X1 U9800 (.Y(n11903), 
	.B1(n6342), 
	.B0(\ram[217][4] ), 
	.A1(n6362), 
	.A0(\ram[216][4] ));
   AOI22X1 U9801 (.Y(n11902), 
	.B1(n6381), 
	.B0(\ram[215][4] ), 
	.A1(n6400), 
	.A0(\ram[214][4] ));
   AOI22X1 U9802 (.Y(n11901), 
	.B1(n6419), 
	.B0(\ram[213][4] ), 
	.A1(n6438), 
	.A0(\ram[212][4] ));
   AOI22X1 U9803 (.Y(n11900), 
	.B1(n6457), 
	.B0(\ram[211][4] ), 
	.A1(n6476), 
	.A0(\ram[210][4] ));
   NAND4X1 U9804 (.Y(n11898), 
	.D(n11907), 
	.C(n11906), 
	.B(n11905), 
	.A(n11904));
   AOI22X1 U9805 (.Y(n11907), 
	.B1(n6495), 
	.B0(\ram[209][4] ), 
	.A1(n6514), 
	.A0(\ram[208][4] ));
   AOI22X1 U9806 (.Y(n11906), 
	.B1(n6533), 
	.B0(\ram[223][4] ), 
	.A1(n6553), 
	.A0(\ram[222][4] ));
   AOI22X1 U9807 (.Y(n11905), 
	.B1(n6572), 
	.B0(\ram[221][4] ), 
	.A1(n6591), 
	.A0(\ram[220][4] ));
   AOI22X1 U9808 (.Y(n11904), 
	.B1(n6610), 
	.B0(\ram[219][4] ), 
	.A1(n6629), 
	.A0(\ram[218][4] ));
   NAND4X1 U9809 (.Y(n11862), 
	.D(n11911), 
	.C(n11910), 
	.B(n11909), 
	.A(n11908));
   OAI21XL U9810 (.Y(n11911), 
	.B0(n7695), 
	.A1(n11913), 
	.A0(n11912));
   NAND4X1 U9811 (.Y(n11913), 
	.D(n11917), 
	.C(n11916), 
	.B(n11915), 
	.A(n11914));
   AOI22X1 U9812 (.Y(n11917), 
	.B1(n6342), 
	.B0(\ram[201][4] ), 
	.A1(n6362), 
	.A0(\ram[200][4] ));
   AOI22X1 U9813 (.Y(n11916), 
	.B1(n6381), 
	.B0(\ram[199][4] ), 
	.A1(n6400), 
	.A0(\ram[198][4] ));
   AOI22X1 U9814 (.Y(n11915), 
	.B1(n6419), 
	.B0(\ram[197][4] ), 
	.A1(n6438), 
	.A0(\ram[196][4] ));
   AOI22X1 U9815 (.Y(n11914), 
	.B1(n6457), 
	.B0(\ram[195][4] ), 
	.A1(n6476), 
	.A0(\ram[194][4] ));
   NAND4X1 U9816 (.Y(n11912), 
	.D(n11921), 
	.C(n11920), 
	.B(n11919), 
	.A(n11918));
   AOI22X1 U9817 (.Y(n11921), 
	.B1(n6495), 
	.B0(\ram[193][4] ), 
	.A1(n6514), 
	.A0(\ram[192][4] ));
   AOI22X1 U9818 (.Y(n11920), 
	.B1(n6533), 
	.B0(\ram[207][4] ), 
	.A1(n6553), 
	.A0(\ram[206][4] ));
   AOI22X1 U9819 (.Y(n11919), 
	.B1(n6572), 
	.B0(\ram[205][4] ), 
	.A1(n6591), 
	.A0(\ram[204][4] ));
   AOI22X1 U9820 (.Y(n11918), 
	.B1(n6610), 
	.B0(\ram[203][4] ), 
	.A1(n6629), 
	.A0(\ram[202][4] ));
   OAI21XL U9821 (.Y(n11910), 
	.B0(n7984), 
	.A1(n11923), 
	.A0(n11922));
   NAND4X1 U9822 (.Y(n11923), 
	.D(n11927), 
	.C(n11926), 
	.B(n11925), 
	.A(n11924));
   AOI22X1 U9823 (.Y(n11927), 
	.B1(n6342), 
	.B0(\ram[185][4] ), 
	.A1(n6362), 
	.A0(\ram[184][4] ));
   AOI22X1 U9824 (.Y(n11926), 
	.B1(n6381), 
	.B0(\ram[183][4] ), 
	.A1(n6400), 
	.A0(\ram[182][4] ));
   AOI22X1 U9825 (.Y(n11925), 
	.B1(n6419), 
	.B0(\ram[181][4] ), 
	.A1(n6438), 
	.A0(\ram[180][4] ));
   AOI22X1 U9826 (.Y(n11924), 
	.B1(n6457), 
	.B0(\ram[179][4] ), 
	.A1(n6476), 
	.A0(\ram[178][4] ));
   NAND4X1 U9827 (.Y(n11922), 
	.D(n11931), 
	.C(n11930), 
	.B(n11929), 
	.A(n11928));
   AOI22X1 U9828 (.Y(n11931), 
	.B1(n6495), 
	.B0(\ram[177][4] ), 
	.A1(n6514), 
	.A0(\ram[176][4] ));
   AOI22X1 U9829 (.Y(n11930), 
	.B1(n6533), 
	.B0(\ram[191][4] ), 
	.A1(n6553), 
	.A0(\ram[190][4] ));
   AOI22X1 U9830 (.Y(n11929), 
	.B1(n6572), 
	.B0(\ram[189][4] ), 
	.A1(n6591), 
	.A0(\ram[188][4] ));
   AOI22X1 U9831 (.Y(n11928), 
	.B1(n6610), 
	.B0(\ram[187][4] ), 
	.A1(n6629), 
	.A0(\ram[186][4] ));
   OAI21XL U9832 (.Y(n11909), 
	.B0(n8273), 
	.A1(n11933), 
	.A0(n11932));
   NAND4X1 U9833 (.Y(n11933), 
	.D(n11937), 
	.C(n11936), 
	.B(n11935), 
	.A(n11934));
   AOI22X1 U9834 (.Y(n11937), 
	.B1(n6342), 
	.B0(\ram[169][4] ), 
	.A1(n6362), 
	.A0(\ram[168][4] ));
   AOI22X1 U9835 (.Y(n11936), 
	.B1(n6381), 
	.B0(\ram[167][4] ), 
	.A1(n6400), 
	.A0(\ram[166][4] ));
   AOI22X1 U9836 (.Y(n11935), 
	.B1(n6419), 
	.B0(\ram[165][4] ), 
	.A1(n6438), 
	.A0(\ram[164][4] ));
   AOI22X1 U9837 (.Y(n11934), 
	.B1(n6457), 
	.B0(\ram[163][4] ), 
	.A1(n6476), 
	.A0(\ram[162][4] ));
   NAND4X1 U9838 (.Y(n11932), 
	.D(n11941), 
	.C(n11940), 
	.B(n11939), 
	.A(n11938));
   AOI22X1 U9839 (.Y(n11941), 
	.B1(n6495), 
	.B0(\ram[161][4] ), 
	.A1(n6514), 
	.A0(\ram[160][4] ));
   AOI22X1 U9840 (.Y(n11940), 
	.B1(n6533), 
	.B0(\ram[175][4] ), 
	.A1(n6553), 
	.A0(\ram[174][4] ));
   AOI22X1 U9841 (.Y(n11939), 
	.B1(n6572), 
	.B0(\ram[173][4] ), 
	.A1(n6591), 
	.A0(\ram[172][4] ));
   AOI22X1 U9842 (.Y(n11938), 
	.B1(n6610), 
	.B0(\ram[171][4] ), 
	.A1(n6629), 
	.A0(\ram[170][4] ));
   OAI21XL U9843 (.Y(n11908), 
	.B0(n8562), 
	.A1(n11943), 
	.A0(n11942));
   NAND4X1 U9844 (.Y(n11943), 
	.D(n11947), 
	.C(n11946), 
	.B(n11945), 
	.A(n11944));
   AOI22X1 U9845 (.Y(n11947), 
	.B1(n6342), 
	.B0(\ram[153][4] ), 
	.A1(n6362), 
	.A0(\ram[152][4] ));
   AOI22X1 U9846 (.Y(n11946), 
	.B1(n6381), 
	.B0(\ram[151][4] ), 
	.A1(n6400), 
	.A0(\ram[150][4] ));
   AOI22X1 U9847 (.Y(n11945), 
	.B1(n6419), 
	.B0(\ram[149][4] ), 
	.A1(n6438), 
	.A0(\ram[148][4] ));
   AOI22X1 U9848 (.Y(n11944), 
	.B1(n6457), 
	.B0(\ram[147][4] ), 
	.A1(n6476), 
	.A0(\ram[146][4] ));
   NAND4X1 U9849 (.Y(n11942), 
	.D(n11951), 
	.C(n11950), 
	.B(n11949), 
	.A(n11948));
   AOI22X1 U9850 (.Y(n11951), 
	.B1(n6495), 
	.B0(\ram[145][4] ), 
	.A1(n6514), 
	.A0(\ram[144][4] ));
   AOI22X1 U9851 (.Y(n11950), 
	.B1(n6533), 
	.B0(\ram[159][4] ), 
	.A1(n6553), 
	.A0(\ram[158][4] ));
   AOI22X1 U9852 (.Y(n11949), 
	.B1(n6572), 
	.B0(\ram[157][4] ), 
	.A1(n6591), 
	.A0(\ram[156][4] ));
   AOI22X1 U9853 (.Y(n11948), 
	.B1(n6610), 
	.B0(\ram[155][4] ), 
	.A1(n6629), 
	.A0(\ram[154][4] ));
   NAND4X1 U9854 (.Y(n11861), 
	.D(n11955), 
	.C(n11954), 
	.B(n11953), 
	.A(n11952));
   OAI21XL U9855 (.Y(n11955), 
	.B0(n8851), 
	.A1(n11957), 
	.A0(n11956));
   NAND4X1 U9856 (.Y(n11957), 
	.D(n11961), 
	.C(n11960), 
	.B(n11959), 
	.A(n11958));
   AOI22X1 U9857 (.Y(n11961), 
	.B1(n6342), 
	.B0(\ram[137][4] ), 
	.A1(n6362), 
	.A0(\ram[136][4] ));
   AOI22X1 U9858 (.Y(n11960), 
	.B1(n6381), 
	.B0(\ram[135][4] ), 
	.A1(n6400), 
	.A0(\ram[134][4] ));
   AOI22X1 U9859 (.Y(n11959), 
	.B1(n6419), 
	.B0(\ram[133][4] ), 
	.A1(n6438), 
	.A0(\ram[132][4] ));
   AOI22X1 U9860 (.Y(n11958), 
	.B1(n6457), 
	.B0(\ram[131][4] ), 
	.A1(n6476), 
	.A0(\ram[130][4] ));
   NAND4X1 U9861 (.Y(n11956), 
	.D(n11965), 
	.C(n11964), 
	.B(n11963), 
	.A(n11962));
   AOI22X1 U9862 (.Y(n11965), 
	.B1(n6495), 
	.B0(\ram[129][4] ), 
	.A1(n6514), 
	.A0(\ram[128][4] ));
   AOI22X1 U9863 (.Y(n11964), 
	.B1(n6533), 
	.B0(\ram[143][4] ), 
	.A1(n6553), 
	.A0(\ram[142][4] ));
   AOI22X1 U9864 (.Y(n11963), 
	.B1(n6572), 
	.B0(\ram[141][4] ), 
	.A1(n6591), 
	.A0(\ram[140][4] ));
   AOI22X1 U9865 (.Y(n11962), 
	.B1(n6610), 
	.B0(\ram[139][4] ), 
	.A1(n6629), 
	.A0(\ram[138][4] ));
   OAI21XL U9866 (.Y(n11954), 
	.B0(n9140), 
	.A1(n11967), 
	.A0(n11966));
   NAND4X1 U9867 (.Y(n11967), 
	.D(n11971), 
	.C(n11970), 
	.B(n11969), 
	.A(n11968));
   AOI22X1 U9868 (.Y(n11971), 
	.B1(n6342), 
	.B0(\ram[121][4] ), 
	.A1(n6362), 
	.A0(\ram[120][4] ));
   AOI22X1 U9869 (.Y(n11970), 
	.B1(n6381), 
	.B0(\ram[119][4] ), 
	.A1(n6400), 
	.A0(\ram[118][4] ));
   AOI22X1 U9870 (.Y(n11969), 
	.B1(n6419), 
	.B0(\ram[117][4] ), 
	.A1(n6438), 
	.A0(\ram[116][4] ));
   AOI22X1 U9871 (.Y(n11968), 
	.B1(n6457), 
	.B0(\ram[115][4] ), 
	.A1(n6476), 
	.A0(\ram[114][4] ));
   NAND4X1 U9872 (.Y(n11966), 
	.D(n11975), 
	.C(n11974), 
	.B(n11973), 
	.A(n11972));
   AOI22X1 U9873 (.Y(n11975), 
	.B1(n6495), 
	.B0(\ram[113][4] ), 
	.A1(n6514), 
	.A0(\ram[112][4] ));
   AOI22X1 U9874 (.Y(n11974), 
	.B1(n6533), 
	.B0(\ram[127][4] ), 
	.A1(n6553), 
	.A0(\ram[126][4] ));
   AOI22X1 U9875 (.Y(n11973), 
	.B1(n6572), 
	.B0(\ram[125][4] ), 
	.A1(n6591), 
	.A0(\ram[124][4] ));
   AOI22X1 U9876 (.Y(n11972), 
	.B1(n6610), 
	.B0(\ram[123][4] ), 
	.A1(n6629), 
	.A0(\ram[122][4] ));
   OAI21XL U9877 (.Y(n11953), 
	.B0(n9429), 
	.A1(n11977), 
	.A0(n11976));
   NAND4X1 U9878 (.Y(n11977), 
	.D(n11981), 
	.C(n11980), 
	.B(n11979), 
	.A(n11978));
   AOI22X1 U9879 (.Y(n11981), 
	.B1(n6342), 
	.B0(\ram[105][4] ), 
	.A1(n6362), 
	.A0(\ram[104][4] ));
   AOI22X1 U9880 (.Y(n11980), 
	.B1(n6381), 
	.B0(\ram[103][4] ), 
	.A1(n6400), 
	.A0(\ram[102][4] ));
   AOI22X1 U9881 (.Y(n11979), 
	.B1(n6419), 
	.B0(\ram[101][4] ), 
	.A1(n6438), 
	.A0(\ram[100][4] ));
   AOI22X1 U9882 (.Y(n11978), 
	.B1(n6457), 
	.B0(\ram[99][4] ), 
	.A1(n6476), 
	.A0(\ram[98][4] ));
   NAND4X1 U9883 (.Y(n11976), 
	.D(n11985), 
	.C(n11984), 
	.B(n11983), 
	.A(n11982));
   AOI22X1 U9884 (.Y(n11985), 
	.B1(n6495), 
	.B0(\ram[97][4] ), 
	.A1(n6514), 
	.A0(\ram[96][4] ));
   AOI22X1 U9885 (.Y(n11984), 
	.B1(n6533), 
	.B0(\ram[111][4] ), 
	.A1(n6553), 
	.A0(\ram[110][4] ));
   AOI22X1 U9886 (.Y(n11983), 
	.B1(n6572), 
	.B0(\ram[109][4] ), 
	.A1(n6591), 
	.A0(\ram[108][4] ));
   AOI22X1 U9887 (.Y(n11982), 
	.B1(n6610), 
	.B0(\ram[107][4] ), 
	.A1(n6629), 
	.A0(\ram[106][4] ));
   OAI21XL U9888 (.Y(n11952), 
	.B0(n9718), 
	.A1(n11987), 
	.A0(n11986));
   NAND4X1 U9889 (.Y(n11987), 
	.D(n11991), 
	.C(n11990), 
	.B(n11989), 
	.A(n11988));
   AOI22X1 U9890 (.Y(n11991), 
	.B1(n6342), 
	.B0(\ram[89][4] ), 
	.A1(n6362), 
	.A0(\ram[88][4] ));
   AOI22X1 U9891 (.Y(n11990), 
	.B1(n6381), 
	.B0(\ram[87][4] ), 
	.A1(n6400), 
	.A0(\ram[86][4] ));
   AOI22X1 U9892 (.Y(n11989), 
	.B1(n6419), 
	.B0(\ram[85][4] ), 
	.A1(n6438), 
	.A0(\ram[84][4] ));
   AOI22X1 U9893 (.Y(n11988), 
	.B1(n6457), 
	.B0(\ram[83][4] ), 
	.A1(n6476), 
	.A0(\ram[82][4] ));
   NAND4X1 U9894 (.Y(n11986), 
	.D(n11995), 
	.C(n11994), 
	.B(n11993), 
	.A(n11992));
   AOI22X1 U9895 (.Y(n11995), 
	.B1(n6495), 
	.B0(\ram[81][4] ), 
	.A1(n6514), 
	.A0(\ram[80][4] ));
   AOI22X1 U9896 (.Y(n11994), 
	.B1(n6533), 
	.B0(\ram[95][4] ), 
	.A1(n6553), 
	.A0(\ram[94][4] ));
   AOI22X1 U9897 (.Y(n11993), 
	.B1(n6572), 
	.B0(\ram[93][4] ), 
	.A1(n6591), 
	.A0(\ram[92][4] ));
   AOI22X1 U9898 (.Y(n11992), 
	.B1(n6610), 
	.B0(\ram[91][4] ), 
	.A1(n6629), 
	.A0(\ram[90][4] ));
   NAND4X1 U9899 (.Y(n11860), 
	.D(n11999), 
	.C(n11998), 
	.B(n11997), 
	.A(n11996));
   OAI21XL U9900 (.Y(n11999), 
	.B0(n10007), 
	.A1(n12001), 
	.A0(n12000));
   NAND4X1 U9901 (.Y(n12001), 
	.D(n12005), 
	.C(n12004), 
	.B(n12003), 
	.A(n12002));
   AOI22X1 U9902 (.Y(n12005), 
	.B1(n6342), 
	.B0(\ram[73][4] ), 
	.A1(n6362), 
	.A0(\ram[72][4] ));
   AOI22X1 U9903 (.Y(n12004), 
	.B1(n6381), 
	.B0(\ram[71][4] ), 
	.A1(n6400), 
	.A0(\ram[70][4] ));
   AOI22X1 U9904 (.Y(n12003), 
	.B1(n6419), 
	.B0(\ram[69][4] ), 
	.A1(n6438), 
	.A0(\ram[68][4] ));
   AOI22X1 U9905 (.Y(n12002), 
	.B1(n6457), 
	.B0(\ram[67][4] ), 
	.A1(n6476), 
	.A0(\ram[66][4] ));
   NAND4X1 U9906 (.Y(n12000), 
	.D(n12009), 
	.C(n12008), 
	.B(n12007), 
	.A(n12006));
   AOI22X1 U9907 (.Y(n12009), 
	.B1(n6495), 
	.B0(\ram[65][4] ), 
	.A1(n6514), 
	.A0(\ram[64][4] ));
   AOI22X1 U9908 (.Y(n12008), 
	.B1(n6533), 
	.B0(\ram[79][4] ), 
	.A1(n6553), 
	.A0(\ram[78][4] ));
   AOI22X1 U9909 (.Y(n12007), 
	.B1(n6572), 
	.B0(\ram[77][4] ), 
	.A1(n6591), 
	.A0(\ram[76][4] ));
   AOI22X1 U9910 (.Y(n12006), 
	.B1(n6610), 
	.B0(\ram[75][4] ), 
	.A1(n6629), 
	.A0(\ram[74][4] ));
   OAI21XL U9911 (.Y(n11998), 
	.B0(n10296), 
	.A1(n12011), 
	.A0(n12010));
   NAND4X1 U9912 (.Y(n12011), 
	.D(n12015), 
	.C(n12014), 
	.B(n12013), 
	.A(n12012));
   AOI22X1 U9913 (.Y(n12015), 
	.B1(n6342), 
	.B0(\ram[57][4] ), 
	.A1(n6362), 
	.A0(\ram[56][4] ));
   AOI22X1 U9914 (.Y(n12014), 
	.B1(n6381), 
	.B0(\ram[55][4] ), 
	.A1(n6400), 
	.A0(\ram[54][4] ));
   AOI22X1 U9915 (.Y(n12013), 
	.B1(n6419), 
	.B0(\ram[53][4] ), 
	.A1(n6438), 
	.A0(\ram[52][4] ));
   AOI22X1 U9916 (.Y(n12012), 
	.B1(n6457), 
	.B0(\ram[51][4] ), 
	.A1(n6476), 
	.A0(\ram[50][4] ));
   NAND4X1 U9917 (.Y(n12010), 
	.D(n12019), 
	.C(n12018), 
	.B(n12017), 
	.A(n12016));
   AOI22X1 U9918 (.Y(n12019), 
	.B1(n6495), 
	.B0(\ram[49][4] ), 
	.A1(n6514), 
	.A0(\ram[48][4] ));
   AOI22X1 U9919 (.Y(n12018), 
	.B1(n6533), 
	.B0(\ram[63][4] ), 
	.A1(n6553), 
	.A0(\ram[62][4] ));
   AOI22X1 U9920 (.Y(n12017), 
	.B1(n6572), 
	.B0(\ram[61][4] ), 
	.A1(n6591), 
	.A0(\ram[60][4] ));
   AOI22X1 U9921 (.Y(n12016), 
	.B1(n6610), 
	.B0(\ram[59][4] ), 
	.A1(n6629), 
	.A0(\ram[58][4] ));
   OAI21XL U9922 (.Y(n11997), 
	.B0(n10585), 
	.A1(n12021), 
	.A0(n12020));
   NAND4X1 U9923 (.Y(n12021), 
	.D(n12025), 
	.C(n12024), 
	.B(n12023), 
	.A(n12022));
   AOI22X1 U9924 (.Y(n12025), 
	.B1(n6342), 
	.B0(\ram[41][4] ), 
	.A1(n6362), 
	.A0(\ram[40][4] ));
   AOI22X1 U9925 (.Y(n12024), 
	.B1(n6381), 
	.B0(\ram[39][4] ), 
	.A1(n6400), 
	.A0(\ram[38][4] ));
   AOI22X1 U9926 (.Y(n12023), 
	.B1(n6419), 
	.B0(\ram[37][4] ), 
	.A1(n6438), 
	.A0(\ram[36][4] ));
   AOI22X1 U9927 (.Y(n12022), 
	.B1(n6457), 
	.B0(\ram[35][4] ), 
	.A1(n6476), 
	.A0(\ram[34][4] ));
   NAND4X1 U9928 (.Y(n12020), 
	.D(n12029), 
	.C(n12028), 
	.B(n12027), 
	.A(n12026));
   AOI22X1 U9929 (.Y(n12029), 
	.B1(n6495), 
	.B0(\ram[33][4] ), 
	.A1(n6514), 
	.A0(\ram[32][4] ));
   AOI22X1 U9930 (.Y(n12028), 
	.B1(n6533), 
	.B0(\ram[47][4] ), 
	.A1(n6553), 
	.A0(\ram[46][4] ));
   AOI22X1 U9931 (.Y(n12027), 
	.B1(n6572), 
	.B0(\ram[45][4] ), 
	.A1(n6591), 
	.A0(\ram[44][4] ));
   AOI22X1 U9932 (.Y(n12026), 
	.B1(n6610), 
	.B0(\ram[43][4] ), 
	.A1(n6629), 
	.A0(\ram[42][4] ));
   OAI21XL U9933 (.Y(n11996), 
	.B0(n6343), 
	.A1(n12031), 
	.A0(n12030));
   NAND4X1 U9934 (.Y(n12031), 
	.D(n12035), 
	.C(n12034), 
	.B(n12033), 
	.A(n12032));
   AOI22X1 U9935 (.Y(n12035), 
	.B1(n6342), 
	.B0(\ram[25][4] ), 
	.A1(n6362), 
	.A0(\ram[24][4] ));
   AOI22X1 U9936 (.Y(n12034), 
	.B1(n6381), 
	.B0(\ram[23][4] ), 
	.A1(n6400), 
	.A0(\ram[22][4] ));
   AOI22X1 U9937 (.Y(n12033), 
	.B1(n6419), 
	.B0(\ram[21][4] ), 
	.A1(n6438), 
	.A0(\ram[20][4] ));
   AOI22X1 U9938 (.Y(n12032), 
	.B1(n6457), 
	.B0(\ram[19][4] ), 
	.A1(n6476), 
	.A0(\ram[18][4] ));
   NAND4X1 U9939 (.Y(n12030), 
	.D(n12039), 
	.C(n12038), 
	.B(n12037), 
	.A(n12036));
   AOI22X1 U9940 (.Y(n12039), 
	.B1(n6495), 
	.B0(\ram[17][4] ), 
	.A1(n6514), 
	.A0(\ram[16][4] ));
   AOI22X1 U9941 (.Y(n12038), 
	.B1(n6533), 
	.B0(\ram[31][4] ), 
	.A1(n6553), 
	.A0(\ram[30][4] ));
   AOI22X1 U9942 (.Y(n12037), 
	.B1(n6572), 
	.B0(\ram[29][4] ), 
	.A1(n6591), 
	.A0(\ram[28][4] ));
   AOI22X1 U9943 (.Y(n12036), 
	.B1(n6610), 
	.B0(\ram[27][4] ), 
	.A1(n6629), 
	.A0(\ram[26][4] ));
   OR4X1 U9944 (.Y(mem_read_data[3]), 
	.D(n12043), 
	.C(n12042), 
	.B(n12041), 
	.A(n12040));
   NAND4X1 U9945 (.Y(n12043), 
	.D(n12047), 
	.C(n12046), 
	.B(n12045), 
	.A(n12044));
   OAI21XL U9946 (.Y(n12047), 
	.B0(n6534), 
	.A1(n12049), 
	.A0(n12048));
   NAND4X1 U9947 (.Y(n12049), 
	.D(n12053), 
	.C(n12052), 
	.B(n12051), 
	.A(n12050));
   AOI22X1 U9948 (.Y(n12053), 
	.B1(n6342), 
	.B0(\ram[9][3] ), 
	.A1(n6362), 
	.A0(\ram[8][3] ));
   AOI22X1 U9949 (.Y(n12052), 
	.B1(n6381), 
	.B0(\ram[7][3] ), 
	.A1(n6400), 
	.A0(\ram[6][3] ));
   AOI22X1 U9950 (.Y(n12051), 
	.B1(n6419), 
	.B0(\ram[5][3] ), 
	.A1(n6438), 
	.A0(\ram[4][3] ));
   AOI22X1 U9951 (.Y(n12050), 
	.B1(n6457), 
	.B0(\ram[3][3] ), 
	.A1(n6476), 
	.A0(\ram[2][3] ));
   NAND4X1 U9952 (.Y(n12048), 
	.D(n12057), 
	.C(n12056), 
	.B(n12055), 
	.A(n12054));
   AOI22X1 U9953 (.Y(n12057), 
	.B1(n6495), 
	.B0(\ram[1][3] ), 
	.A1(n6514), 
	.A0(\ram[0][3] ));
   AOI22X1 U9954 (.Y(n12056), 
	.B1(n6533), 
	.B0(\ram[15][3] ), 
	.A1(n6553), 
	.A0(\ram[14][3] ));
   AOI22X1 U9955 (.Y(n12055), 
	.B1(n6572), 
	.B0(\ram[13][3] ), 
	.A1(n6591), 
	.A0(\ram[12][3] ));
   AOI22X1 U9956 (.Y(n12054), 
	.B1(n6610), 
	.B0(\ram[11][3] ), 
	.A1(n6629), 
	.A0(\ram[10][3] ));
   OAI21XL U9957 (.Y(n12046), 
	.B0(n6828), 
	.A1(n12059), 
	.A0(n12058));
   NAND4X1 U9958 (.Y(n12059), 
	.D(n12063), 
	.C(n12062), 
	.B(n12061), 
	.A(n12060));
   AOI22X1 U9959 (.Y(n12063), 
	.B1(n6342), 
	.B0(\ram[249][3] ), 
	.A1(n6362), 
	.A0(\ram[248][3] ));
   AOI22X1 U9960 (.Y(n12062), 
	.B1(n6381), 
	.B0(\ram[247][3] ), 
	.A1(n6400), 
	.A0(\ram[246][3] ));
   AOI22X1 U9961 (.Y(n12061), 
	.B1(n6419), 
	.B0(\ram[245][3] ), 
	.A1(n6438), 
	.A0(\ram[244][3] ));
   AOI22X1 U9962 (.Y(n12060), 
	.B1(n6457), 
	.B0(\ram[243][3] ), 
	.A1(n6476), 
	.A0(\ram[242][3] ));
   NAND4X1 U9963 (.Y(n12058), 
	.D(n12067), 
	.C(n12066), 
	.B(n12065), 
	.A(n12064));
   AOI22X1 U9964 (.Y(n12067), 
	.B1(n6495), 
	.B0(\ram[241][3] ), 
	.A1(n6514), 
	.A0(\ram[240][3] ));
   AOI22X1 U9965 (.Y(n12066), 
	.B1(n6533), 
	.B0(\ram[255][3] ), 
	.A1(n6553), 
	.A0(\ram[254][3] ));
   AOI22X1 U9966 (.Y(n12065), 
	.B1(n6572), 
	.B0(\ram[253][3] ), 
	.A1(n6591), 
	.A0(\ram[252][3] ));
   AOI22X1 U9967 (.Y(n12064), 
	.B1(n6610), 
	.B0(\ram[251][3] ), 
	.A1(n6629), 
	.A0(\ram[250][3] ));
   OAI21XL U9968 (.Y(n12045), 
	.B0(n7117), 
	.A1(n12069), 
	.A0(n12068));
   NAND4X1 U9969 (.Y(n12069), 
	.D(n12073), 
	.C(n12072), 
	.B(n12071), 
	.A(n12070));
   AOI22X1 U9970 (.Y(n12073), 
	.B1(n6342), 
	.B0(\ram[233][3] ), 
	.A1(n6362), 
	.A0(\ram[232][3] ));
   AOI22X1 U9971 (.Y(n12072), 
	.B1(n6381), 
	.B0(\ram[231][3] ), 
	.A1(n6400), 
	.A0(\ram[230][3] ));
   AOI22X1 U9972 (.Y(n12071), 
	.B1(n6419), 
	.B0(\ram[229][3] ), 
	.A1(n6438), 
	.A0(\ram[228][3] ));
   AOI22X1 U9973 (.Y(n12070), 
	.B1(n6457), 
	.B0(\ram[227][3] ), 
	.A1(n6476), 
	.A0(\ram[226][3] ));
   NAND4X1 U9974 (.Y(n12068), 
	.D(n12077), 
	.C(n12076), 
	.B(n12075), 
	.A(n12074));
   AOI22X1 U9975 (.Y(n12077), 
	.B1(n6495), 
	.B0(\ram[225][3] ), 
	.A1(n6514), 
	.A0(\ram[224][3] ));
   AOI22X1 U9976 (.Y(n12076), 
	.B1(n6533), 
	.B0(\ram[239][3] ), 
	.A1(n6553), 
	.A0(\ram[238][3] ));
   AOI22X1 U9977 (.Y(n12075), 
	.B1(n6572), 
	.B0(\ram[237][3] ), 
	.A1(n6591), 
	.A0(\ram[236][3] ));
   AOI22X1 U9978 (.Y(n12074), 
	.B1(n6610), 
	.B0(\ram[235][3] ), 
	.A1(n6629), 
	.A0(\ram[234][3] ));
   OAI21XL U9979 (.Y(n12044), 
	.B0(n7406), 
	.A1(n12079), 
	.A0(n12078));
   NAND4X1 U9980 (.Y(n12079), 
	.D(n12083), 
	.C(n12082), 
	.B(n12081), 
	.A(n12080));
   AOI22X1 U9981 (.Y(n12083), 
	.B1(n6342), 
	.B0(\ram[217][3] ), 
	.A1(n6362), 
	.A0(\ram[216][3] ));
   AOI22X1 U9982 (.Y(n12082), 
	.B1(n6381), 
	.B0(\ram[215][3] ), 
	.A1(n6400), 
	.A0(\ram[214][3] ));
   AOI22X1 U9983 (.Y(n12081), 
	.B1(n6419), 
	.B0(\ram[213][3] ), 
	.A1(n6438), 
	.A0(\ram[212][3] ));
   AOI22X1 U9984 (.Y(n12080), 
	.B1(n6457), 
	.B0(\ram[211][3] ), 
	.A1(n6476), 
	.A0(\ram[210][3] ));
   NAND4X1 U9985 (.Y(n12078), 
	.D(n12087), 
	.C(n12086), 
	.B(n12085), 
	.A(n12084));
   AOI22X1 U9986 (.Y(n12087), 
	.B1(n6495), 
	.B0(\ram[209][3] ), 
	.A1(n6514), 
	.A0(\ram[208][3] ));
   AOI22X1 U9987 (.Y(n12086), 
	.B1(n6533), 
	.B0(\ram[223][3] ), 
	.A1(n6553), 
	.A0(\ram[222][3] ));
   AOI22X1 U9988 (.Y(n12085), 
	.B1(n6572), 
	.B0(\ram[221][3] ), 
	.A1(n6591), 
	.A0(\ram[220][3] ));
   AOI22X1 U9989 (.Y(n12084), 
	.B1(n6610), 
	.B0(\ram[219][3] ), 
	.A1(n6629), 
	.A0(\ram[218][3] ));
   NAND4X1 U9990 (.Y(n12042), 
	.D(n12091), 
	.C(n12090), 
	.B(n12089), 
	.A(n12088));
   OAI21XL U9991 (.Y(n12091), 
	.B0(n7695), 
	.A1(n12093), 
	.A0(n12092));
   NAND4X1 U9992 (.Y(n12093), 
	.D(n12097), 
	.C(n12096), 
	.B(n12095), 
	.A(n12094));
   AOI22X1 U9993 (.Y(n12097), 
	.B1(n6342), 
	.B0(\ram[201][3] ), 
	.A1(n6362), 
	.A0(\ram[200][3] ));
   AOI22X1 U9994 (.Y(n12096), 
	.B1(n6381), 
	.B0(\ram[199][3] ), 
	.A1(n6400), 
	.A0(\ram[198][3] ));
   AOI22X1 U9995 (.Y(n12095), 
	.B1(n6419), 
	.B0(\ram[197][3] ), 
	.A1(n6438), 
	.A0(\ram[196][3] ));
   AOI22X1 U9996 (.Y(n12094), 
	.B1(n6457), 
	.B0(\ram[195][3] ), 
	.A1(n6476), 
	.A0(\ram[194][3] ));
   NAND4X1 U9997 (.Y(n12092), 
	.D(n12101), 
	.C(n12100), 
	.B(n12099), 
	.A(n12098));
   AOI22X1 U9998 (.Y(n12101), 
	.B1(n6495), 
	.B0(\ram[193][3] ), 
	.A1(n6514), 
	.A0(\ram[192][3] ));
   AOI22X1 U9999 (.Y(n12100), 
	.B1(n6533), 
	.B0(\ram[207][3] ), 
	.A1(n6553), 
	.A0(\ram[206][3] ));
   AOI22X1 U10000 (.Y(n12099), 
	.B1(n6572), 
	.B0(\ram[205][3] ), 
	.A1(n6591), 
	.A0(\ram[204][3] ));
   AOI22X1 U10001 (.Y(n12098), 
	.B1(n6610), 
	.B0(\ram[203][3] ), 
	.A1(n6629), 
	.A0(\ram[202][3] ));
   OAI21XL U10002 (.Y(n12090), 
	.B0(n7984), 
	.A1(n12103), 
	.A0(n12102));
   NAND4X1 U10003 (.Y(n12103), 
	.D(n12107), 
	.C(n12106), 
	.B(n12105), 
	.A(n12104));
   AOI22X1 U10004 (.Y(n12107), 
	.B1(n6342), 
	.B0(\ram[185][3] ), 
	.A1(n6362), 
	.A0(\ram[184][3] ));
   AOI22X1 U10005 (.Y(n12106), 
	.B1(n6381), 
	.B0(\ram[183][3] ), 
	.A1(n6400), 
	.A0(\ram[182][3] ));
   AOI22X1 U10006 (.Y(n12105), 
	.B1(n6419), 
	.B0(\ram[181][3] ), 
	.A1(n6438), 
	.A0(\ram[180][3] ));
   AOI22X1 U10007 (.Y(n12104), 
	.B1(n6457), 
	.B0(\ram[179][3] ), 
	.A1(n6476), 
	.A0(\ram[178][3] ));
   NAND4X1 U10008 (.Y(n12102), 
	.D(n12111), 
	.C(n12110), 
	.B(n12109), 
	.A(n12108));
   AOI22X1 U10009 (.Y(n12111), 
	.B1(n6495), 
	.B0(\ram[177][3] ), 
	.A1(n6514), 
	.A0(\ram[176][3] ));
   AOI22X1 U10010 (.Y(n12110), 
	.B1(n6533), 
	.B0(\ram[191][3] ), 
	.A1(n6553), 
	.A0(\ram[190][3] ));
   AOI22X1 U10011 (.Y(n12109), 
	.B1(n6572), 
	.B0(\ram[189][3] ), 
	.A1(n6591), 
	.A0(\ram[188][3] ));
   AOI22X1 U10012 (.Y(n12108), 
	.B1(n6610), 
	.B0(\ram[187][3] ), 
	.A1(n6629), 
	.A0(\ram[186][3] ));
   OAI21XL U10013 (.Y(n12089), 
	.B0(n8273), 
	.A1(n12113), 
	.A0(n12112));
   NAND4X1 U10014 (.Y(n12113), 
	.D(n12117), 
	.C(n12116), 
	.B(n12115), 
	.A(n12114));
   AOI22X1 U10015 (.Y(n12117), 
	.B1(n6342), 
	.B0(\ram[169][3] ), 
	.A1(n6362), 
	.A0(\ram[168][3] ));
   AOI22X1 U10016 (.Y(n12116), 
	.B1(n6381), 
	.B0(\ram[167][3] ), 
	.A1(n6400), 
	.A0(\ram[166][3] ));
   AOI22X1 U10017 (.Y(n12115), 
	.B1(n6419), 
	.B0(\ram[165][3] ), 
	.A1(n6438), 
	.A0(\ram[164][3] ));
   AOI22X1 U10018 (.Y(n12114), 
	.B1(n6457), 
	.B0(\ram[163][3] ), 
	.A1(n6476), 
	.A0(\ram[162][3] ));
   NAND4X1 U10019 (.Y(n12112), 
	.D(n12121), 
	.C(n12120), 
	.B(n12119), 
	.A(n12118));
   AOI22X1 U10020 (.Y(n12121), 
	.B1(n6495), 
	.B0(\ram[161][3] ), 
	.A1(n6514), 
	.A0(\ram[160][3] ));
   AOI22X1 U10021 (.Y(n12120), 
	.B1(n6533), 
	.B0(\ram[175][3] ), 
	.A1(n6553), 
	.A0(\ram[174][3] ));
   AOI22X1 U10022 (.Y(n12119), 
	.B1(n6572), 
	.B0(\ram[173][3] ), 
	.A1(n6591), 
	.A0(\ram[172][3] ));
   AOI22X1 U10023 (.Y(n12118), 
	.B1(n6610), 
	.B0(\ram[171][3] ), 
	.A1(n6629), 
	.A0(\ram[170][3] ));
   OAI21XL U10024 (.Y(n12088), 
	.B0(n8562), 
	.A1(n12123), 
	.A0(n12122));
   NAND4X1 U10025 (.Y(n12123), 
	.D(n12127), 
	.C(n12126), 
	.B(n12125), 
	.A(n12124));
   AOI22X1 U10026 (.Y(n12127), 
	.B1(n6342), 
	.B0(\ram[153][3] ), 
	.A1(n6362), 
	.A0(\ram[152][3] ));
   AOI22X1 U10027 (.Y(n12126), 
	.B1(n6381), 
	.B0(\ram[151][3] ), 
	.A1(n6400), 
	.A0(\ram[150][3] ));
   AOI22X1 U10028 (.Y(n12125), 
	.B1(n6419), 
	.B0(\ram[149][3] ), 
	.A1(n6438), 
	.A0(\ram[148][3] ));
   AOI22X1 U10029 (.Y(n12124), 
	.B1(n6457), 
	.B0(\ram[147][3] ), 
	.A1(n6476), 
	.A0(\ram[146][3] ));
   NAND4X1 U10030 (.Y(n12122), 
	.D(n12131), 
	.C(n12130), 
	.B(n12129), 
	.A(n12128));
   AOI22X1 U10031 (.Y(n12131), 
	.B1(n6495), 
	.B0(\ram[145][3] ), 
	.A1(n6514), 
	.A0(\ram[144][3] ));
   AOI22X1 U10032 (.Y(n12130), 
	.B1(n6533), 
	.B0(\ram[159][3] ), 
	.A1(n6553), 
	.A0(\ram[158][3] ));
   AOI22X1 U10033 (.Y(n12129), 
	.B1(n6572), 
	.B0(\ram[157][3] ), 
	.A1(n6591), 
	.A0(\ram[156][3] ));
   AOI22X1 U10034 (.Y(n12128), 
	.B1(n6610), 
	.B0(\ram[155][3] ), 
	.A1(n6629), 
	.A0(\ram[154][3] ));
   NAND4X1 U10035 (.Y(n12041), 
	.D(n12135), 
	.C(n12134), 
	.B(n12133), 
	.A(n12132));
   OAI21XL U10036 (.Y(n12135), 
	.B0(n8851), 
	.A1(n12137), 
	.A0(n12136));
   NAND4X1 U10037 (.Y(n12137), 
	.D(n12141), 
	.C(n12140), 
	.B(n12139), 
	.A(n12138));
   AOI22X1 U10038 (.Y(n12141), 
	.B1(n6342), 
	.B0(\ram[137][3] ), 
	.A1(n6362), 
	.A0(\ram[136][3] ));
   AOI22X1 U10039 (.Y(n12140), 
	.B1(n6381), 
	.B0(\ram[135][3] ), 
	.A1(n6400), 
	.A0(\ram[134][3] ));
   AOI22X1 U10040 (.Y(n12139), 
	.B1(n6419), 
	.B0(\ram[133][3] ), 
	.A1(n6438), 
	.A0(\ram[132][3] ));
   AOI22X1 U10041 (.Y(n12138), 
	.B1(n6457), 
	.B0(\ram[131][3] ), 
	.A1(n6476), 
	.A0(\ram[130][3] ));
   NAND4X1 U10042 (.Y(n12136), 
	.D(n12145), 
	.C(n12144), 
	.B(n12143), 
	.A(n12142));
   AOI22X1 U10043 (.Y(n12145), 
	.B1(n6495), 
	.B0(\ram[129][3] ), 
	.A1(n6514), 
	.A0(\ram[128][3] ));
   AOI22X1 U10044 (.Y(n12144), 
	.B1(n6533), 
	.B0(\ram[143][3] ), 
	.A1(n6553), 
	.A0(\ram[142][3] ));
   AOI22X1 U10045 (.Y(n12143), 
	.B1(n6572), 
	.B0(\ram[141][3] ), 
	.A1(n6591), 
	.A0(\ram[140][3] ));
   AOI22X1 U10046 (.Y(n12142), 
	.B1(n6610), 
	.B0(\ram[139][3] ), 
	.A1(n6629), 
	.A0(\ram[138][3] ));
   OAI21XL U10047 (.Y(n12134), 
	.B0(n9140), 
	.A1(n12147), 
	.A0(n12146));
   NAND4X1 U10048 (.Y(n12147), 
	.D(n12151), 
	.C(n12150), 
	.B(n12149), 
	.A(n12148));
   AOI22X1 U10049 (.Y(n12151), 
	.B1(n6342), 
	.B0(\ram[121][3] ), 
	.A1(n6362), 
	.A0(\ram[120][3] ));
   AOI22X1 U10050 (.Y(n12150), 
	.B1(n6381), 
	.B0(\ram[119][3] ), 
	.A1(n6400), 
	.A0(\ram[118][3] ));
   AOI22X1 U10051 (.Y(n12149), 
	.B1(n6419), 
	.B0(\ram[117][3] ), 
	.A1(n6438), 
	.A0(\ram[116][3] ));
   AOI22X1 U10052 (.Y(n12148), 
	.B1(n6457), 
	.B0(\ram[115][3] ), 
	.A1(n6476), 
	.A0(\ram[114][3] ));
   NAND4X1 U10053 (.Y(n12146), 
	.D(n12155), 
	.C(n12154), 
	.B(n12153), 
	.A(n12152));
   AOI22X1 U10054 (.Y(n12155), 
	.B1(n6495), 
	.B0(\ram[113][3] ), 
	.A1(n6514), 
	.A0(\ram[112][3] ));
   AOI22X1 U10055 (.Y(n12154), 
	.B1(n6533), 
	.B0(\ram[127][3] ), 
	.A1(n6553), 
	.A0(\ram[126][3] ));
   AOI22X1 U10056 (.Y(n12153), 
	.B1(n6572), 
	.B0(\ram[125][3] ), 
	.A1(n6591), 
	.A0(\ram[124][3] ));
   AOI22X1 U10057 (.Y(n12152), 
	.B1(n6610), 
	.B0(\ram[123][3] ), 
	.A1(n6629), 
	.A0(\ram[122][3] ));
   OAI21XL U10058 (.Y(n12133), 
	.B0(n9429), 
	.A1(n12157), 
	.A0(n12156));
   NAND4X1 U10059 (.Y(n12157), 
	.D(n12161), 
	.C(n12160), 
	.B(n12159), 
	.A(n12158));
   AOI22X1 U10060 (.Y(n12161), 
	.B1(n6342), 
	.B0(\ram[105][3] ), 
	.A1(n6362), 
	.A0(\ram[104][3] ));
   AOI22X1 U10061 (.Y(n12160), 
	.B1(n6381), 
	.B0(\ram[103][3] ), 
	.A1(n6400), 
	.A0(\ram[102][3] ));
   AOI22X1 U10062 (.Y(n12159), 
	.B1(n6419), 
	.B0(\ram[101][3] ), 
	.A1(n6438), 
	.A0(\ram[100][3] ));
   AOI22X1 U10063 (.Y(n12158), 
	.B1(n6457), 
	.B0(\ram[99][3] ), 
	.A1(n6476), 
	.A0(\ram[98][3] ));
   NAND4X1 U10064 (.Y(n12156), 
	.D(n12165), 
	.C(n12164), 
	.B(n12163), 
	.A(n12162));
   AOI22X1 U10065 (.Y(n12165), 
	.B1(n6495), 
	.B0(\ram[97][3] ), 
	.A1(n6514), 
	.A0(\ram[96][3] ));
   AOI22X1 U10066 (.Y(n12164), 
	.B1(n6533), 
	.B0(\ram[111][3] ), 
	.A1(n6553), 
	.A0(\ram[110][3] ));
   AOI22X1 U10067 (.Y(n12163), 
	.B1(n6572), 
	.B0(\ram[109][3] ), 
	.A1(n6591), 
	.A0(\ram[108][3] ));
   AOI22X1 U10068 (.Y(n12162), 
	.B1(n6610), 
	.B0(\ram[107][3] ), 
	.A1(n6629), 
	.A0(\ram[106][3] ));
   OAI21XL U10069 (.Y(n12132), 
	.B0(n9718), 
	.A1(n12167), 
	.A0(n12166));
   NAND4X1 U10070 (.Y(n12167), 
	.D(n12171), 
	.C(n12170), 
	.B(n12169), 
	.A(n12168));
   AOI22X1 U10071 (.Y(n12171), 
	.B1(n6342), 
	.B0(\ram[89][3] ), 
	.A1(n6362), 
	.A0(\ram[88][3] ));
   AOI22X1 U10072 (.Y(n12170), 
	.B1(n6381), 
	.B0(\ram[87][3] ), 
	.A1(n6400), 
	.A0(\ram[86][3] ));
   AOI22X1 U10073 (.Y(n12169), 
	.B1(n6419), 
	.B0(\ram[85][3] ), 
	.A1(n6438), 
	.A0(\ram[84][3] ));
   AOI22X1 U10074 (.Y(n12168), 
	.B1(n6457), 
	.B0(\ram[83][3] ), 
	.A1(n6476), 
	.A0(\ram[82][3] ));
   NAND4X1 U10075 (.Y(n12166), 
	.D(n12175), 
	.C(n12174), 
	.B(n12173), 
	.A(n12172));
   AOI22X1 U10076 (.Y(n12175), 
	.B1(n6495), 
	.B0(\ram[81][3] ), 
	.A1(n6514), 
	.A0(\ram[80][3] ));
   AOI22X1 U10077 (.Y(n12174), 
	.B1(n6533), 
	.B0(\ram[95][3] ), 
	.A1(n6553), 
	.A0(\ram[94][3] ));
   AOI22X1 U10078 (.Y(n12173), 
	.B1(n6572), 
	.B0(\ram[93][3] ), 
	.A1(n6591), 
	.A0(\ram[92][3] ));
   AOI22X1 U10079 (.Y(n12172), 
	.B1(n6610), 
	.B0(\ram[91][3] ), 
	.A1(n6629), 
	.A0(\ram[90][3] ));
   NAND4X1 U10080 (.Y(n12040), 
	.D(n12179), 
	.C(n12178), 
	.B(n12177), 
	.A(n12176));
   OAI21XL U10081 (.Y(n12179), 
	.B0(n10007), 
	.A1(n12181), 
	.A0(n12180));
   NAND4X1 U10082 (.Y(n12181), 
	.D(n12185), 
	.C(n12184), 
	.B(n12183), 
	.A(n12182));
   AOI22X1 U10083 (.Y(n12185), 
	.B1(n6342), 
	.B0(\ram[73][3] ), 
	.A1(n6362), 
	.A0(\ram[72][3] ));
   AOI22X1 U10084 (.Y(n12184), 
	.B1(n6381), 
	.B0(\ram[71][3] ), 
	.A1(n6400), 
	.A0(\ram[70][3] ));
   AOI22X1 U10085 (.Y(n12183), 
	.B1(n6419), 
	.B0(\ram[69][3] ), 
	.A1(n6438), 
	.A0(\ram[68][3] ));
   AOI22X1 U10086 (.Y(n12182), 
	.B1(n6457), 
	.B0(\ram[67][3] ), 
	.A1(n6476), 
	.A0(\ram[66][3] ));
   NAND4X1 U10087 (.Y(n12180), 
	.D(n12189), 
	.C(n12188), 
	.B(n12187), 
	.A(n12186));
   AOI22X1 U10088 (.Y(n12189), 
	.B1(n6495), 
	.B0(\ram[65][3] ), 
	.A1(n6514), 
	.A0(\ram[64][3] ));
   AOI22X1 U10089 (.Y(n12188), 
	.B1(n6533), 
	.B0(\ram[79][3] ), 
	.A1(n6553), 
	.A0(\ram[78][3] ));
   AOI22X1 U10090 (.Y(n12187), 
	.B1(n6572), 
	.B0(\ram[77][3] ), 
	.A1(n6591), 
	.A0(\ram[76][3] ));
   AOI22X1 U10091 (.Y(n12186), 
	.B1(n6610), 
	.B0(\ram[75][3] ), 
	.A1(n6629), 
	.A0(\ram[74][3] ));
   OAI21XL U10092 (.Y(n12178), 
	.B0(n10296), 
	.A1(n12191), 
	.A0(n12190));
   NAND4X1 U10093 (.Y(n12191), 
	.D(n12195), 
	.C(n12194), 
	.B(n12193), 
	.A(n12192));
   AOI22X1 U10094 (.Y(n12195), 
	.B1(n6342), 
	.B0(\ram[57][3] ), 
	.A1(n6362), 
	.A0(\ram[56][3] ));
   AOI22X1 U10095 (.Y(n12194), 
	.B1(n6381), 
	.B0(\ram[55][3] ), 
	.A1(n6400), 
	.A0(\ram[54][3] ));
   AOI22X1 U10096 (.Y(n12193), 
	.B1(n6419), 
	.B0(\ram[53][3] ), 
	.A1(n6438), 
	.A0(\ram[52][3] ));
   AOI22X1 U10097 (.Y(n12192), 
	.B1(n6457), 
	.B0(\ram[51][3] ), 
	.A1(n6476), 
	.A0(\ram[50][3] ));
   NAND4X1 U10098 (.Y(n12190), 
	.D(n12199), 
	.C(n12198), 
	.B(n12197), 
	.A(n12196));
   AOI22X1 U10099 (.Y(n12199), 
	.B1(n6495), 
	.B0(\ram[49][3] ), 
	.A1(n6514), 
	.A0(\ram[48][3] ));
   AOI22X1 U10100 (.Y(n12198), 
	.B1(n6533), 
	.B0(\ram[63][3] ), 
	.A1(n6553), 
	.A0(\ram[62][3] ));
   AOI22X1 U10101 (.Y(n12197), 
	.B1(n6572), 
	.B0(\ram[61][3] ), 
	.A1(n6591), 
	.A0(\ram[60][3] ));
   AOI22X1 U10102 (.Y(n12196), 
	.B1(n6610), 
	.B0(\ram[59][3] ), 
	.A1(n6629), 
	.A0(\ram[58][3] ));
   OAI21XL U10103 (.Y(n12177), 
	.B0(n10585), 
	.A1(n12201), 
	.A0(n12200));
   NAND4X1 U10104 (.Y(n12201), 
	.D(n12205), 
	.C(n12204), 
	.B(n12203), 
	.A(n12202));
   AOI22X1 U10105 (.Y(n12205), 
	.B1(n6342), 
	.B0(\ram[41][3] ), 
	.A1(n6362), 
	.A0(\ram[40][3] ));
   AOI22X1 U10106 (.Y(n12204), 
	.B1(n6381), 
	.B0(\ram[39][3] ), 
	.A1(n6400), 
	.A0(\ram[38][3] ));
   AOI22X1 U10107 (.Y(n12203), 
	.B1(n6419), 
	.B0(\ram[37][3] ), 
	.A1(n6438), 
	.A0(\ram[36][3] ));
   AOI22X1 U10108 (.Y(n12202), 
	.B1(n6457), 
	.B0(\ram[35][3] ), 
	.A1(n6476), 
	.A0(\ram[34][3] ));
   NAND4X1 U10109 (.Y(n12200), 
	.D(n12209), 
	.C(n12208), 
	.B(n12207), 
	.A(n12206));
   AOI22X1 U10110 (.Y(n12209), 
	.B1(n6495), 
	.B0(\ram[33][3] ), 
	.A1(n6514), 
	.A0(\ram[32][3] ));
   AOI22X1 U10111 (.Y(n12208), 
	.B1(n6533), 
	.B0(\ram[47][3] ), 
	.A1(n6553), 
	.A0(\ram[46][3] ));
   AOI22X1 U10112 (.Y(n12207), 
	.B1(n6572), 
	.B0(\ram[45][3] ), 
	.A1(n6591), 
	.A0(\ram[44][3] ));
   AOI22X1 U10113 (.Y(n12206), 
	.B1(n6610), 
	.B0(\ram[43][3] ), 
	.A1(n6629), 
	.A0(\ram[42][3] ));
   OAI21XL U10114 (.Y(n12176), 
	.B0(n6343), 
	.A1(n12211), 
	.A0(n12210));
   NAND4X1 U10115 (.Y(n12211), 
	.D(n12215), 
	.C(n12214), 
	.B(n12213), 
	.A(n12212));
   AOI22X1 U10116 (.Y(n12215), 
	.B1(n6342), 
	.B0(\ram[25][3] ), 
	.A1(n6362), 
	.A0(\ram[24][3] ));
   AOI22X1 U10117 (.Y(n12214), 
	.B1(n6381), 
	.B0(\ram[23][3] ), 
	.A1(n6400), 
	.A0(\ram[22][3] ));
   AOI22X1 U10118 (.Y(n12213), 
	.B1(n6419), 
	.B0(\ram[21][3] ), 
	.A1(n6438), 
	.A0(\ram[20][3] ));
   AOI22X1 U10119 (.Y(n12212), 
	.B1(n6457), 
	.B0(\ram[19][3] ), 
	.A1(n6476), 
	.A0(\ram[18][3] ));
   NAND4X1 U10120 (.Y(n12210), 
	.D(n12219), 
	.C(n12218), 
	.B(n12217), 
	.A(n12216));
   AOI22X1 U10121 (.Y(n12219), 
	.B1(n6495), 
	.B0(\ram[17][3] ), 
	.A1(n6514), 
	.A0(\ram[16][3] ));
   AOI22X1 U10122 (.Y(n12218), 
	.B1(n6533), 
	.B0(\ram[31][3] ), 
	.A1(n6553), 
	.A0(\ram[30][3] ));
   AOI22X1 U10123 (.Y(n12217), 
	.B1(n6572), 
	.B0(\ram[29][3] ), 
	.A1(n6591), 
	.A0(\ram[28][3] ));
   AOI22X1 U10124 (.Y(n12216), 
	.B1(n6610), 
	.B0(\ram[27][3] ), 
	.A1(n6629), 
	.A0(\ram[26][3] ));
   OR4X1 U10125 (.Y(mem_read_data[2]), 
	.D(n12223), 
	.C(n12222), 
	.B(n12221), 
	.A(n12220));
   NAND4X1 U10126 (.Y(n12223), 
	.D(n12227), 
	.C(n12226), 
	.B(n12225), 
	.A(n12224));
   OAI21XL U10127 (.Y(n12227), 
	.B0(n6534), 
	.A1(n12229), 
	.A0(n12228));
   NAND4X1 U10128 (.Y(n12229), 
	.D(n12233), 
	.C(n12232), 
	.B(n12231), 
	.A(n12230));
   AOI22X1 U10129 (.Y(n12233), 
	.B1(n6342), 
	.B0(\ram[9][2] ), 
	.A1(n6362), 
	.A0(\ram[8][2] ));
   AOI22X1 U10130 (.Y(n12232), 
	.B1(n6381), 
	.B0(\ram[7][2] ), 
	.A1(n6400), 
	.A0(\ram[6][2] ));
   AOI22X1 U10131 (.Y(n12231), 
	.B1(n6419), 
	.B0(\ram[5][2] ), 
	.A1(n6438), 
	.A0(\ram[4][2] ));
   AOI22X1 U10132 (.Y(n12230), 
	.B1(n6457), 
	.B0(\ram[3][2] ), 
	.A1(n6476), 
	.A0(\ram[2][2] ));
   NAND4X1 U10133 (.Y(n12228), 
	.D(n12237), 
	.C(n12236), 
	.B(n12235), 
	.A(n12234));
   AOI22X1 U10134 (.Y(n12237), 
	.B1(n6495), 
	.B0(\ram[1][2] ), 
	.A1(n6514), 
	.A0(\ram[0][2] ));
   AOI22X1 U10135 (.Y(n12236), 
	.B1(n6533), 
	.B0(\ram[15][2] ), 
	.A1(n6553), 
	.A0(\ram[14][2] ));
   AOI22X1 U10136 (.Y(n12235), 
	.B1(n6572), 
	.B0(\ram[13][2] ), 
	.A1(n6591), 
	.A0(\ram[12][2] ));
   AOI22X1 U10137 (.Y(n12234), 
	.B1(n6610), 
	.B0(\ram[11][2] ), 
	.A1(n6629), 
	.A0(\ram[10][2] ));
   OAI21XL U10138 (.Y(n12226), 
	.B0(n6828), 
	.A1(n12239), 
	.A0(n12238));
   NAND4X1 U10139 (.Y(n12239), 
	.D(n12243), 
	.C(n12242), 
	.B(n12241), 
	.A(n12240));
   AOI22X1 U10140 (.Y(n12243), 
	.B1(n6342), 
	.B0(\ram[249][2] ), 
	.A1(n6362), 
	.A0(\ram[248][2] ));
   AOI22X1 U10141 (.Y(n12242), 
	.B1(n6381), 
	.B0(\ram[247][2] ), 
	.A1(n6400), 
	.A0(\ram[246][2] ));
   AOI22X1 U10142 (.Y(n12241), 
	.B1(n6419), 
	.B0(\ram[245][2] ), 
	.A1(n6438), 
	.A0(\ram[244][2] ));
   AOI22X1 U10143 (.Y(n12240), 
	.B1(n6457), 
	.B0(\ram[243][2] ), 
	.A1(n6476), 
	.A0(\ram[242][2] ));
   NAND4X1 U10144 (.Y(n12238), 
	.D(n12247), 
	.C(n12246), 
	.B(n12245), 
	.A(n12244));
   AOI22X1 U10145 (.Y(n12247), 
	.B1(n6495), 
	.B0(\ram[241][2] ), 
	.A1(n6514), 
	.A0(\ram[240][2] ));
   AOI22X1 U10146 (.Y(n12246), 
	.B1(n6533), 
	.B0(\ram[255][2] ), 
	.A1(n6553), 
	.A0(\ram[254][2] ));
   AOI22X1 U10147 (.Y(n12245), 
	.B1(n6572), 
	.B0(\ram[253][2] ), 
	.A1(n6591), 
	.A0(\ram[252][2] ));
   AOI22X1 U10148 (.Y(n12244), 
	.B1(n6610), 
	.B0(\ram[251][2] ), 
	.A1(n6629), 
	.A0(\ram[250][2] ));
   OAI21XL U10149 (.Y(n12225), 
	.B0(n7117), 
	.A1(n12249), 
	.A0(n12248));
   NAND4X1 U10150 (.Y(n12249), 
	.D(n12253), 
	.C(n12252), 
	.B(n12251), 
	.A(n12250));
   AOI22X1 U10151 (.Y(n12253), 
	.B1(n6342), 
	.B0(\ram[233][2] ), 
	.A1(n6362), 
	.A0(\ram[232][2] ));
   AOI22X1 U10152 (.Y(n12252), 
	.B1(n6381), 
	.B0(\ram[231][2] ), 
	.A1(n6400), 
	.A0(\ram[230][2] ));
   AOI22X1 U10153 (.Y(n12251), 
	.B1(n6419), 
	.B0(\ram[229][2] ), 
	.A1(n6438), 
	.A0(\ram[228][2] ));
   AOI22X1 U10154 (.Y(n12250), 
	.B1(n6457), 
	.B0(\ram[227][2] ), 
	.A1(n6476), 
	.A0(\ram[226][2] ));
   NAND4X1 U10155 (.Y(n12248), 
	.D(n12257), 
	.C(n12256), 
	.B(n12255), 
	.A(n12254));
   AOI22X1 U10156 (.Y(n12257), 
	.B1(n6495), 
	.B0(\ram[225][2] ), 
	.A1(n6514), 
	.A0(\ram[224][2] ));
   AOI22X1 U10157 (.Y(n12256), 
	.B1(n6533), 
	.B0(\ram[239][2] ), 
	.A1(n6553), 
	.A0(\ram[238][2] ));
   AOI22X1 U10158 (.Y(n12255), 
	.B1(n6572), 
	.B0(\ram[237][2] ), 
	.A1(n6591), 
	.A0(\ram[236][2] ));
   AOI22X1 U10159 (.Y(n12254), 
	.B1(n6610), 
	.B0(\ram[235][2] ), 
	.A1(n6629), 
	.A0(\ram[234][2] ));
   OAI21XL U10160 (.Y(n12224), 
	.B0(n7406), 
	.A1(n12259), 
	.A0(n12258));
   NAND4X1 U10161 (.Y(n12259), 
	.D(n12263), 
	.C(n12262), 
	.B(n12261), 
	.A(n12260));
   AOI22X1 U10162 (.Y(n12263), 
	.B1(n6342), 
	.B0(\ram[217][2] ), 
	.A1(n6362), 
	.A0(\ram[216][2] ));
   AOI22X1 U10163 (.Y(n12262), 
	.B1(n6381), 
	.B0(\ram[215][2] ), 
	.A1(n6400), 
	.A0(\ram[214][2] ));
   AOI22X1 U10164 (.Y(n12261), 
	.B1(n6419), 
	.B0(\ram[213][2] ), 
	.A1(n6438), 
	.A0(\ram[212][2] ));
   AOI22X1 U10165 (.Y(n12260), 
	.B1(n6457), 
	.B0(\ram[211][2] ), 
	.A1(n6476), 
	.A0(\ram[210][2] ));
   NAND4X1 U10166 (.Y(n12258), 
	.D(n12267), 
	.C(n12266), 
	.B(n12265), 
	.A(n12264));
   AOI22X1 U10167 (.Y(n12267), 
	.B1(n6495), 
	.B0(\ram[209][2] ), 
	.A1(n6514), 
	.A0(\ram[208][2] ));
   AOI22X1 U10168 (.Y(n12266), 
	.B1(n6533), 
	.B0(\ram[223][2] ), 
	.A1(n6553), 
	.A0(\ram[222][2] ));
   AOI22X1 U10169 (.Y(n12265), 
	.B1(n6572), 
	.B0(\ram[221][2] ), 
	.A1(n6591), 
	.A0(\ram[220][2] ));
   AOI22X1 U10170 (.Y(n12264), 
	.B1(n6610), 
	.B0(\ram[219][2] ), 
	.A1(n6629), 
	.A0(\ram[218][2] ));
   NAND4X1 U10171 (.Y(n12222), 
	.D(n12271), 
	.C(n12270), 
	.B(n12269), 
	.A(n12268));
   OAI21XL U10172 (.Y(n12271), 
	.B0(n7695), 
	.A1(n12273), 
	.A0(n12272));
   NAND4X1 U10173 (.Y(n12273), 
	.D(n12277), 
	.C(n12276), 
	.B(n12275), 
	.A(n12274));
   AOI22X1 U10174 (.Y(n12277), 
	.B1(n6342), 
	.B0(\ram[201][2] ), 
	.A1(n6362), 
	.A0(\ram[200][2] ));
   AOI22X1 U10175 (.Y(n12276), 
	.B1(n6381), 
	.B0(\ram[199][2] ), 
	.A1(n6400), 
	.A0(\ram[198][2] ));
   AOI22X1 U10176 (.Y(n12275), 
	.B1(n6419), 
	.B0(\ram[197][2] ), 
	.A1(n6438), 
	.A0(\ram[196][2] ));
   AOI22X1 U10177 (.Y(n12274), 
	.B1(n6457), 
	.B0(\ram[195][2] ), 
	.A1(n6476), 
	.A0(\ram[194][2] ));
   NAND4X1 U10178 (.Y(n12272), 
	.D(n12281), 
	.C(n12280), 
	.B(n12279), 
	.A(n12278));
   AOI22X1 U10179 (.Y(n12281), 
	.B1(n6495), 
	.B0(\ram[193][2] ), 
	.A1(n6514), 
	.A0(\ram[192][2] ));
   AOI22X1 U10180 (.Y(n12280), 
	.B1(n6533), 
	.B0(\ram[207][2] ), 
	.A1(n6553), 
	.A0(\ram[206][2] ));
   AOI22X1 U10181 (.Y(n12279), 
	.B1(n6572), 
	.B0(\ram[205][2] ), 
	.A1(n6591), 
	.A0(\ram[204][2] ));
   AOI22X1 U10182 (.Y(n12278), 
	.B1(n6610), 
	.B0(\ram[203][2] ), 
	.A1(n6629), 
	.A0(\ram[202][2] ));
   OAI21XL U10183 (.Y(n12270), 
	.B0(n7984), 
	.A1(n12283), 
	.A0(n12282));
   NAND4X1 U10184 (.Y(n12283), 
	.D(n12287), 
	.C(n12286), 
	.B(n12285), 
	.A(n12284));
   AOI22X1 U10185 (.Y(n12287), 
	.B1(n6342), 
	.B0(\ram[185][2] ), 
	.A1(n6362), 
	.A0(\ram[184][2] ));
   AOI22X1 U10186 (.Y(n12286), 
	.B1(n6381), 
	.B0(\ram[183][2] ), 
	.A1(n6400), 
	.A0(\ram[182][2] ));
   AOI22X1 U10187 (.Y(n12285), 
	.B1(n6419), 
	.B0(\ram[181][2] ), 
	.A1(n6438), 
	.A0(\ram[180][2] ));
   AOI22X1 U10188 (.Y(n12284), 
	.B1(n6457), 
	.B0(\ram[179][2] ), 
	.A1(n6476), 
	.A0(\ram[178][2] ));
   NAND4X1 U10189 (.Y(n12282), 
	.D(n12291), 
	.C(n12290), 
	.B(n12289), 
	.A(n12288));
   AOI22X1 U10190 (.Y(n12291), 
	.B1(n6495), 
	.B0(\ram[177][2] ), 
	.A1(n6514), 
	.A0(\ram[176][2] ));
   AOI22X1 U10191 (.Y(n12290), 
	.B1(n6533), 
	.B0(\ram[191][2] ), 
	.A1(n6553), 
	.A0(\ram[190][2] ));
   AOI22X1 U10192 (.Y(n12289), 
	.B1(n6572), 
	.B0(\ram[189][2] ), 
	.A1(n6591), 
	.A0(\ram[188][2] ));
   AOI22X1 U10193 (.Y(n12288), 
	.B1(n6610), 
	.B0(\ram[187][2] ), 
	.A1(n6629), 
	.A0(\ram[186][2] ));
   OAI21XL U10194 (.Y(n12269), 
	.B0(n8273), 
	.A1(n12293), 
	.A0(n12292));
   NAND4X1 U10195 (.Y(n12293), 
	.D(n12297), 
	.C(n12296), 
	.B(n12295), 
	.A(n12294));
   AOI22X1 U10196 (.Y(n12297), 
	.B1(n6342), 
	.B0(\ram[169][2] ), 
	.A1(n6362), 
	.A0(\ram[168][2] ));
   AOI22X1 U10197 (.Y(n12296), 
	.B1(n6381), 
	.B0(\ram[167][2] ), 
	.A1(n6400), 
	.A0(\ram[166][2] ));
   AOI22X1 U10198 (.Y(n12295), 
	.B1(n6419), 
	.B0(\ram[165][2] ), 
	.A1(n6438), 
	.A0(\ram[164][2] ));
   AOI22X1 U10199 (.Y(n12294), 
	.B1(n6457), 
	.B0(\ram[163][2] ), 
	.A1(n6476), 
	.A0(\ram[162][2] ));
   NAND4X1 U10200 (.Y(n12292), 
	.D(n12301), 
	.C(n12300), 
	.B(n12299), 
	.A(n12298));
   AOI22X1 U10201 (.Y(n12301), 
	.B1(n6495), 
	.B0(\ram[161][2] ), 
	.A1(n6514), 
	.A0(\ram[160][2] ));
   AOI22X1 U10202 (.Y(n12300), 
	.B1(n6533), 
	.B0(\ram[175][2] ), 
	.A1(n6553), 
	.A0(\ram[174][2] ));
   AOI22X1 U10203 (.Y(n12299), 
	.B1(n6572), 
	.B0(\ram[173][2] ), 
	.A1(n6591), 
	.A0(\ram[172][2] ));
   AOI22X1 U10204 (.Y(n12298), 
	.B1(n6610), 
	.B0(\ram[171][2] ), 
	.A1(n6629), 
	.A0(\ram[170][2] ));
   OAI21XL U10205 (.Y(n12268), 
	.B0(n8562), 
	.A1(n12303), 
	.A0(n12302));
   NAND4X1 U10206 (.Y(n12303), 
	.D(n12307), 
	.C(n12306), 
	.B(n12305), 
	.A(n12304));
   AOI22X1 U10207 (.Y(n12307), 
	.B1(n6342), 
	.B0(\ram[153][2] ), 
	.A1(n6362), 
	.A0(\ram[152][2] ));
   AOI22X1 U10208 (.Y(n12306), 
	.B1(n6381), 
	.B0(\ram[151][2] ), 
	.A1(n6400), 
	.A0(\ram[150][2] ));
   AOI22X1 U10209 (.Y(n12305), 
	.B1(n6419), 
	.B0(\ram[149][2] ), 
	.A1(n6438), 
	.A0(\ram[148][2] ));
   AOI22X1 U10210 (.Y(n12304), 
	.B1(n6457), 
	.B0(\ram[147][2] ), 
	.A1(n6476), 
	.A0(\ram[146][2] ));
   NAND4X1 U10211 (.Y(n12302), 
	.D(n12311), 
	.C(n12310), 
	.B(n12309), 
	.A(n12308));
   AOI22X1 U10212 (.Y(n12311), 
	.B1(n6495), 
	.B0(\ram[145][2] ), 
	.A1(n6514), 
	.A0(\ram[144][2] ));
   AOI22X1 U10213 (.Y(n12310), 
	.B1(n6533), 
	.B0(\ram[159][2] ), 
	.A1(n6553), 
	.A0(\ram[158][2] ));
   AOI22X1 U10214 (.Y(n12309), 
	.B1(n6572), 
	.B0(\ram[157][2] ), 
	.A1(n6591), 
	.A0(\ram[156][2] ));
   AOI22X1 U10215 (.Y(n12308), 
	.B1(n6610), 
	.B0(\ram[155][2] ), 
	.A1(n6629), 
	.A0(\ram[154][2] ));
   NAND4X1 U10216 (.Y(n12221), 
	.D(n12315), 
	.C(n12314), 
	.B(n12313), 
	.A(n12312));
   OAI21XL U10217 (.Y(n12315), 
	.B0(n8851), 
	.A1(n12317), 
	.A0(n12316));
   NAND4X1 U10218 (.Y(n12317), 
	.D(n12321), 
	.C(n12320), 
	.B(n12319), 
	.A(n12318));
   AOI22X1 U10219 (.Y(n12321), 
	.B1(n6342), 
	.B0(\ram[137][2] ), 
	.A1(n6362), 
	.A0(\ram[136][2] ));
   AOI22X1 U10220 (.Y(n12320), 
	.B1(n6381), 
	.B0(\ram[135][2] ), 
	.A1(n6400), 
	.A0(\ram[134][2] ));
   AOI22X1 U10221 (.Y(n12319), 
	.B1(n6419), 
	.B0(\ram[133][2] ), 
	.A1(n6438), 
	.A0(\ram[132][2] ));
   AOI22X1 U10222 (.Y(n12318), 
	.B1(n6457), 
	.B0(\ram[131][2] ), 
	.A1(n6476), 
	.A0(\ram[130][2] ));
   NAND4X1 U10223 (.Y(n12316), 
	.D(n12325), 
	.C(n12324), 
	.B(n12323), 
	.A(n12322));
   AOI22X1 U10224 (.Y(n12325), 
	.B1(n6495), 
	.B0(\ram[129][2] ), 
	.A1(n6514), 
	.A0(\ram[128][2] ));
   AOI22X1 U10225 (.Y(n12324), 
	.B1(n6533), 
	.B0(\ram[143][2] ), 
	.A1(n6553), 
	.A0(\ram[142][2] ));
   AOI22X1 U10226 (.Y(n12323), 
	.B1(n6572), 
	.B0(\ram[141][2] ), 
	.A1(n6591), 
	.A0(\ram[140][2] ));
   AOI22X1 U10227 (.Y(n12322), 
	.B1(n6610), 
	.B0(\ram[139][2] ), 
	.A1(n6629), 
	.A0(\ram[138][2] ));
   OAI21XL U10228 (.Y(n12314), 
	.B0(n9140), 
	.A1(n12327), 
	.A0(n12326));
   NAND4X1 U10229 (.Y(n12327), 
	.D(n12331), 
	.C(n12330), 
	.B(n12329), 
	.A(n12328));
   AOI22X1 U10230 (.Y(n12331), 
	.B1(n6342), 
	.B0(\ram[121][2] ), 
	.A1(n6362), 
	.A0(\ram[120][2] ));
   AOI22X1 U10231 (.Y(n12330), 
	.B1(n6381), 
	.B0(\ram[119][2] ), 
	.A1(n6400), 
	.A0(\ram[118][2] ));
   AOI22X1 U10232 (.Y(n12329), 
	.B1(n6419), 
	.B0(\ram[117][2] ), 
	.A1(n6438), 
	.A0(\ram[116][2] ));
   AOI22X1 U10233 (.Y(n12328), 
	.B1(n6457), 
	.B0(\ram[115][2] ), 
	.A1(n6476), 
	.A0(\ram[114][2] ));
   NAND4X1 U10234 (.Y(n12326), 
	.D(n12335), 
	.C(n12334), 
	.B(n12333), 
	.A(n12332));
   AOI22X1 U10235 (.Y(n12335), 
	.B1(n6495), 
	.B0(\ram[113][2] ), 
	.A1(n6514), 
	.A0(\ram[112][2] ));
   AOI22X1 U10236 (.Y(n12334), 
	.B1(n6533), 
	.B0(\ram[127][2] ), 
	.A1(n6553), 
	.A0(\ram[126][2] ));
   AOI22X1 U10237 (.Y(n12333), 
	.B1(n6572), 
	.B0(\ram[125][2] ), 
	.A1(n6591), 
	.A0(\ram[124][2] ));
   AOI22X1 U10238 (.Y(n12332), 
	.B1(n6610), 
	.B0(\ram[123][2] ), 
	.A1(n6629), 
	.A0(\ram[122][2] ));
   OAI21XL U10239 (.Y(n12313), 
	.B0(n9429), 
	.A1(n12337), 
	.A0(n12336));
   NAND4X1 U10240 (.Y(n12337), 
	.D(n12341), 
	.C(n12340), 
	.B(n12339), 
	.A(n12338));
   AOI22X1 U10241 (.Y(n12341), 
	.B1(n6342), 
	.B0(\ram[105][2] ), 
	.A1(n6362), 
	.A0(\ram[104][2] ));
   AOI22X1 U10242 (.Y(n12340), 
	.B1(n6381), 
	.B0(\ram[103][2] ), 
	.A1(n6400), 
	.A0(\ram[102][2] ));
   AOI22X1 U10243 (.Y(n12339), 
	.B1(n6419), 
	.B0(\ram[101][2] ), 
	.A1(n6438), 
	.A0(\ram[100][2] ));
   AOI22X1 U10244 (.Y(n12338), 
	.B1(n6457), 
	.B0(\ram[99][2] ), 
	.A1(n6476), 
	.A0(\ram[98][2] ));
   NAND4X1 U10245 (.Y(n12336), 
	.D(n12345), 
	.C(n12344), 
	.B(n12343), 
	.A(n12342));
   AOI22X1 U10246 (.Y(n12345), 
	.B1(n6495), 
	.B0(\ram[97][2] ), 
	.A1(n6514), 
	.A0(\ram[96][2] ));
   AOI22X1 U10247 (.Y(n12344), 
	.B1(n6533), 
	.B0(\ram[111][2] ), 
	.A1(n6553), 
	.A0(\ram[110][2] ));
   AOI22X1 U10248 (.Y(n12343), 
	.B1(n6572), 
	.B0(\ram[109][2] ), 
	.A1(n6591), 
	.A0(\ram[108][2] ));
   AOI22X1 U10249 (.Y(n12342), 
	.B1(n6610), 
	.B0(\ram[107][2] ), 
	.A1(n6629), 
	.A0(\ram[106][2] ));
   OAI21XL U10250 (.Y(n12312), 
	.B0(n9718), 
	.A1(n12347), 
	.A0(n12346));
   NAND4X1 U10251 (.Y(n12347), 
	.D(n12351), 
	.C(n12350), 
	.B(n12349), 
	.A(n12348));
   AOI22X1 U10252 (.Y(n12351), 
	.B1(n6342), 
	.B0(\ram[89][2] ), 
	.A1(n6362), 
	.A0(\ram[88][2] ));
   AOI22X1 U10253 (.Y(n12350), 
	.B1(n6381), 
	.B0(\ram[87][2] ), 
	.A1(n6400), 
	.A0(\ram[86][2] ));
   AOI22X1 U10254 (.Y(n12349), 
	.B1(n6419), 
	.B0(\ram[85][2] ), 
	.A1(n6438), 
	.A0(\ram[84][2] ));
   AOI22X1 U10255 (.Y(n12348), 
	.B1(n6457), 
	.B0(\ram[83][2] ), 
	.A1(n6476), 
	.A0(\ram[82][2] ));
   NAND4X1 U10256 (.Y(n12346), 
	.D(n12355), 
	.C(n12354), 
	.B(n12353), 
	.A(n12352));
   AOI22X1 U10257 (.Y(n12355), 
	.B1(n6495), 
	.B0(\ram[81][2] ), 
	.A1(n6514), 
	.A0(\ram[80][2] ));
   AOI22X1 U10258 (.Y(n12354), 
	.B1(n6533), 
	.B0(\ram[95][2] ), 
	.A1(n6553), 
	.A0(\ram[94][2] ));
   AOI22X1 U10259 (.Y(n12353), 
	.B1(n6572), 
	.B0(\ram[93][2] ), 
	.A1(n6591), 
	.A0(\ram[92][2] ));
   AOI22X1 U10260 (.Y(n12352), 
	.B1(n6610), 
	.B0(\ram[91][2] ), 
	.A1(n6629), 
	.A0(\ram[90][2] ));
   NAND4X1 U10261 (.Y(n12220), 
	.D(n12359), 
	.C(n12358), 
	.B(n12357), 
	.A(n12356));
   OAI21XL U10262 (.Y(n12359), 
	.B0(n10007), 
	.A1(n12361), 
	.A0(n12360));
   NAND4X1 U10263 (.Y(n12361), 
	.D(n12365), 
	.C(n12364), 
	.B(n12363), 
	.A(n12362));
   AOI22X1 U10264 (.Y(n12365), 
	.B1(n6342), 
	.B0(\ram[73][2] ), 
	.A1(n6362), 
	.A0(\ram[72][2] ));
   AOI22X1 U10265 (.Y(n12364), 
	.B1(n6381), 
	.B0(\ram[71][2] ), 
	.A1(n6400), 
	.A0(\ram[70][2] ));
   AOI22X1 U10266 (.Y(n12363), 
	.B1(n6419), 
	.B0(\ram[69][2] ), 
	.A1(n6438), 
	.A0(\ram[68][2] ));
   AOI22X1 U10267 (.Y(n12362), 
	.B1(n6457), 
	.B0(\ram[67][2] ), 
	.A1(n6476), 
	.A0(\ram[66][2] ));
   NAND4X1 U10268 (.Y(n12360), 
	.D(n12369), 
	.C(n12368), 
	.B(n12367), 
	.A(n12366));
   AOI22X1 U10269 (.Y(n12369), 
	.B1(n6495), 
	.B0(\ram[65][2] ), 
	.A1(n6514), 
	.A0(\ram[64][2] ));
   AOI22X1 U10270 (.Y(n12368), 
	.B1(n6533), 
	.B0(\ram[79][2] ), 
	.A1(n6553), 
	.A0(\ram[78][2] ));
   AOI22X1 U10271 (.Y(n12367), 
	.B1(n6572), 
	.B0(\ram[77][2] ), 
	.A1(n6591), 
	.A0(\ram[76][2] ));
   AOI22X1 U10272 (.Y(n12366), 
	.B1(n6610), 
	.B0(\ram[75][2] ), 
	.A1(n6629), 
	.A0(\ram[74][2] ));
   OAI21XL U10273 (.Y(n12358), 
	.B0(n10296), 
	.A1(n12371), 
	.A0(n12370));
   NAND4X1 U10274 (.Y(n12371), 
	.D(n12375), 
	.C(n12374), 
	.B(n12373), 
	.A(n12372));
   AOI22X1 U10275 (.Y(n12375), 
	.B1(n6342), 
	.B0(\ram[57][2] ), 
	.A1(n6362), 
	.A0(\ram[56][2] ));
   AOI22X1 U10276 (.Y(n12374), 
	.B1(n6381), 
	.B0(\ram[55][2] ), 
	.A1(n6400), 
	.A0(\ram[54][2] ));
   AOI22X1 U10277 (.Y(n12373), 
	.B1(n6419), 
	.B0(\ram[53][2] ), 
	.A1(n6438), 
	.A0(\ram[52][2] ));
   AOI22X1 U10278 (.Y(n12372), 
	.B1(n6457), 
	.B0(\ram[51][2] ), 
	.A1(n6476), 
	.A0(\ram[50][2] ));
   NAND4X1 U10279 (.Y(n12370), 
	.D(n12379), 
	.C(n12378), 
	.B(n12377), 
	.A(n12376));
   AOI22X1 U10280 (.Y(n12379), 
	.B1(n6495), 
	.B0(\ram[49][2] ), 
	.A1(n6514), 
	.A0(\ram[48][2] ));
   AOI22X1 U10281 (.Y(n12378), 
	.B1(n6533), 
	.B0(\ram[63][2] ), 
	.A1(n6553), 
	.A0(\ram[62][2] ));
   AOI22X1 U10282 (.Y(n12377), 
	.B1(n6572), 
	.B0(\ram[61][2] ), 
	.A1(n6591), 
	.A0(\ram[60][2] ));
   AOI22X1 U10283 (.Y(n12376), 
	.B1(n6610), 
	.B0(\ram[59][2] ), 
	.A1(n6629), 
	.A0(\ram[58][2] ));
   OAI21XL U10284 (.Y(n12357), 
	.B0(n10585), 
	.A1(n12381), 
	.A0(n12380));
   NAND4X1 U10285 (.Y(n12381), 
	.D(n12385), 
	.C(n12384), 
	.B(n12383), 
	.A(n12382));
   AOI22X1 U10286 (.Y(n12385), 
	.B1(n6342), 
	.B0(\ram[41][2] ), 
	.A1(n6362), 
	.A0(\ram[40][2] ));
   AOI22X1 U10287 (.Y(n12384), 
	.B1(n6381), 
	.B0(\ram[39][2] ), 
	.A1(n6400), 
	.A0(\ram[38][2] ));
   AOI22X1 U10288 (.Y(n12383), 
	.B1(n6419), 
	.B0(\ram[37][2] ), 
	.A1(n6438), 
	.A0(\ram[36][2] ));
   AOI22X1 U10289 (.Y(n12382), 
	.B1(n6457), 
	.B0(\ram[35][2] ), 
	.A1(n6476), 
	.A0(\ram[34][2] ));
   NAND4X1 U10290 (.Y(n12380), 
	.D(n12389), 
	.C(n12388), 
	.B(n12387), 
	.A(n12386));
   AOI22X1 U10291 (.Y(n12389), 
	.B1(n6495), 
	.B0(\ram[33][2] ), 
	.A1(n6514), 
	.A0(\ram[32][2] ));
   AOI22X1 U10292 (.Y(n12388), 
	.B1(n6533), 
	.B0(\ram[47][2] ), 
	.A1(n6553), 
	.A0(\ram[46][2] ));
   AOI22X1 U10293 (.Y(n12387), 
	.B1(n6572), 
	.B0(\ram[45][2] ), 
	.A1(n6591), 
	.A0(\ram[44][2] ));
   AOI22X1 U10294 (.Y(n12386), 
	.B1(n6610), 
	.B0(\ram[43][2] ), 
	.A1(n6629), 
	.A0(\ram[42][2] ));
   OAI21XL U10295 (.Y(n12356), 
	.B0(n6343), 
	.A1(n12391), 
	.A0(n12390));
   NAND4X1 U10296 (.Y(n12391), 
	.D(n12395), 
	.C(n12394), 
	.B(n12393), 
	.A(n12392));
   AOI22X1 U10297 (.Y(n12395), 
	.B1(n6342), 
	.B0(\ram[25][2] ), 
	.A1(n6362), 
	.A0(\ram[24][2] ));
   AOI22X1 U10298 (.Y(n12394), 
	.B1(n6381), 
	.B0(\ram[23][2] ), 
	.A1(n6400), 
	.A0(\ram[22][2] ));
   AOI22X1 U10299 (.Y(n12393), 
	.B1(n6419), 
	.B0(\ram[21][2] ), 
	.A1(n6438), 
	.A0(\ram[20][2] ));
   AOI22X1 U10300 (.Y(n12392), 
	.B1(n6457), 
	.B0(\ram[19][2] ), 
	.A1(n6476), 
	.A0(\ram[18][2] ));
   NAND4X1 U10301 (.Y(n12390), 
	.D(n12399), 
	.C(n12398), 
	.B(n12397), 
	.A(n12396));
   AOI22X1 U10302 (.Y(n12399), 
	.B1(n6495), 
	.B0(\ram[17][2] ), 
	.A1(n6514), 
	.A0(\ram[16][2] ));
   AOI22X1 U10303 (.Y(n12398), 
	.B1(n6533), 
	.B0(\ram[31][2] ), 
	.A1(n6553), 
	.A0(\ram[30][2] ));
   AOI22X1 U10304 (.Y(n12397), 
	.B1(n6572), 
	.B0(\ram[29][2] ), 
	.A1(n6591), 
	.A0(\ram[28][2] ));
   AOI22X1 U10305 (.Y(n12396), 
	.B1(n6610), 
	.B0(\ram[27][2] ), 
	.A1(n6629), 
	.A0(\ram[26][2] ));
   OR4X1 U10306 (.Y(mem_read_data[1]), 
	.D(n12403), 
	.C(n12402), 
	.B(n12401), 
	.A(n12400));
   NAND4X1 U10307 (.Y(n12403), 
	.D(n12407), 
	.C(n12406), 
	.B(n12405), 
	.A(n12404));
   OAI21XL U10308 (.Y(n12407), 
	.B0(n6534), 
	.A1(n12409), 
	.A0(n12408));
   NAND4X1 U10309 (.Y(n12409), 
	.D(n12413), 
	.C(n12412), 
	.B(n12411), 
	.A(n12410));
   AOI22X1 U10310 (.Y(n12413), 
	.B1(n6342), 
	.B0(\ram[9][1] ), 
	.A1(n6362), 
	.A0(\ram[8][1] ));
   AOI22X1 U10311 (.Y(n12412), 
	.B1(n6381), 
	.B0(\ram[7][1] ), 
	.A1(n6400), 
	.A0(\ram[6][1] ));
   AOI22X1 U10312 (.Y(n12411), 
	.B1(n6419), 
	.B0(\ram[5][1] ), 
	.A1(n6438), 
	.A0(\ram[4][1] ));
   AOI22X1 U10313 (.Y(n12410), 
	.B1(n6457), 
	.B0(\ram[3][1] ), 
	.A1(n6476), 
	.A0(\ram[2][1] ));
   NAND4X1 U10314 (.Y(n12408), 
	.D(n12417), 
	.C(n12416), 
	.B(n12415), 
	.A(n12414));
   AOI22X1 U10315 (.Y(n12417), 
	.B1(n6495), 
	.B0(\ram[1][1] ), 
	.A1(n6514), 
	.A0(\ram[0][1] ));
   AOI22X1 U10316 (.Y(n12416), 
	.B1(n6533), 
	.B0(\ram[15][1] ), 
	.A1(n6553), 
	.A0(\ram[14][1] ));
   AOI22X1 U10317 (.Y(n12415), 
	.B1(n6572), 
	.B0(\ram[13][1] ), 
	.A1(n6591), 
	.A0(\ram[12][1] ));
   AOI22X1 U10318 (.Y(n12414), 
	.B1(n6610), 
	.B0(\ram[11][1] ), 
	.A1(n6629), 
	.A0(\ram[10][1] ));
   OAI21XL U10319 (.Y(n12406), 
	.B0(n6828), 
	.A1(n12419), 
	.A0(n12418));
   NAND4X1 U10320 (.Y(n12419), 
	.D(n12423), 
	.C(n12422), 
	.B(n12421), 
	.A(n12420));
   AOI22X1 U10321 (.Y(n12423), 
	.B1(n6342), 
	.B0(\ram[249][1] ), 
	.A1(n6362), 
	.A0(\ram[248][1] ));
   AOI22X1 U10322 (.Y(n12422), 
	.B1(n6381), 
	.B0(\ram[247][1] ), 
	.A1(n6400), 
	.A0(\ram[246][1] ));
   AOI22X1 U10323 (.Y(n12421), 
	.B1(n6419), 
	.B0(\ram[245][1] ), 
	.A1(n6438), 
	.A0(\ram[244][1] ));
   AOI22X1 U10324 (.Y(n12420), 
	.B1(n6457), 
	.B0(\ram[243][1] ), 
	.A1(n6476), 
	.A0(\ram[242][1] ));
   NAND4X1 U10325 (.Y(n12418), 
	.D(n12427), 
	.C(n12426), 
	.B(n12425), 
	.A(n12424));
   AOI22X1 U10326 (.Y(n12427), 
	.B1(n6495), 
	.B0(\ram[241][1] ), 
	.A1(n6514), 
	.A0(\ram[240][1] ));
   AOI22X1 U10327 (.Y(n12426), 
	.B1(n6533), 
	.B0(\ram[255][1] ), 
	.A1(n6553), 
	.A0(\ram[254][1] ));
   AOI22X1 U10328 (.Y(n12425), 
	.B1(n6572), 
	.B0(\ram[253][1] ), 
	.A1(n6591), 
	.A0(\ram[252][1] ));
   AOI22X1 U10329 (.Y(n12424), 
	.B1(n6610), 
	.B0(\ram[251][1] ), 
	.A1(n6629), 
	.A0(\ram[250][1] ));
   OAI21XL U10330 (.Y(n12405), 
	.B0(n7117), 
	.A1(n12429), 
	.A0(n12428));
   NAND4X1 U10331 (.Y(n12429), 
	.D(n12433), 
	.C(n12432), 
	.B(n12431), 
	.A(n12430));
   AOI22X1 U10332 (.Y(n12433), 
	.B1(n6342), 
	.B0(\ram[233][1] ), 
	.A1(n6362), 
	.A0(\ram[232][1] ));
   AOI22X1 U10333 (.Y(n12432), 
	.B1(n6381), 
	.B0(\ram[231][1] ), 
	.A1(n6400), 
	.A0(\ram[230][1] ));
   AOI22X1 U10334 (.Y(n12431), 
	.B1(n6419), 
	.B0(\ram[229][1] ), 
	.A1(n6438), 
	.A0(\ram[228][1] ));
   AOI22X1 U10335 (.Y(n12430), 
	.B1(n6457), 
	.B0(\ram[227][1] ), 
	.A1(n6476), 
	.A0(\ram[226][1] ));
   NAND4X1 U10336 (.Y(n12428), 
	.D(n12437), 
	.C(n12436), 
	.B(n12435), 
	.A(n12434));
   AOI22X1 U10337 (.Y(n12437), 
	.B1(n6495), 
	.B0(\ram[225][1] ), 
	.A1(n6514), 
	.A0(\ram[224][1] ));
   AOI22X1 U10338 (.Y(n12436), 
	.B1(n6533), 
	.B0(\ram[239][1] ), 
	.A1(n6553), 
	.A0(\ram[238][1] ));
   AOI22X1 U10339 (.Y(n12435), 
	.B1(n6572), 
	.B0(\ram[237][1] ), 
	.A1(n6591), 
	.A0(\ram[236][1] ));
   AOI22X1 U10340 (.Y(n12434), 
	.B1(n6610), 
	.B0(\ram[235][1] ), 
	.A1(n6629), 
	.A0(\ram[234][1] ));
   OAI21XL U10341 (.Y(n12404), 
	.B0(n7406), 
	.A1(n12439), 
	.A0(n12438));
   NAND4X1 U10342 (.Y(n12439), 
	.D(n12443), 
	.C(n12442), 
	.B(n12441), 
	.A(n12440));
   AOI22X1 U10343 (.Y(n12443), 
	.B1(n6342), 
	.B0(\ram[217][1] ), 
	.A1(n6362), 
	.A0(\ram[216][1] ));
   AOI22X1 U10344 (.Y(n12442), 
	.B1(n6381), 
	.B0(\ram[215][1] ), 
	.A1(n6400), 
	.A0(\ram[214][1] ));
   AOI22X1 U10345 (.Y(n12441), 
	.B1(n6419), 
	.B0(\ram[213][1] ), 
	.A1(n6438), 
	.A0(\ram[212][1] ));
   AOI22X1 U10346 (.Y(n12440), 
	.B1(n6457), 
	.B0(\ram[211][1] ), 
	.A1(n6476), 
	.A0(\ram[210][1] ));
   NAND4X1 U10347 (.Y(n12438), 
	.D(n12447), 
	.C(n12446), 
	.B(n12445), 
	.A(n12444));
   AOI22X1 U10348 (.Y(n12447), 
	.B1(n6495), 
	.B0(\ram[209][1] ), 
	.A1(n6514), 
	.A0(\ram[208][1] ));
   AOI22X1 U10349 (.Y(n12446), 
	.B1(n6533), 
	.B0(\ram[223][1] ), 
	.A1(n6553), 
	.A0(\ram[222][1] ));
   AOI22X1 U10350 (.Y(n12445), 
	.B1(n6572), 
	.B0(\ram[221][1] ), 
	.A1(n6591), 
	.A0(\ram[220][1] ));
   AOI22X1 U10351 (.Y(n12444), 
	.B1(n6610), 
	.B0(\ram[219][1] ), 
	.A1(n6629), 
	.A0(\ram[218][1] ));
   NAND4X1 U10352 (.Y(n12402), 
	.D(n12451), 
	.C(n12450), 
	.B(n12449), 
	.A(n12448));
   OAI21XL U10353 (.Y(n12451), 
	.B0(n7695), 
	.A1(n12453), 
	.A0(n12452));
   NAND4X1 U10354 (.Y(n12453), 
	.D(n12457), 
	.C(n12456), 
	.B(n12455), 
	.A(n12454));
   AOI22X1 U10355 (.Y(n12457), 
	.B1(n6342), 
	.B0(\ram[201][1] ), 
	.A1(n6362), 
	.A0(\ram[200][1] ));
   AOI22X1 U10356 (.Y(n12456), 
	.B1(n6381), 
	.B0(\ram[199][1] ), 
	.A1(n6400), 
	.A0(\ram[198][1] ));
   AOI22X1 U10357 (.Y(n12455), 
	.B1(n6419), 
	.B0(\ram[197][1] ), 
	.A1(n6438), 
	.A0(\ram[196][1] ));
   AOI22X1 U10358 (.Y(n12454), 
	.B1(n6457), 
	.B0(\ram[195][1] ), 
	.A1(n6476), 
	.A0(\ram[194][1] ));
   NAND4X1 U10359 (.Y(n12452), 
	.D(n12461), 
	.C(n12460), 
	.B(n12459), 
	.A(n12458));
   AOI22X1 U10360 (.Y(n12461), 
	.B1(n6495), 
	.B0(\ram[193][1] ), 
	.A1(n6514), 
	.A0(\ram[192][1] ));
   AOI22X1 U10361 (.Y(n12460), 
	.B1(n6533), 
	.B0(\ram[207][1] ), 
	.A1(n6553), 
	.A0(\ram[206][1] ));
   AOI22X1 U10362 (.Y(n12459), 
	.B1(n6572), 
	.B0(\ram[205][1] ), 
	.A1(n6591), 
	.A0(\ram[204][1] ));
   AOI22X1 U10363 (.Y(n12458), 
	.B1(n6610), 
	.B0(\ram[203][1] ), 
	.A1(n6629), 
	.A0(\ram[202][1] ));
   OAI21XL U10364 (.Y(n12450), 
	.B0(n7984), 
	.A1(n12463), 
	.A0(n12462));
   NAND4X1 U10365 (.Y(n12463), 
	.D(n12467), 
	.C(n12466), 
	.B(n12465), 
	.A(n12464));
   AOI22X1 U10366 (.Y(n12467), 
	.B1(n6342), 
	.B0(\ram[185][1] ), 
	.A1(n6362), 
	.A0(\ram[184][1] ));
   AOI22X1 U10367 (.Y(n12466), 
	.B1(n6381), 
	.B0(\ram[183][1] ), 
	.A1(n6400), 
	.A0(\ram[182][1] ));
   AOI22X1 U10368 (.Y(n12465), 
	.B1(n6419), 
	.B0(\ram[181][1] ), 
	.A1(n6438), 
	.A0(\ram[180][1] ));
   AOI22X1 U10369 (.Y(n12464), 
	.B1(n6457), 
	.B0(\ram[179][1] ), 
	.A1(n6476), 
	.A0(\ram[178][1] ));
   NAND4X1 U10370 (.Y(n12462), 
	.D(n12471), 
	.C(n12470), 
	.B(n12469), 
	.A(n12468));
   AOI22X1 U10371 (.Y(n12471), 
	.B1(n6495), 
	.B0(\ram[177][1] ), 
	.A1(n6514), 
	.A0(\ram[176][1] ));
   AOI22X1 U10372 (.Y(n12470), 
	.B1(n6533), 
	.B0(\ram[191][1] ), 
	.A1(n6553), 
	.A0(\ram[190][1] ));
   AOI22X1 U10373 (.Y(n12469), 
	.B1(n6572), 
	.B0(\ram[189][1] ), 
	.A1(n6591), 
	.A0(\ram[188][1] ));
   AOI22X1 U10374 (.Y(n12468), 
	.B1(n6610), 
	.B0(\ram[187][1] ), 
	.A1(n6629), 
	.A0(\ram[186][1] ));
   OAI21XL U10375 (.Y(n12449), 
	.B0(n8273), 
	.A1(n12473), 
	.A0(n12472));
   NAND4X1 U10376 (.Y(n12473), 
	.D(n12477), 
	.C(n12476), 
	.B(n12475), 
	.A(n12474));
   AOI22X1 U10377 (.Y(n12477), 
	.B1(n6342), 
	.B0(\ram[169][1] ), 
	.A1(n6362), 
	.A0(\ram[168][1] ));
   AOI22X1 U10378 (.Y(n12476), 
	.B1(n6381), 
	.B0(\ram[167][1] ), 
	.A1(n6400), 
	.A0(\ram[166][1] ));
   AOI22X1 U10379 (.Y(n12475), 
	.B1(n6419), 
	.B0(\ram[165][1] ), 
	.A1(n6438), 
	.A0(\ram[164][1] ));
   AOI22X1 U10380 (.Y(n12474), 
	.B1(n6457), 
	.B0(\ram[163][1] ), 
	.A1(n6476), 
	.A0(\ram[162][1] ));
   NAND4X1 U10381 (.Y(n12472), 
	.D(n12481), 
	.C(n12480), 
	.B(n12479), 
	.A(n12478));
   AOI22X1 U10382 (.Y(n12481), 
	.B1(n6495), 
	.B0(\ram[161][1] ), 
	.A1(n6514), 
	.A0(\ram[160][1] ));
   AOI22X1 U10383 (.Y(n12480), 
	.B1(n6533), 
	.B0(\ram[175][1] ), 
	.A1(n6553), 
	.A0(\ram[174][1] ));
   AOI22X1 U10384 (.Y(n12479), 
	.B1(n6572), 
	.B0(\ram[173][1] ), 
	.A1(n6591), 
	.A0(\ram[172][1] ));
   AOI22X1 U10385 (.Y(n12478), 
	.B1(n6610), 
	.B0(\ram[171][1] ), 
	.A1(n6629), 
	.A0(\ram[170][1] ));
   OAI21XL U10386 (.Y(n12448), 
	.B0(n8562), 
	.A1(n12483), 
	.A0(n12482));
   NAND4X1 U10387 (.Y(n12483), 
	.D(n12487), 
	.C(n12486), 
	.B(n12485), 
	.A(n12484));
   AOI22X1 U10388 (.Y(n12487), 
	.B1(n6342), 
	.B0(\ram[153][1] ), 
	.A1(n6362), 
	.A0(\ram[152][1] ));
   AOI22X1 U10389 (.Y(n12486), 
	.B1(n6381), 
	.B0(\ram[151][1] ), 
	.A1(n6400), 
	.A0(\ram[150][1] ));
   AOI22X1 U10390 (.Y(n12485), 
	.B1(n6419), 
	.B0(\ram[149][1] ), 
	.A1(n6438), 
	.A0(\ram[148][1] ));
   AOI22X1 U10391 (.Y(n12484), 
	.B1(n6457), 
	.B0(\ram[147][1] ), 
	.A1(n6476), 
	.A0(\ram[146][1] ));
   NAND4X1 U10392 (.Y(n12482), 
	.D(n12491), 
	.C(n12490), 
	.B(n12489), 
	.A(n12488));
   AOI22X1 U10393 (.Y(n12491), 
	.B1(n6495), 
	.B0(\ram[145][1] ), 
	.A1(n6514), 
	.A0(\ram[144][1] ));
   AOI22X1 U10394 (.Y(n12490), 
	.B1(n6533), 
	.B0(\ram[159][1] ), 
	.A1(n6553), 
	.A0(\ram[158][1] ));
   AOI22X1 U10395 (.Y(n12489), 
	.B1(n6572), 
	.B0(\ram[157][1] ), 
	.A1(n6591), 
	.A0(\ram[156][1] ));
   AOI22X1 U10396 (.Y(n12488), 
	.B1(n6610), 
	.B0(\ram[155][1] ), 
	.A1(n6629), 
	.A0(\ram[154][1] ));
   NAND4X1 U10397 (.Y(n12401), 
	.D(n12495), 
	.C(n12494), 
	.B(n12493), 
	.A(n12492));
   OAI21XL U10398 (.Y(n12495), 
	.B0(n8851), 
	.A1(n12497), 
	.A0(n12496));
   NAND4X1 U10399 (.Y(n12497), 
	.D(n12501), 
	.C(n12500), 
	.B(n12499), 
	.A(n12498));
   AOI22X1 U10400 (.Y(n12501), 
	.B1(n6342), 
	.B0(\ram[137][1] ), 
	.A1(n6362), 
	.A0(\ram[136][1] ));
   AOI22X1 U10401 (.Y(n12500), 
	.B1(n6381), 
	.B0(\ram[135][1] ), 
	.A1(n6400), 
	.A0(\ram[134][1] ));
   AOI22X1 U10402 (.Y(n12499), 
	.B1(n6419), 
	.B0(\ram[133][1] ), 
	.A1(n6438), 
	.A0(\ram[132][1] ));
   AOI22X1 U10403 (.Y(n12498), 
	.B1(n6457), 
	.B0(\ram[131][1] ), 
	.A1(n6476), 
	.A0(\ram[130][1] ));
   NAND4X1 U10404 (.Y(n12496), 
	.D(n12505), 
	.C(n12504), 
	.B(n12503), 
	.A(n12502));
   AOI22X1 U10405 (.Y(n12505), 
	.B1(n6495), 
	.B0(\ram[129][1] ), 
	.A1(n6514), 
	.A0(\ram[128][1] ));
   AOI22X1 U10406 (.Y(n12504), 
	.B1(n6533), 
	.B0(\ram[143][1] ), 
	.A1(n6553), 
	.A0(\ram[142][1] ));
   AOI22X1 U10407 (.Y(n12503), 
	.B1(n6572), 
	.B0(\ram[141][1] ), 
	.A1(n6591), 
	.A0(\ram[140][1] ));
   AOI22X1 U10408 (.Y(n12502), 
	.B1(n6610), 
	.B0(\ram[139][1] ), 
	.A1(n6629), 
	.A0(\ram[138][1] ));
   OAI21XL U10409 (.Y(n12494), 
	.B0(n9140), 
	.A1(n12507), 
	.A0(n12506));
   NAND4X1 U10410 (.Y(n12507), 
	.D(n12511), 
	.C(n12510), 
	.B(n12509), 
	.A(n12508));
   AOI22X1 U10411 (.Y(n12511), 
	.B1(n6342), 
	.B0(\ram[121][1] ), 
	.A1(n6362), 
	.A0(\ram[120][1] ));
   AOI22X1 U10412 (.Y(n12510), 
	.B1(n6381), 
	.B0(\ram[119][1] ), 
	.A1(n6400), 
	.A0(\ram[118][1] ));
   AOI22X1 U10413 (.Y(n12509), 
	.B1(n6419), 
	.B0(\ram[117][1] ), 
	.A1(n6438), 
	.A0(\ram[116][1] ));
   AOI22X1 U10414 (.Y(n12508), 
	.B1(n6457), 
	.B0(\ram[115][1] ), 
	.A1(n6476), 
	.A0(\ram[114][1] ));
   NAND4X1 U10415 (.Y(n12506), 
	.D(n12515), 
	.C(n12514), 
	.B(n12513), 
	.A(n12512));
   AOI22X1 U10416 (.Y(n12515), 
	.B1(n6495), 
	.B0(\ram[113][1] ), 
	.A1(n6514), 
	.A0(\ram[112][1] ));
   AOI22X1 U10417 (.Y(n12514), 
	.B1(n6533), 
	.B0(\ram[127][1] ), 
	.A1(n6553), 
	.A0(\ram[126][1] ));
   AOI22X1 U10418 (.Y(n12513), 
	.B1(n6572), 
	.B0(\ram[125][1] ), 
	.A1(n6591), 
	.A0(\ram[124][1] ));
   AOI22X1 U10419 (.Y(n12512), 
	.B1(n6610), 
	.B0(\ram[123][1] ), 
	.A1(n6629), 
	.A0(\ram[122][1] ));
   OAI21XL U10420 (.Y(n12493), 
	.B0(n9429), 
	.A1(n12517), 
	.A0(n12516));
   NAND4X1 U10421 (.Y(n12517), 
	.D(n12521), 
	.C(n12520), 
	.B(n12519), 
	.A(n12518));
   AOI22X1 U10422 (.Y(n12521), 
	.B1(n6342), 
	.B0(\ram[105][1] ), 
	.A1(n6362), 
	.A0(\ram[104][1] ));
   AOI22X1 U10423 (.Y(n12520), 
	.B1(n6381), 
	.B0(\ram[103][1] ), 
	.A1(n6400), 
	.A0(\ram[102][1] ));
   AOI22X1 U10424 (.Y(n12519), 
	.B1(n6419), 
	.B0(\ram[101][1] ), 
	.A1(n6438), 
	.A0(\ram[100][1] ));
   AOI22X1 U10425 (.Y(n12518), 
	.B1(n6457), 
	.B0(\ram[99][1] ), 
	.A1(n6476), 
	.A0(\ram[98][1] ));
   NAND4X1 U10426 (.Y(n12516), 
	.D(n12525), 
	.C(n12524), 
	.B(n12523), 
	.A(n12522));
   AOI22X1 U10427 (.Y(n12525), 
	.B1(n6495), 
	.B0(\ram[97][1] ), 
	.A1(n6514), 
	.A0(\ram[96][1] ));
   AOI22X1 U10428 (.Y(n12524), 
	.B1(n6533), 
	.B0(\ram[111][1] ), 
	.A1(n6553), 
	.A0(\ram[110][1] ));
   AOI22X1 U10429 (.Y(n12523), 
	.B1(n6572), 
	.B0(\ram[109][1] ), 
	.A1(n6591), 
	.A0(\ram[108][1] ));
   AOI22X1 U10430 (.Y(n12522), 
	.B1(n6610), 
	.B0(\ram[107][1] ), 
	.A1(n6629), 
	.A0(\ram[106][1] ));
   OAI21XL U10431 (.Y(n12492), 
	.B0(n9718), 
	.A1(n12527), 
	.A0(n12526));
   NAND4X1 U10432 (.Y(n12527), 
	.D(n12531), 
	.C(n12530), 
	.B(n12529), 
	.A(n12528));
   AOI22X1 U10433 (.Y(n12531), 
	.B1(n6342), 
	.B0(\ram[89][1] ), 
	.A1(n6362), 
	.A0(\ram[88][1] ));
   AOI22X1 U10434 (.Y(n12530), 
	.B1(n6381), 
	.B0(\ram[87][1] ), 
	.A1(n6400), 
	.A0(\ram[86][1] ));
   AOI22X1 U10435 (.Y(n12529), 
	.B1(n6419), 
	.B0(\ram[85][1] ), 
	.A1(n6438), 
	.A0(\ram[84][1] ));
   AOI22X1 U10436 (.Y(n12528), 
	.B1(n6457), 
	.B0(\ram[83][1] ), 
	.A1(n6476), 
	.A0(\ram[82][1] ));
   NAND4X1 U10437 (.Y(n12526), 
	.D(n12535), 
	.C(n12534), 
	.B(n12533), 
	.A(n12532));
   AOI22X1 U10438 (.Y(n12535), 
	.B1(n6495), 
	.B0(\ram[81][1] ), 
	.A1(n6514), 
	.A0(\ram[80][1] ));
   AOI22X1 U10439 (.Y(n12534), 
	.B1(n6533), 
	.B0(\ram[95][1] ), 
	.A1(n6553), 
	.A0(\ram[94][1] ));
   AOI22X1 U10440 (.Y(n12533), 
	.B1(n6572), 
	.B0(\ram[93][1] ), 
	.A1(n6591), 
	.A0(\ram[92][1] ));
   AOI22X1 U10441 (.Y(n12532), 
	.B1(n6610), 
	.B0(\ram[91][1] ), 
	.A1(n6629), 
	.A0(\ram[90][1] ));
   NAND4X1 U10442 (.Y(n12400), 
	.D(n12539), 
	.C(n12538), 
	.B(n12537), 
	.A(n12536));
   OAI21XL U10443 (.Y(n12539), 
	.B0(n10007), 
	.A1(n12541), 
	.A0(n12540));
   NAND4X1 U10444 (.Y(n12541), 
	.D(n12545), 
	.C(n12544), 
	.B(n12543), 
	.A(n12542));
   AOI22X1 U10445 (.Y(n12545), 
	.B1(n6342), 
	.B0(\ram[73][1] ), 
	.A1(n6362), 
	.A0(\ram[72][1] ));
   AOI22X1 U10446 (.Y(n12544), 
	.B1(n6381), 
	.B0(\ram[71][1] ), 
	.A1(n6400), 
	.A0(\ram[70][1] ));
   AOI22X1 U10447 (.Y(n12543), 
	.B1(n6419), 
	.B0(\ram[69][1] ), 
	.A1(n6438), 
	.A0(\ram[68][1] ));
   AOI22X1 U10448 (.Y(n12542), 
	.B1(n6457), 
	.B0(\ram[67][1] ), 
	.A1(n6476), 
	.A0(\ram[66][1] ));
   NAND4X1 U10449 (.Y(n12540), 
	.D(n12549), 
	.C(n12548), 
	.B(n12547), 
	.A(n12546));
   AOI22X1 U10450 (.Y(n12549), 
	.B1(n6495), 
	.B0(\ram[65][1] ), 
	.A1(n6514), 
	.A0(\ram[64][1] ));
   AOI22X1 U10451 (.Y(n12548), 
	.B1(n6533), 
	.B0(\ram[79][1] ), 
	.A1(n6553), 
	.A0(\ram[78][1] ));
   AOI22X1 U10452 (.Y(n12547), 
	.B1(n6572), 
	.B0(\ram[77][1] ), 
	.A1(n6591), 
	.A0(\ram[76][1] ));
   AOI22X1 U10453 (.Y(n12546), 
	.B1(n6610), 
	.B0(\ram[75][1] ), 
	.A1(n6629), 
	.A0(\ram[74][1] ));
   OAI21XL U10454 (.Y(n12538), 
	.B0(n10296), 
	.A1(n12551), 
	.A0(n12550));
   NAND4X1 U10455 (.Y(n12551), 
	.D(n12555), 
	.C(n12554), 
	.B(n12553), 
	.A(n12552));
   AOI22X1 U10456 (.Y(n12555), 
	.B1(n6342), 
	.B0(\ram[57][1] ), 
	.A1(n6362), 
	.A0(\ram[56][1] ));
   AOI22X1 U10457 (.Y(n12554), 
	.B1(n6381), 
	.B0(\ram[55][1] ), 
	.A1(n6400), 
	.A0(\ram[54][1] ));
   AOI22X1 U10458 (.Y(n12553), 
	.B1(n6419), 
	.B0(\ram[53][1] ), 
	.A1(n6438), 
	.A0(\ram[52][1] ));
   AOI22X1 U10459 (.Y(n12552), 
	.B1(n6457), 
	.B0(\ram[51][1] ), 
	.A1(n6476), 
	.A0(\ram[50][1] ));
   NAND4X1 U10460 (.Y(n12550), 
	.D(n12559), 
	.C(n12558), 
	.B(n12557), 
	.A(n12556));
   AOI22X1 U10461 (.Y(n12559), 
	.B1(n6495), 
	.B0(\ram[49][1] ), 
	.A1(n6514), 
	.A0(\ram[48][1] ));
   AOI22X1 U10462 (.Y(n12558), 
	.B1(n6533), 
	.B0(\ram[63][1] ), 
	.A1(n6553), 
	.A0(\ram[62][1] ));
   AOI22X1 U10463 (.Y(n12557), 
	.B1(n6572), 
	.B0(\ram[61][1] ), 
	.A1(n6591), 
	.A0(\ram[60][1] ));
   AOI22X1 U10464 (.Y(n12556), 
	.B1(n6610), 
	.B0(\ram[59][1] ), 
	.A1(n6629), 
	.A0(\ram[58][1] ));
   OAI21XL U10465 (.Y(n12537), 
	.B0(n10585), 
	.A1(n12561), 
	.A0(n12560));
   NAND4X1 U10466 (.Y(n12561), 
	.D(n12565), 
	.C(n12564), 
	.B(n12563), 
	.A(n12562));
   AOI22X1 U10467 (.Y(n12565), 
	.B1(n6342), 
	.B0(\ram[41][1] ), 
	.A1(n6362), 
	.A0(\ram[40][1] ));
   AOI22X1 U10468 (.Y(n12564), 
	.B1(n6381), 
	.B0(\ram[39][1] ), 
	.A1(n6400), 
	.A0(\ram[38][1] ));
   AOI22X1 U10469 (.Y(n12563), 
	.B1(n6419), 
	.B0(\ram[37][1] ), 
	.A1(n6438), 
	.A0(\ram[36][1] ));
   AOI22X1 U10470 (.Y(n12562), 
	.B1(n6457), 
	.B0(\ram[35][1] ), 
	.A1(n6476), 
	.A0(\ram[34][1] ));
   NAND4X1 U10471 (.Y(n12560), 
	.D(n12569), 
	.C(n12568), 
	.B(n12567), 
	.A(n12566));
   AOI22X1 U10472 (.Y(n12569), 
	.B1(n6495), 
	.B0(\ram[33][1] ), 
	.A1(n6514), 
	.A0(\ram[32][1] ));
   AOI22X1 U10473 (.Y(n12568), 
	.B1(n6533), 
	.B0(\ram[47][1] ), 
	.A1(n6553), 
	.A0(\ram[46][1] ));
   AOI22X1 U10474 (.Y(n12567), 
	.B1(n6572), 
	.B0(\ram[45][1] ), 
	.A1(n6591), 
	.A0(\ram[44][1] ));
   AOI22X1 U10475 (.Y(n12566), 
	.B1(n6610), 
	.B0(\ram[43][1] ), 
	.A1(n6629), 
	.A0(\ram[42][1] ));
   OAI21XL U10476 (.Y(n12536), 
	.B0(n6343), 
	.A1(n12571), 
	.A0(n12570));
   NAND4X1 U10477 (.Y(n12571), 
	.D(n12575), 
	.C(n12574), 
	.B(n12573), 
	.A(n12572));
   AOI22X1 U10478 (.Y(n12575), 
	.B1(n6342), 
	.B0(\ram[25][1] ), 
	.A1(n6362), 
	.A0(\ram[24][1] ));
   AOI22X1 U10479 (.Y(n12574), 
	.B1(n6381), 
	.B0(\ram[23][1] ), 
	.A1(n6400), 
	.A0(\ram[22][1] ));
   AOI22X1 U10480 (.Y(n12573), 
	.B1(n6419), 
	.B0(\ram[21][1] ), 
	.A1(n6438), 
	.A0(\ram[20][1] ));
   AOI22X1 U10481 (.Y(n12572), 
	.B1(n6457), 
	.B0(\ram[19][1] ), 
	.A1(n6476), 
	.A0(\ram[18][1] ));
   NAND4X1 U10482 (.Y(n12570), 
	.D(n12579), 
	.C(n12578), 
	.B(n12577), 
	.A(n12576));
   AOI22X1 U10483 (.Y(n12579), 
	.B1(n6495), 
	.B0(\ram[17][1] ), 
	.A1(n6514), 
	.A0(\ram[16][1] ));
   AOI22X1 U10484 (.Y(n12578), 
	.B1(n6533), 
	.B0(\ram[31][1] ), 
	.A1(n6553), 
	.A0(\ram[30][1] ));
   AOI22X1 U10485 (.Y(n12577), 
	.B1(n6572), 
	.B0(\ram[29][1] ), 
	.A1(n6591), 
	.A0(\ram[28][1] ));
   AOI22X1 U10486 (.Y(n12576), 
	.B1(n6610), 
	.B0(\ram[27][1] ), 
	.A1(n6629), 
	.A0(\ram[26][1] ));
   OR4X1 U10487 (.Y(mem_read_data[15]), 
	.D(n12583), 
	.C(n12582), 
	.B(n12581), 
	.A(n12580));
   NAND4X1 U10488 (.Y(n12583), 
	.D(n12587), 
	.C(n12586), 
	.B(n12585), 
	.A(n12584));
   OAI21XL U10489 (.Y(n12587), 
	.B0(n6534), 
	.A1(n12589), 
	.A0(n12588));
   NAND4X1 U10490 (.Y(n12589), 
	.D(n12593), 
	.C(n12592), 
	.B(n12591), 
	.A(n12590));
   AOI22X1 U10491 (.Y(n12593), 
	.B1(n6342), 
	.B0(\ram[9][15] ), 
	.A1(n6362), 
	.A0(\ram[8][15] ));
   AOI22X1 U10492 (.Y(n12592), 
	.B1(n6381), 
	.B0(\ram[7][15] ), 
	.A1(n6400), 
	.A0(\ram[6][15] ));
   AOI22X1 U10493 (.Y(n12591), 
	.B1(n6419), 
	.B0(\ram[5][15] ), 
	.A1(n6438), 
	.A0(\ram[4][15] ));
   AOI22X1 U10494 (.Y(n12590), 
	.B1(n6457), 
	.B0(\ram[3][15] ), 
	.A1(n6476), 
	.A0(\ram[2][15] ));
   NAND4X1 U10495 (.Y(n12588), 
	.D(n12597), 
	.C(n12596), 
	.B(n12595), 
	.A(n12594));
   AOI22X1 U10496 (.Y(n12597), 
	.B1(n6495), 
	.B0(\ram[1][15] ), 
	.A1(n6514), 
	.A0(\ram[0][15] ));
   AOI22X1 U10497 (.Y(n12596), 
	.B1(n6533), 
	.B0(\ram[15][15] ), 
	.A1(n6553), 
	.A0(\ram[14][15] ));
   AOI22X1 U10498 (.Y(n12595), 
	.B1(n6572), 
	.B0(\ram[13][15] ), 
	.A1(n6591), 
	.A0(\ram[12][15] ));
   AOI22X1 U10499 (.Y(n12594), 
	.B1(n6610), 
	.B0(\ram[11][15] ), 
	.A1(n6629), 
	.A0(\ram[10][15] ));
   OAI21XL U10500 (.Y(n12586), 
	.B0(n6828), 
	.A1(n12599), 
	.A0(n12598));
   NAND4X1 U10501 (.Y(n12599), 
	.D(n12603), 
	.C(n12602), 
	.B(n12601), 
	.A(n12600));
   AOI22X1 U10502 (.Y(n12603), 
	.B1(n6342), 
	.B0(\ram[249][15] ), 
	.A1(n6362), 
	.A0(\ram[248][15] ));
   AOI22X1 U10503 (.Y(n12602), 
	.B1(n6381), 
	.B0(\ram[247][15] ), 
	.A1(n6400), 
	.A0(\ram[246][15] ));
   AOI22X1 U10504 (.Y(n12601), 
	.B1(n6419), 
	.B0(\ram[245][15] ), 
	.A1(n6438), 
	.A0(\ram[244][15] ));
   AOI22X1 U10505 (.Y(n12600), 
	.B1(n6457), 
	.B0(\ram[243][15] ), 
	.A1(n6476), 
	.A0(\ram[242][15] ));
   NAND4X1 U10506 (.Y(n12598), 
	.D(n12607), 
	.C(n12606), 
	.B(n12605), 
	.A(n12604));
   AOI22X1 U10507 (.Y(n12607), 
	.B1(n6495), 
	.B0(\ram[241][15] ), 
	.A1(n6514), 
	.A0(\ram[240][15] ));
   AOI22X1 U10508 (.Y(n12606), 
	.B1(n6533), 
	.B0(\ram[255][15] ), 
	.A1(n6553), 
	.A0(\ram[254][15] ));
   AOI22X1 U10509 (.Y(n12605), 
	.B1(n6572), 
	.B0(\ram[253][15] ), 
	.A1(n6591), 
	.A0(\ram[252][15] ));
   AOI22X1 U10510 (.Y(n12604), 
	.B1(n6610), 
	.B0(\ram[251][15] ), 
	.A1(n6629), 
	.A0(\ram[250][15] ));
   OAI21XL U10511 (.Y(n12585), 
	.B0(n7117), 
	.A1(n12609), 
	.A0(n12608));
   NAND4X1 U10512 (.Y(n12609), 
	.D(n12613), 
	.C(n12612), 
	.B(n12611), 
	.A(n12610));
   AOI22X1 U10513 (.Y(n12613), 
	.B1(n6342), 
	.B0(\ram[233][15] ), 
	.A1(n6362), 
	.A0(\ram[232][15] ));
   AOI22X1 U10514 (.Y(n12612), 
	.B1(n6381), 
	.B0(\ram[231][15] ), 
	.A1(n6400), 
	.A0(\ram[230][15] ));
   AOI22X1 U10515 (.Y(n12611), 
	.B1(n6419), 
	.B0(\ram[229][15] ), 
	.A1(n6438), 
	.A0(\ram[228][15] ));
   AOI22X1 U10516 (.Y(n12610), 
	.B1(n6457), 
	.B0(\ram[227][15] ), 
	.A1(n6476), 
	.A0(\ram[226][15] ));
   NAND4X1 U10517 (.Y(n12608), 
	.D(n12617), 
	.C(n12616), 
	.B(n12615), 
	.A(n12614));
   AOI22X1 U10518 (.Y(n12617), 
	.B1(n6495), 
	.B0(\ram[225][15] ), 
	.A1(n6514), 
	.A0(\ram[224][15] ));
   AOI22X1 U10519 (.Y(n12616), 
	.B1(n6533), 
	.B0(\ram[239][15] ), 
	.A1(n6553), 
	.A0(\ram[238][15] ));
   AOI22X1 U10520 (.Y(n12615), 
	.B1(n6572), 
	.B0(\ram[237][15] ), 
	.A1(n6591), 
	.A0(\ram[236][15] ));
   AOI22X1 U10521 (.Y(n12614), 
	.B1(n6610), 
	.B0(\ram[235][15] ), 
	.A1(n6629), 
	.A0(\ram[234][15] ));
   OAI21XL U10522 (.Y(n12584), 
	.B0(n7406), 
	.A1(n12619), 
	.A0(n12618));
   NAND4X1 U10523 (.Y(n12619), 
	.D(n12623), 
	.C(n12622), 
	.B(n12621), 
	.A(n12620));
   AOI22X1 U10524 (.Y(n12623), 
	.B1(n6342), 
	.B0(\ram[217][15] ), 
	.A1(n6362), 
	.A0(\ram[216][15] ));
   AOI22X1 U10525 (.Y(n12622), 
	.B1(n6381), 
	.B0(\ram[215][15] ), 
	.A1(n6400), 
	.A0(\ram[214][15] ));
   AOI22X1 U10526 (.Y(n12621), 
	.B1(n6419), 
	.B0(\ram[213][15] ), 
	.A1(n6438), 
	.A0(\ram[212][15] ));
   AOI22X1 U10527 (.Y(n12620), 
	.B1(n6457), 
	.B0(\ram[211][15] ), 
	.A1(n6476), 
	.A0(\ram[210][15] ));
   NAND4X1 U10528 (.Y(n12618), 
	.D(n12627), 
	.C(n12626), 
	.B(n12625), 
	.A(n12624));
   AOI22X1 U10529 (.Y(n12627), 
	.B1(n6495), 
	.B0(\ram[209][15] ), 
	.A1(n6514), 
	.A0(\ram[208][15] ));
   AOI22X1 U10530 (.Y(n12626), 
	.B1(n6533), 
	.B0(\ram[223][15] ), 
	.A1(n6553), 
	.A0(\ram[222][15] ));
   AOI22X1 U10531 (.Y(n12625), 
	.B1(n6572), 
	.B0(\ram[221][15] ), 
	.A1(n6591), 
	.A0(\ram[220][15] ));
   AOI22X1 U10532 (.Y(n12624), 
	.B1(n6610), 
	.B0(\ram[219][15] ), 
	.A1(n6629), 
	.A0(\ram[218][15] ));
   NAND4X1 U10533 (.Y(n12582), 
	.D(n12631), 
	.C(n12630), 
	.B(n12629), 
	.A(n12628));
   OAI21XL U10534 (.Y(n12631), 
	.B0(n7695), 
	.A1(n12633), 
	.A0(n12632));
   NAND4X1 U10535 (.Y(n12633), 
	.D(n12637), 
	.C(n12636), 
	.B(n12635), 
	.A(n12634));
   AOI22X1 U10536 (.Y(n12637), 
	.B1(n6342), 
	.B0(\ram[201][15] ), 
	.A1(n6362), 
	.A0(\ram[200][15] ));
   AOI22X1 U10537 (.Y(n12636), 
	.B1(n6381), 
	.B0(\ram[199][15] ), 
	.A1(n6400), 
	.A0(\ram[198][15] ));
   AOI22X1 U10538 (.Y(n12635), 
	.B1(n6419), 
	.B0(\ram[197][15] ), 
	.A1(n6438), 
	.A0(\ram[196][15] ));
   AOI22X1 U10539 (.Y(n12634), 
	.B1(n6457), 
	.B0(\ram[195][15] ), 
	.A1(n6476), 
	.A0(\ram[194][15] ));
   NAND4X1 U10540 (.Y(n12632), 
	.D(n12641), 
	.C(n12640), 
	.B(n12639), 
	.A(n12638));
   AOI22X1 U10541 (.Y(n12641), 
	.B1(n6495), 
	.B0(\ram[193][15] ), 
	.A1(n6514), 
	.A0(\ram[192][15] ));
   AOI22X1 U10542 (.Y(n12640), 
	.B1(n6533), 
	.B0(\ram[207][15] ), 
	.A1(n6553), 
	.A0(\ram[206][15] ));
   AOI22X1 U10543 (.Y(n12639), 
	.B1(n6572), 
	.B0(\ram[205][15] ), 
	.A1(n6591), 
	.A0(\ram[204][15] ));
   AOI22X1 U10544 (.Y(n12638), 
	.B1(n6610), 
	.B0(\ram[203][15] ), 
	.A1(n6629), 
	.A0(\ram[202][15] ));
   OAI21XL U10545 (.Y(n12630), 
	.B0(n7984), 
	.A1(n12643), 
	.A0(n12642));
   NAND4X1 U10546 (.Y(n12643), 
	.D(n12647), 
	.C(n12646), 
	.B(n12645), 
	.A(n12644));
   AOI22X1 U10547 (.Y(n12647), 
	.B1(n6342), 
	.B0(\ram[185][15] ), 
	.A1(n6362), 
	.A0(\ram[184][15] ));
   AOI22X1 U10548 (.Y(n12646), 
	.B1(n6381), 
	.B0(\ram[183][15] ), 
	.A1(n6400), 
	.A0(\ram[182][15] ));
   AOI22X1 U10549 (.Y(n12645), 
	.B1(n6419), 
	.B0(\ram[181][15] ), 
	.A1(n6438), 
	.A0(\ram[180][15] ));
   AOI22X1 U10550 (.Y(n12644), 
	.B1(n6457), 
	.B0(\ram[179][15] ), 
	.A1(n6476), 
	.A0(\ram[178][15] ));
   NAND4X1 U10551 (.Y(n12642), 
	.D(n12651), 
	.C(n12650), 
	.B(n12649), 
	.A(n12648));
   AOI22X1 U10552 (.Y(n12651), 
	.B1(n6495), 
	.B0(\ram[177][15] ), 
	.A1(n6514), 
	.A0(\ram[176][15] ));
   AOI22X1 U10553 (.Y(n12650), 
	.B1(n6533), 
	.B0(\ram[191][15] ), 
	.A1(n6553), 
	.A0(\ram[190][15] ));
   AOI22X1 U10554 (.Y(n12649), 
	.B1(n6572), 
	.B0(\ram[189][15] ), 
	.A1(n6591), 
	.A0(\ram[188][15] ));
   AOI22X1 U10555 (.Y(n12648), 
	.B1(n6610), 
	.B0(\ram[187][15] ), 
	.A1(n6629), 
	.A0(\ram[186][15] ));
   OAI21XL U10556 (.Y(n12629), 
	.B0(n8273), 
	.A1(n12653), 
	.A0(n12652));
   NAND4X1 U10557 (.Y(n12653), 
	.D(n12657), 
	.C(n12656), 
	.B(n12655), 
	.A(n12654));
   AOI22X1 U10558 (.Y(n12657), 
	.B1(n6342), 
	.B0(\ram[169][15] ), 
	.A1(n6362), 
	.A0(\ram[168][15] ));
   AOI22X1 U10559 (.Y(n12656), 
	.B1(n6381), 
	.B0(\ram[167][15] ), 
	.A1(n6400), 
	.A0(\ram[166][15] ));
   AOI22X1 U10560 (.Y(n12655), 
	.B1(n6419), 
	.B0(\ram[165][15] ), 
	.A1(n6438), 
	.A0(\ram[164][15] ));
   AOI22X1 U10561 (.Y(n12654), 
	.B1(n6457), 
	.B0(\ram[163][15] ), 
	.A1(n6476), 
	.A0(\ram[162][15] ));
   NAND4X1 U10562 (.Y(n12652), 
	.D(n12661), 
	.C(n12660), 
	.B(n12659), 
	.A(n12658));
   AOI22X1 U10563 (.Y(n12661), 
	.B1(n6495), 
	.B0(\ram[161][15] ), 
	.A1(n6514), 
	.A0(\ram[160][15] ));
   AOI22X1 U10564 (.Y(n12660), 
	.B1(n6533), 
	.B0(\ram[175][15] ), 
	.A1(n6553), 
	.A0(\ram[174][15] ));
   AOI22X1 U10565 (.Y(n12659), 
	.B1(n6572), 
	.B0(\ram[173][15] ), 
	.A1(n6591), 
	.A0(\ram[172][15] ));
   AOI22X1 U10566 (.Y(n12658), 
	.B1(n6610), 
	.B0(\ram[171][15] ), 
	.A1(n6629), 
	.A0(\ram[170][15] ));
   OAI21XL U10567 (.Y(n12628), 
	.B0(n8562), 
	.A1(n12663), 
	.A0(n12662));
   NAND4X1 U10568 (.Y(n12663), 
	.D(n12667), 
	.C(n12666), 
	.B(n12665), 
	.A(n12664));
   AOI22X1 U10569 (.Y(n12667), 
	.B1(n6342), 
	.B0(\ram[153][15] ), 
	.A1(n6362), 
	.A0(\ram[152][15] ));
   AOI22X1 U10570 (.Y(n12666), 
	.B1(n6381), 
	.B0(\ram[151][15] ), 
	.A1(n6400), 
	.A0(\ram[150][15] ));
   AOI22X1 U10571 (.Y(n12665), 
	.B1(n6419), 
	.B0(\ram[149][15] ), 
	.A1(n6438), 
	.A0(\ram[148][15] ));
   AOI22X1 U10572 (.Y(n12664), 
	.B1(n6457), 
	.B0(\ram[147][15] ), 
	.A1(n6476), 
	.A0(\ram[146][15] ));
   NAND4X1 U10573 (.Y(n12662), 
	.D(n12671), 
	.C(n12670), 
	.B(n12669), 
	.A(n12668));
   AOI22X1 U10574 (.Y(n12671), 
	.B1(n6495), 
	.B0(\ram[145][15] ), 
	.A1(n6514), 
	.A0(\ram[144][15] ));
   AOI22X1 U10575 (.Y(n12670), 
	.B1(n6533), 
	.B0(\ram[159][15] ), 
	.A1(n6553), 
	.A0(\ram[158][15] ));
   AOI22X1 U10576 (.Y(n12669), 
	.B1(n6572), 
	.B0(\ram[157][15] ), 
	.A1(n6591), 
	.A0(\ram[156][15] ));
   AOI22X1 U10577 (.Y(n12668), 
	.B1(n6610), 
	.B0(\ram[155][15] ), 
	.A1(n6629), 
	.A0(\ram[154][15] ));
   NAND4X1 U10578 (.Y(n12581), 
	.D(n12675), 
	.C(n12674), 
	.B(n12673), 
	.A(n12672));
   OAI21XL U10579 (.Y(n12675), 
	.B0(n8851), 
	.A1(n12677), 
	.A0(n12676));
   NAND4X1 U10580 (.Y(n12677), 
	.D(n12681), 
	.C(n12680), 
	.B(n12679), 
	.A(n12678));
   AOI22X1 U10581 (.Y(n12681), 
	.B1(n6342), 
	.B0(\ram[137][15] ), 
	.A1(n6362), 
	.A0(\ram[136][15] ));
   AOI22X1 U10582 (.Y(n12680), 
	.B1(n6381), 
	.B0(\ram[135][15] ), 
	.A1(n6400), 
	.A0(\ram[134][15] ));
   AOI22X1 U10583 (.Y(n12679), 
	.B1(n6419), 
	.B0(\ram[133][15] ), 
	.A1(n6438), 
	.A0(\ram[132][15] ));
   AOI22X1 U10584 (.Y(n12678), 
	.B1(n6457), 
	.B0(\ram[131][15] ), 
	.A1(n6476), 
	.A0(\ram[130][15] ));
   NAND4X1 U10585 (.Y(n12676), 
	.D(n12685), 
	.C(n12684), 
	.B(n12683), 
	.A(n12682));
   AOI22X1 U10586 (.Y(n12685), 
	.B1(n6495), 
	.B0(\ram[129][15] ), 
	.A1(n6514), 
	.A0(\ram[128][15] ));
   AOI22X1 U10587 (.Y(n12684), 
	.B1(n6533), 
	.B0(\ram[143][15] ), 
	.A1(n6553), 
	.A0(\ram[142][15] ));
   AOI22X1 U10588 (.Y(n12683), 
	.B1(n6572), 
	.B0(\ram[141][15] ), 
	.A1(n6591), 
	.A0(\ram[140][15] ));
   AOI22X1 U10589 (.Y(n12682), 
	.B1(n6610), 
	.B0(\ram[139][15] ), 
	.A1(n6629), 
	.A0(\ram[138][15] ));
   OAI21XL U10590 (.Y(n12674), 
	.B0(n9140), 
	.A1(n12687), 
	.A0(n12686));
   NAND4X1 U10591 (.Y(n12687), 
	.D(n12691), 
	.C(n12690), 
	.B(n12689), 
	.A(n12688));
   AOI22X1 U10592 (.Y(n12691), 
	.B1(n6342), 
	.B0(\ram[121][15] ), 
	.A1(n6362), 
	.A0(\ram[120][15] ));
   AOI22X1 U10593 (.Y(n12690), 
	.B1(n6381), 
	.B0(\ram[119][15] ), 
	.A1(n6400), 
	.A0(\ram[118][15] ));
   AOI22X1 U10594 (.Y(n12689), 
	.B1(n6419), 
	.B0(\ram[117][15] ), 
	.A1(n6438), 
	.A0(\ram[116][15] ));
   AOI22X1 U10595 (.Y(n12688), 
	.B1(n6457), 
	.B0(\ram[115][15] ), 
	.A1(n6476), 
	.A0(\ram[114][15] ));
   NAND4X1 U10596 (.Y(n12686), 
	.D(n12695), 
	.C(n12694), 
	.B(n12693), 
	.A(n12692));
   AOI22X1 U10597 (.Y(n12695), 
	.B1(n6495), 
	.B0(\ram[113][15] ), 
	.A1(n6514), 
	.A0(\ram[112][15] ));
   AOI22X1 U10598 (.Y(n12694), 
	.B1(n6533), 
	.B0(\ram[127][15] ), 
	.A1(n6553), 
	.A0(\ram[126][15] ));
   AOI22X1 U10599 (.Y(n12693), 
	.B1(n6572), 
	.B0(\ram[125][15] ), 
	.A1(n6591), 
	.A0(\ram[124][15] ));
   AOI22X1 U10600 (.Y(n12692), 
	.B1(n6610), 
	.B0(\ram[123][15] ), 
	.A1(n6629), 
	.A0(\ram[122][15] ));
   OAI21XL U10601 (.Y(n12673), 
	.B0(n9429), 
	.A1(n12697), 
	.A0(n12696));
   NAND4X1 U10602 (.Y(n12697), 
	.D(n12701), 
	.C(n12700), 
	.B(n12699), 
	.A(n12698));
   AOI22X1 U10603 (.Y(n12701), 
	.B1(n6342), 
	.B0(\ram[105][15] ), 
	.A1(n6362), 
	.A0(\ram[104][15] ));
   AOI22X1 U10604 (.Y(n12700), 
	.B1(n6381), 
	.B0(\ram[103][15] ), 
	.A1(n6400), 
	.A0(\ram[102][15] ));
   AOI22X1 U10605 (.Y(n12699), 
	.B1(n6419), 
	.B0(\ram[101][15] ), 
	.A1(n6438), 
	.A0(\ram[100][15] ));
   AOI22X1 U10606 (.Y(n12698), 
	.B1(n6457), 
	.B0(\ram[99][15] ), 
	.A1(n6476), 
	.A0(\ram[98][15] ));
   NAND4X1 U10607 (.Y(n12696), 
	.D(n12705), 
	.C(n12704), 
	.B(n12703), 
	.A(n12702));
   AOI22X1 U10608 (.Y(n12705), 
	.B1(n6495), 
	.B0(\ram[97][15] ), 
	.A1(n6514), 
	.A0(\ram[96][15] ));
   AOI22X1 U10609 (.Y(n12704), 
	.B1(n6533), 
	.B0(\ram[111][15] ), 
	.A1(n6553), 
	.A0(\ram[110][15] ));
   AOI22X1 U10610 (.Y(n12703), 
	.B1(n6572), 
	.B0(\ram[109][15] ), 
	.A1(n6591), 
	.A0(\ram[108][15] ));
   AOI22X1 U10611 (.Y(n12702), 
	.B1(n6610), 
	.B0(\ram[107][15] ), 
	.A1(n6629), 
	.A0(\ram[106][15] ));
   OAI21XL U10612 (.Y(n12672), 
	.B0(n9718), 
	.A1(n12707), 
	.A0(n12706));
   NAND4X1 U10613 (.Y(n12707), 
	.D(n12711), 
	.C(n12710), 
	.B(n12709), 
	.A(n12708));
   AOI22X1 U10614 (.Y(n12711), 
	.B1(n6342), 
	.B0(\ram[89][15] ), 
	.A1(n6362), 
	.A0(\ram[88][15] ));
   AOI22X1 U10615 (.Y(n12710), 
	.B1(n6381), 
	.B0(\ram[87][15] ), 
	.A1(n6400), 
	.A0(\ram[86][15] ));
   AOI22X1 U10616 (.Y(n12709), 
	.B1(n6419), 
	.B0(\ram[85][15] ), 
	.A1(n6438), 
	.A0(\ram[84][15] ));
   AOI22X1 U10617 (.Y(n12708), 
	.B1(n6457), 
	.B0(\ram[83][15] ), 
	.A1(n6476), 
	.A0(\ram[82][15] ));
   NAND4X1 U10618 (.Y(n12706), 
	.D(n12715), 
	.C(n12714), 
	.B(n12713), 
	.A(n12712));
   AOI22X1 U10619 (.Y(n12715), 
	.B1(n6495), 
	.B0(\ram[81][15] ), 
	.A1(n6514), 
	.A0(\ram[80][15] ));
   AOI22X1 U10620 (.Y(n12714), 
	.B1(n6533), 
	.B0(\ram[95][15] ), 
	.A1(n6553), 
	.A0(\ram[94][15] ));
   AOI22X1 U10621 (.Y(n12713), 
	.B1(n6572), 
	.B0(\ram[93][15] ), 
	.A1(n6591), 
	.A0(\ram[92][15] ));
   AOI22X1 U10622 (.Y(n12712), 
	.B1(n6610), 
	.B0(\ram[91][15] ), 
	.A1(n6629), 
	.A0(\ram[90][15] ));
   NAND4X1 U10623 (.Y(n12580), 
	.D(n12719), 
	.C(n12718), 
	.B(n12717), 
	.A(n12716));
   OAI21XL U10624 (.Y(n12719), 
	.B0(n10007), 
	.A1(n12721), 
	.A0(n12720));
   NAND4X1 U10625 (.Y(n12721), 
	.D(n12725), 
	.C(n12724), 
	.B(n12723), 
	.A(n12722));
   AOI22X1 U10626 (.Y(n12725), 
	.B1(n6342), 
	.B0(\ram[73][15] ), 
	.A1(n6362), 
	.A0(\ram[72][15] ));
   AOI22X1 U10627 (.Y(n12724), 
	.B1(n6381), 
	.B0(\ram[71][15] ), 
	.A1(n6400), 
	.A0(\ram[70][15] ));
   AOI22X1 U10628 (.Y(n12723), 
	.B1(n6419), 
	.B0(\ram[69][15] ), 
	.A1(n6438), 
	.A0(\ram[68][15] ));
   AOI22X1 U10629 (.Y(n12722), 
	.B1(n6457), 
	.B0(\ram[67][15] ), 
	.A1(n6476), 
	.A0(\ram[66][15] ));
   NAND4X1 U10630 (.Y(n12720), 
	.D(n12729), 
	.C(n12728), 
	.B(n12727), 
	.A(n12726));
   AOI22X1 U10631 (.Y(n12729), 
	.B1(n6495), 
	.B0(\ram[65][15] ), 
	.A1(n6514), 
	.A0(\ram[64][15] ));
   AOI22X1 U10632 (.Y(n12728), 
	.B1(n6533), 
	.B0(\ram[79][15] ), 
	.A1(n6553), 
	.A0(\ram[78][15] ));
   AOI22X1 U10633 (.Y(n12727), 
	.B1(n6572), 
	.B0(\ram[77][15] ), 
	.A1(n6591), 
	.A0(\ram[76][15] ));
   AOI22X1 U10634 (.Y(n12726), 
	.B1(n6610), 
	.B0(\ram[75][15] ), 
	.A1(n6629), 
	.A0(\ram[74][15] ));
   OAI21XL U10635 (.Y(n12718), 
	.B0(n10296), 
	.A1(n12731), 
	.A0(n12730));
   NAND4X1 U10636 (.Y(n12731), 
	.D(n12735), 
	.C(n12734), 
	.B(n12733), 
	.A(n12732));
   AOI22X1 U10637 (.Y(n12735), 
	.B1(n6342), 
	.B0(\ram[57][15] ), 
	.A1(n6362), 
	.A0(\ram[56][15] ));
   AOI22X1 U10638 (.Y(n12734), 
	.B1(n6381), 
	.B0(\ram[55][15] ), 
	.A1(n6400), 
	.A0(\ram[54][15] ));
   AOI22X1 U10639 (.Y(n12733), 
	.B1(n6419), 
	.B0(\ram[53][15] ), 
	.A1(n6438), 
	.A0(\ram[52][15] ));
   AOI22X1 U10640 (.Y(n12732), 
	.B1(n6457), 
	.B0(\ram[51][15] ), 
	.A1(n6476), 
	.A0(\ram[50][15] ));
   NAND4X1 U10641 (.Y(n12730), 
	.D(n12739), 
	.C(n12738), 
	.B(n12737), 
	.A(n12736));
   AOI22X1 U10642 (.Y(n12739), 
	.B1(n6495), 
	.B0(\ram[49][15] ), 
	.A1(n6514), 
	.A0(\ram[48][15] ));
   AOI22X1 U10643 (.Y(n12738), 
	.B1(n6533), 
	.B0(\ram[63][15] ), 
	.A1(n6553), 
	.A0(\ram[62][15] ));
   AOI22X1 U10644 (.Y(n12737), 
	.B1(n6572), 
	.B0(\ram[61][15] ), 
	.A1(n6591), 
	.A0(\ram[60][15] ));
   AOI22X1 U10645 (.Y(n12736), 
	.B1(n6610), 
	.B0(\ram[59][15] ), 
	.A1(n6629), 
	.A0(\ram[58][15] ));
   OAI21XL U10646 (.Y(n12717), 
	.B0(n10585), 
	.A1(n12741), 
	.A0(n12740));
   NAND4X1 U10647 (.Y(n12741), 
	.D(n12745), 
	.C(n12744), 
	.B(n12743), 
	.A(n12742));
   AOI22X1 U10648 (.Y(n12745), 
	.B1(n6342), 
	.B0(\ram[41][15] ), 
	.A1(n6362), 
	.A0(\ram[40][15] ));
   AOI22X1 U10649 (.Y(n12744), 
	.B1(n6381), 
	.B0(\ram[39][15] ), 
	.A1(n6400), 
	.A0(\ram[38][15] ));
   AOI22X1 U10650 (.Y(n12743), 
	.B1(n6419), 
	.B0(\ram[37][15] ), 
	.A1(n6438), 
	.A0(\ram[36][15] ));
   AOI22X1 U10651 (.Y(n12742), 
	.B1(n6457), 
	.B0(\ram[35][15] ), 
	.A1(n6476), 
	.A0(\ram[34][15] ));
   NAND4X1 U10652 (.Y(n12740), 
	.D(n12749), 
	.C(n12748), 
	.B(n12747), 
	.A(n12746));
   AOI22X1 U10653 (.Y(n12749), 
	.B1(n6495), 
	.B0(\ram[33][15] ), 
	.A1(n6514), 
	.A0(\ram[32][15] ));
   AOI22X1 U10654 (.Y(n12748), 
	.B1(n6533), 
	.B0(\ram[47][15] ), 
	.A1(n6553), 
	.A0(\ram[46][15] ));
   AOI22X1 U10655 (.Y(n12747), 
	.B1(n6572), 
	.B0(\ram[45][15] ), 
	.A1(n6591), 
	.A0(\ram[44][15] ));
   AOI22X1 U10656 (.Y(n12746), 
	.B1(n6610), 
	.B0(\ram[43][15] ), 
	.A1(n6629), 
	.A0(\ram[42][15] ));
   OAI21XL U10657 (.Y(n12716), 
	.B0(n6343), 
	.A1(n12751), 
	.A0(n12750));
   NAND4X1 U10658 (.Y(n12751), 
	.D(n12755), 
	.C(n12754), 
	.B(n12753), 
	.A(n12752));
   AOI22X1 U10659 (.Y(n12755), 
	.B1(n6342), 
	.B0(\ram[25][15] ), 
	.A1(n6362), 
	.A0(\ram[24][15] ));
   AOI22X1 U10660 (.Y(n12754), 
	.B1(n6381), 
	.B0(\ram[23][15] ), 
	.A1(n6400), 
	.A0(\ram[22][15] ));
   AOI22X1 U10661 (.Y(n12753), 
	.B1(n6419), 
	.B0(\ram[21][15] ), 
	.A1(n6438), 
	.A0(\ram[20][15] ));
   AOI22X1 U10662 (.Y(n12752), 
	.B1(n6457), 
	.B0(\ram[19][15] ), 
	.A1(n6476), 
	.A0(\ram[18][15] ));
   NAND4X1 U10663 (.Y(n12750), 
	.D(n12759), 
	.C(n12758), 
	.B(n12757), 
	.A(n12756));
   AOI22X1 U10664 (.Y(n12759), 
	.B1(n6495), 
	.B0(\ram[17][15] ), 
	.A1(n6514), 
	.A0(\ram[16][15] ));
   AOI22X1 U10665 (.Y(n12758), 
	.B1(n6533), 
	.B0(\ram[31][15] ), 
	.A1(n6553), 
	.A0(\ram[30][15] ));
   AOI22X1 U10666 (.Y(n12757), 
	.B1(n6572), 
	.B0(\ram[29][15] ), 
	.A1(n6591), 
	.A0(\ram[28][15] ));
   AOI22X1 U10667 (.Y(n12756), 
	.B1(n6610), 
	.B0(\ram[27][15] ), 
	.A1(n6629), 
	.A0(\ram[26][15] ));
   OR4X1 U10668 (.Y(mem_read_data[14]), 
	.D(n12763), 
	.C(n12762), 
	.B(n12761), 
	.A(n12760));
   NAND4X1 U10669 (.Y(n12763), 
	.D(n12767), 
	.C(n12766), 
	.B(n12765), 
	.A(n12764));
   OAI21XL U10670 (.Y(n12767), 
	.B0(n6534), 
	.A1(n12769), 
	.A0(n12768));
   NAND4X1 U10671 (.Y(n12769), 
	.D(n12773), 
	.C(n12772), 
	.B(n12771), 
	.A(n12770));
   AOI22X1 U10672 (.Y(n12773), 
	.B1(n6342), 
	.B0(\ram[9][14] ), 
	.A1(n6362), 
	.A0(\ram[8][14] ));
   AOI22X1 U10673 (.Y(n12772), 
	.B1(n6381), 
	.B0(\ram[7][14] ), 
	.A1(n6400), 
	.A0(\ram[6][14] ));
   AOI22X1 U10674 (.Y(n12771), 
	.B1(n6419), 
	.B0(\ram[5][14] ), 
	.A1(n6438), 
	.A0(\ram[4][14] ));
   AOI22X1 U10675 (.Y(n12770), 
	.B1(n6457), 
	.B0(\ram[3][14] ), 
	.A1(n6476), 
	.A0(\ram[2][14] ));
   NAND4X1 U10676 (.Y(n12768), 
	.D(n12777), 
	.C(n12776), 
	.B(n12775), 
	.A(n12774));
   AOI22X1 U10677 (.Y(n12777), 
	.B1(n6495), 
	.B0(\ram[1][14] ), 
	.A1(n6514), 
	.A0(\ram[0][14] ));
   AOI22X1 U10678 (.Y(n12776), 
	.B1(n6533), 
	.B0(\ram[15][14] ), 
	.A1(n6553), 
	.A0(\ram[14][14] ));
   AOI22X1 U10679 (.Y(n12775), 
	.B1(n6572), 
	.B0(\ram[13][14] ), 
	.A1(n6591), 
	.A0(\ram[12][14] ));
   AOI22X1 U10680 (.Y(n12774), 
	.B1(n6610), 
	.B0(\ram[11][14] ), 
	.A1(n6629), 
	.A0(\ram[10][14] ));
   OAI21XL U10681 (.Y(n12766), 
	.B0(n6828), 
	.A1(n12779), 
	.A0(n12778));
   NAND4X1 U10682 (.Y(n12779), 
	.D(n12783), 
	.C(n12782), 
	.B(n12781), 
	.A(n12780));
   AOI22X1 U10683 (.Y(n12783), 
	.B1(n6342), 
	.B0(\ram[249][14] ), 
	.A1(n6362), 
	.A0(\ram[248][14] ));
   AOI22X1 U10684 (.Y(n12782), 
	.B1(n6381), 
	.B0(\ram[247][14] ), 
	.A1(n6400), 
	.A0(\ram[246][14] ));
   AOI22X1 U10685 (.Y(n12781), 
	.B1(n6419), 
	.B0(\ram[245][14] ), 
	.A1(n6438), 
	.A0(\ram[244][14] ));
   AOI22X1 U10686 (.Y(n12780), 
	.B1(n6457), 
	.B0(\ram[243][14] ), 
	.A1(n6476), 
	.A0(\ram[242][14] ));
   NAND4X1 U10687 (.Y(n12778), 
	.D(n12787), 
	.C(n12786), 
	.B(n12785), 
	.A(n12784));
   AOI22X1 U10688 (.Y(n12787), 
	.B1(n6495), 
	.B0(\ram[241][14] ), 
	.A1(n6514), 
	.A0(\ram[240][14] ));
   AOI22X1 U10689 (.Y(n12786), 
	.B1(n6533), 
	.B0(\ram[255][14] ), 
	.A1(n6553), 
	.A0(\ram[254][14] ));
   AOI22X1 U10690 (.Y(n12785), 
	.B1(n6572), 
	.B0(\ram[253][14] ), 
	.A1(n6591), 
	.A0(\ram[252][14] ));
   AOI22X1 U10691 (.Y(n12784), 
	.B1(n6610), 
	.B0(\ram[251][14] ), 
	.A1(n6629), 
	.A0(\ram[250][14] ));
   OAI21XL U10692 (.Y(n12765), 
	.B0(n7117), 
	.A1(n12789), 
	.A0(n12788));
   NAND4X1 U10693 (.Y(n12789), 
	.D(n12793), 
	.C(n12792), 
	.B(n12791), 
	.A(n12790));
   AOI22X1 U10694 (.Y(n12793), 
	.B1(n6342), 
	.B0(\ram[233][14] ), 
	.A1(n6362), 
	.A0(\ram[232][14] ));
   AOI22X1 U10695 (.Y(n12792), 
	.B1(n6381), 
	.B0(\ram[231][14] ), 
	.A1(n6400), 
	.A0(\ram[230][14] ));
   AOI22X1 U10696 (.Y(n12791), 
	.B1(n6419), 
	.B0(\ram[229][14] ), 
	.A1(n6438), 
	.A0(\ram[228][14] ));
   AOI22X1 U10697 (.Y(n12790), 
	.B1(n6457), 
	.B0(\ram[227][14] ), 
	.A1(n6476), 
	.A0(\ram[226][14] ));
   NAND4X1 U10698 (.Y(n12788), 
	.D(n12797), 
	.C(n12796), 
	.B(n12795), 
	.A(n12794));
   AOI22X1 U10699 (.Y(n12797), 
	.B1(n6495), 
	.B0(\ram[225][14] ), 
	.A1(n6514), 
	.A0(\ram[224][14] ));
   AOI22X1 U10700 (.Y(n12796), 
	.B1(n6533), 
	.B0(\ram[239][14] ), 
	.A1(n6553), 
	.A0(\ram[238][14] ));
   AOI22X1 U10701 (.Y(n12795), 
	.B1(n6572), 
	.B0(\ram[237][14] ), 
	.A1(n6591), 
	.A0(\ram[236][14] ));
   AOI22X1 U10702 (.Y(n12794), 
	.B1(n6610), 
	.B0(\ram[235][14] ), 
	.A1(n6629), 
	.A0(\ram[234][14] ));
   OAI21XL U10703 (.Y(n12764), 
	.B0(n7406), 
	.A1(n12799), 
	.A0(n12798));
   NAND4X1 U10704 (.Y(n12799), 
	.D(n12803), 
	.C(n12802), 
	.B(n12801), 
	.A(n12800));
   AOI22X1 U10705 (.Y(n12803), 
	.B1(n6342), 
	.B0(\ram[217][14] ), 
	.A1(n6362), 
	.A0(\ram[216][14] ));
   AOI22X1 U10706 (.Y(n12802), 
	.B1(n6381), 
	.B0(\ram[215][14] ), 
	.A1(n6400), 
	.A0(\ram[214][14] ));
   AOI22X1 U10707 (.Y(n12801), 
	.B1(n6419), 
	.B0(\ram[213][14] ), 
	.A1(n6438), 
	.A0(\ram[212][14] ));
   AOI22X1 U10708 (.Y(n12800), 
	.B1(n6457), 
	.B0(\ram[211][14] ), 
	.A1(n6476), 
	.A0(\ram[210][14] ));
   NAND4X1 U10709 (.Y(n12798), 
	.D(n12807), 
	.C(n12806), 
	.B(n12805), 
	.A(n12804));
   AOI22X1 U10710 (.Y(n12807), 
	.B1(n6495), 
	.B0(\ram[209][14] ), 
	.A1(n6514), 
	.A0(\ram[208][14] ));
   AOI22X1 U10711 (.Y(n12806), 
	.B1(n6533), 
	.B0(\ram[223][14] ), 
	.A1(n6553), 
	.A0(\ram[222][14] ));
   AOI22X1 U10712 (.Y(n12805), 
	.B1(n6572), 
	.B0(\ram[221][14] ), 
	.A1(n6591), 
	.A0(\ram[220][14] ));
   AOI22X1 U10713 (.Y(n12804), 
	.B1(n6610), 
	.B0(\ram[219][14] ), 
	.A1(n6629), 
	.A0(\ram[218][14] ));
   NAND4X1 U10714 (.Y(n12762), 
	.D(n12811), 
	.C(n12810), 
	.B(n12809), 
	.A(n12808));
   OAI21XL U10715 (.Y(n12811), 
	.B0(n7695), 
	.A1(n12813), 
	.A0(n12812));
   NAND4X1 U10716 (.Y(n12813), 
	.D(n12817), 
	.C(n12816), 
	.B(n12815), 
	.A(n12814));
   AOI22X1 U10717 (.Y(n12817), 
	.B1(n6342), 
	.B0(\ram[201][14] ), 
	.A1(n6362), 
	.A0(\ram[200][14] ));
   AOI22X1 U10718 (.Y(n12816), 
	.B1(n6381), 
	.B0(\ram[199][14] ), 
	.A1(n6400), 
	.A0(\ram[198][14] ));
   AOI22X1 U10719 (.Y(n12815), 
	.B1(n6419), 
	.B0(\ram[197][14] ), 
	.A1(n6438), 
	.A0(\ram[196][14] ));
   AOI22X1 U10720 (.Y(n12814), 
	.B1(n6457), 
	.B0(\ram[195][14] ), 
	.A1(n6476), 
	.A0(\ram[194][14] ));
   NAND4X1 U10721 (.Y(n12812), 
	.D(n12821), 
	.C(n12820), 
	.B(n12819), 
	.A(n12818));
   AOI22X1 U10722 (.Y(n12821), 
	.B1(n6495), 
	.B0(\ram[193][14] ), 
	.A1(n6514), 
	.A0(\ram[192][14] ));
   AOI22X1 U10723 (.Y(n12820), 
	.B1(n6533), 
	.B0(\ram[207][14] ), 
	.A1(n6553), 
	.A0(\ram[206][14] ));
   AOI22X1 U10724 (.Y(n12819), 
	.B1(n6572), 
	.B0(\ram[205][14] ), 
	.A1(n6591), 
	.A0(\ram[204][14] ));
   AOI22X1 U10725 (.Y(n12818), 
	.B1(n6610), 
	.B0(\ram[203][14] ), 
	.A1(n6629), 
	.A0(\ram[202][14] ));
   OAI21XL U10726 (.Y(n12810), 
	.B0(n7984), 
	.A1(n12823), 
	.A0(n12822));
   NAND4X1 U10727 (.Y(n12823), 
	.D(n12827), 
	.C(n12826), 
	.B(n12825), 
	.A(n12824));
   AOI22X1 U10728 (.Y(n12827), 
	.B1(n6342), 
	.B0(\ram[185][14] ), 
	.A1(n6362), 
	.A0(\ram[184][14] ));
   AOI22X1 U10729 (.Y(n12826), 
	.B1(n6381), 
	.B0(\ram[183][14] ), 
	.A1(n6400), 
	.A0(\ram[182][14] ));
   AOI22X1 U10730 (.Y(n12825), 
	.B1(n6419), 
	.B0(\ram[181][14] ), 
	.A1(n6438), 
	.A0(\ram[180][14] ));
   AOI22X1 U10731 (.Y(n12824), 
	.B1(n6457), 
	.B0(\ram[179][14] ), 
	.A1(n6476), 
	.A0(\ram[178][14] ));
   NAND4X1 U10732 (.Y(n12822), 
	.D(n12831), 
	.C(n12830), 
	.B(n12829), 
	.A(n12828));
   AOI22X1 U10733 (.Y(n12831), 
	.B1(n6495), 
	.B0(\ram[177][14] ), 
	.A1(n6514), 
	.A0(\ram[176][14] ));
   AOI22X1 U10734 (.Y(n12830), 
	.B1(n6533), 
	.B0(\ram[191][14] ), 
	.A1(n6553), 
	.A0(\ram[190][14] ));
   AOI22X1 U10735 (.Y(n12829), 
	.B1(n6572), 
	.B0(\ram[189][14] ), 
	.A1(n6591), 
	.A0(\ram[188][14] ));
   AOI22X1 U10736 (.Y(n12828), 
	.B1(n6610), 
	.B0(\ram[187][14] ), 
	.A1(n6629), 
	.A0(\ram[186][14] ));
   OAI21XL U10737 (.Y(n12809), 
	.B0(n8273), 
	.A1(n12833), 
	.A0(n12832));
   NAND4X1 U10738 (.Y(n12833), 
	.D(n12837), 
	.C(n12836), 
	.B(n12835), 
	.A(n12834));
   AOI22X1 U10739 (.Y(n12837), 
	.B1(n6342), 
	.B0(\ram[169][14] ), 
	.A1(n6362), 
	.A0(\ram[168][14] ));
   AOI22X1 U10740 (.Y(n12836), 
	.B1(n6381), 
	.B0(\ram[167][14] ), 
	.A1(n6400), 
	.A0(\ram[166][14] ));
   AOI22X1 U10741 (.Y(n12835), 
	.B1(n6419), 
	.B0(\ram[165][14] ), 
	.A1(n6438), 
	.A0(\ram[164][14] ));
   AOI22X1 U10742 (.Y(n12834), 
	.B1(n6457), 
	.B0(\ram[163][14] ), 
	.A1(n6476), 
	.A0(\ram[162][14] ));
   NAND4X1 U10743 (.Y(n12832), 
	.D(n12841), 
	.C(n12840), 
	.B(n12839), 
	.A(n12838));
   AOI22X1 U10744 (.Y(n12841), 
	.B1(n6495), 
	.B0(\ram[161][14] ), 
	.A1(n6514), 
	.A0(\ram[160][14] ));
   AOI22X1 U10745 (.Y(n12840), 
	.B1(n6533), 
	.B0(\ram[175][14] ), 
	.A1(n6553), 
	.A0(\ram[174][14] ));
   AOI22X1 U10746 (.Y(n12839), 
	.B1(n6572), 
	.B0(\ram[173][14] ), 
	.A1(n6591), 
	.A0(\ram[172][14] ));
   AOI22X1 U10747 (.Y(n12838), 
	.B1(n6610), 
	.B0(\ram[171][14] ), 
	.A1(n6629), 
	.A0(\ram[170][14] ));
   OAI21XL U10748 (.Y(n12808), 
	.B0(n8562), 
	.A1(n12843), 
	.A0(n12842));
   NAND4X1 U10749 (.Y(n12843), 
	.D(n12847), 
	.C(n12846), 
	.B(n12845), 
	.A(n12844));
   AOI22X1 U10750 (.Y(n12847), 
	.B1(n6342), 
	.B0(\ram[153][14] ), 
	.A1(n6362), 
	.A0(\ram[152][14] ));
   AOI22X1 U10751 (.Y(n12846), 
	.B1(n6381), 
	.B0(\ram[151][14] ), 
	.A1(n6400), 
	.A0(\ram[150][14] ));
   AOI22X1 U10752 (.Y(n12845), 
	.B1(n6419), 
	.B0(\ram[149][14] ), 
	.A1(n6438), 
	.A0(\ram[148][14] ));
   AOI22X1 U10753 (.Y(n12844), 
	.B1(n6457), 
	.B0(\ram[147][14] ), 
	.A1(n6476), 
	.A0(\ram[146][14] ));
   NAND4X1 U10754 (.Y(n12842), 
	.D(n12851), 
	.C(n12850), 
	.B(n12849), 
	.A(n12848));
   AOI22X1 U10755 (.Y(n12851), 
	.B1(n6495), 
	.B0(\ram[145][14] ), 
	.A1(n6514), 
	.A0(\ram[144][14] ));
   AOI22X1 U10756 (.Y(n12850), 
	.B1(n6533), 
	.B0(\ram[159][14] ), 
	.A1(n6553), 
	.A0(\ram[158][14] ));
   AOI22X1 U10757 (.Y(n12849), 
	.B1(n6572), 
	.B0(\ram[157][14] ), 
	.A1(n6591), 
	.A0(\ram[156][14] ));
   AOI22X1 U10758 (.Y(n12848), 
	.B1(n6610), 
	.B0(\ram[155][14] ), 
	.A1(n6629), 
	.A0(\ram[154][14] ));
   NAND4X1 U10759 (.Y(n12761), 
	.D(n12855), 
	.C(n12854), 
	.B(n12853), 
	.A(n12852));
   OAI21XL U10760 (.Y(n12855), 
	.B0(n8851), 
	.A1(n12857), 
	.A0(n12856));
   NAND4X1 U10761 (.Y(n12857), 
	.D(n12861), 
	.C(n12860), 
	.B(n12859), 
	.A(n12858));
   AOI22X1 U10762 (.Y(n12861), 
	.B1(n6342), 
	.B0(\ram[137][14] ), 
	.A1(n6362), 
	.A0(\ram[136][14] ));
   AOI22X1 U10763 (.Y(n12860), 
	.B1(n6381), 
	.B0(\ram[135][14] ), 
	.A1(n6400), 
	.A0(\ram[134][14] ));
   AOI22X1 U10764 (.Y(n12859), 
	.B1(n6419), 
	.B0(\ram[133][14] ), 
	.A1(n6438), 
	.A0(\ram[132][14] ));
   AOI22X1 U10765 (.Y(n12858), 
	.B1(n6457), 
	.B0(\ram[131][14] ), 
	.A1(n6476), 
	.A0(\ram[130][14] ));
   NAND4X1 U10766 (.Y(n12856), 
	.D(n12865), 
	.C(n12864), 
	.B(n12863), 
	.A(n12862));
   AOI22X1 U10767 (.Y(n12865), 
	.B1(n6495), 
	.B0(\ram[129][14] ), 
	.A1(n6514), 
	.A0(\ram[128][14] ));
   AOI22X1 U10768 (.Y(n12864), 
	.B1(n6533), 
	.B0(\ram[143][14] ), 
	.A1(n6553), 
	.A0(\ram[142][14] ));
   AOI22X1 U10769 (.Y(n12863), 
	.B1(n6572), 
	.B0(\ram[141][14] ), 
	.A1(n6591), 
	.A0(\ram[140][14] ));
   AOI22X1 U10770 (.Y(n12862), 
	.B1(n6610), 
	.B0(\ram[139][14] ), 
	.A1(n6629), 
	.A0(\ram[138][14] ));
   OAI21XL U10771 (.Y(n12854), 
	.B0(n9140), 
	.A1(n12867), 
	.A0(n12866));
   NAND4X1 U10772 (.Y(n12867), 
	.D(n12871), 
	.C(n12870), 
	.B(n12869), 
	.A(n12868));
   AOI22X1 U10773 (.Y(n12871), 
	.B1(n6342), 
	.B0(\ram[121][14] ), 
	.A1(n6362), 
	.A0(\ram[120][14] ));
   AOI22X1 U10774 (.Y(n12870), 
	.B1(n6381), 
	.B0(\ram[119][14] ), 
	.A1(n6400), 
	.A0(\ram[118][14] ));
   AOI22X1 U10775 (.Y(n12869), 
	.B1(n6419), 
	.B0(\ram[117][14] ), 
	.A1(n6438), 
	.A0(\ram[116][14] ));
   AOI22X1 U10776 (.Y(n12868), 
	.B1(n6457), 
	.B0(\ram[115][14] ), 
	.A1(n6476), 
	.A0(\ram[114][14] ));
   NAND4X1 U10777 (.Y(n12866), 
	.D(n12875), 
	.C(n12874), 
	.B(n12873), 
	.A(n12872));
   AOI22X1 U10778 (.Y(n12875), 
	.B1(n6495), 
	.B0(\ram[113][14] ), 
	.A1(n6514), 
	.A0(\ram[112][14] ));
   AOI22X1 U10779 (.Y(n12874), 
	.B1(n6533), 
	.B0(\ram[127][14] ), 
	.A1(n6553), 
	.A0(\ram[126][14] ));
   AOI22X1 U10780 (.Y(n12873), 
	.B1(n6572), 
	.B0(\ram[125][14] ), 
	.A1(n6591), 
	.A0(\ram[124][14] ));
   AOI22X1 U10781 (.Y(n12872), 
	.B1(n6610), 
	.B0(\ram[123][14] ), 
	.A1(n6629), 
	.A0(\ram[122][14] ));
   OAI21XL U10782 (.Y(n12853), 
	.B0(n9429), 
	.A1(n12877), 
	.A0(n12876));
   NAND4X1 U10783 (.Y(n12877), 
	.D(n12881), 
	.C(n12880), 
	.B(n12879), 
	.A(n12878));
   AOI22X1 U10784 (.Y(n12881), 
	.B1(n6342), 
	.B0(\ram[105][14] ), 
	.A1(n6362), 
	.A0(\ram[104][14] ));
   AOI22X1 U10785 (.Y(n12880), 
	.B1(n6381), 
	.B0(\ram[103][14] ), 
	.A1(n6400), 
	.A0(\ram[102][14] ));
   AOI22X1 U10786 (.Y(n12879), 
	.B1(n6419), 
	.B0(\ram[101][14] ), 
	.A1(n6438), 
	.A0(\ram[100][14] ));
   AOI22X1 U10787 (.Y(n12878), 
	.B1(n6457), 
	.B0(\ram[99][14] ), 
	.A1(n6476), 
	.A0(\ram[98][14] ));
   NAND4X1 U10788 (.Y(n12876), 
	.D(n12885), 
	.C(n12884), 
	.B(n12883), 
	.A(n12882));
   AOI22X1 U10789 (.Y(n12885), 
	.B1(n6495), 
	.B0(\ram[97][14] ), 
	.A1(n6514), 
	.A0(\ram[96][14] ));
   AOI22X1 U10790 (.Y(n12884), 
	.B1(n6533), 
	.B0(\ram[111][14] ), 
	.A1(n6553), 
	.A0(\ram[110][14] ));
   AOI22X1 U10791 (.Y(n12883), 
	.B1(n6572), 
	.B0(\ram[109][14] ), 
	.A1(n6591), 
	.A0(\ram[108][14] ));
   AOI22X1 U10792 (.Y(n12882), 
	.B1(n6610), 
	.B0(\ram[107][14] ), 
	.A1(n6629), 
	.A0(\ram[106][14] ));
   OAI21XL U10793 (.Y(n12852), 
	.B0(n9718), 
	.A1(n12887), 
	.A0(n12886));
   NAND4X1 U10794 (.Y(n12887), 
	.D(n12891), 
	.C(n12890), 
	.B(n12889), 
	.A(n12888));
   AOI22X1 U10795 (.Y(n12891), 
	.B1(n6342), 
	.B0(\ram[89][14] ), 
	.A1(n6362), 
	.A0(\ram[88][14] ));
   AOI22X1 U10796 (.Y(n12890), 
	.B1(n6381), 
	.B0(\ram[87][14] ), 
	.A1(n6400), 
	.A0(\ram[86][14] ));
   AOI22X1 U10797 (.Y(n12889), 
	.B1(n6419), 
	.B0(\ram[85][14] ), 
	.A1(n6438), 
	.A0(\ram[84][14] ));
   AOI22X1 U10798 (.Y(n12888), 
	.B1(n6457), 
	.B0(\ram[83][14] ), 
	.A1(n6476), 
	.A0(\ram[82][14] ));
   NAND4X1 U10799 (.Y(n12886), 
	.D(n12895), 
	.C(n12894), 
	.B(n12893), 
	.A(n12892));
   AOI22X1 U10800 (.Y(n12895), 
	.B1(n6495), 
	.B0(\ram[81][14] ), 
	.A1(n6514), 
	.A0(\ram[80][14] ));
   AOI22X1 U10801 (.Y(n12894), 
	.B1(n6533), 
	.B0(\ram[95][14] ), 
	.A1(n6553), 
	.A0(\ram[94][14] ));
   AOI22X1 U10802 (.Y(n12893), 
	.B1(n6572), 
	.B0(\ram[93][14] ), 
	.A1(n6591), 
	.A0(\ram[92][14] ));
   AOI22X1 U10803 (.Y(n12892), 
	.B1(n6610), 
	.B0(\ram[91][14] ), 
	.A1(n6629), 
	.A0(\ram[90][14] ));
   NAND4X1 U10804 (.Y(n12760), 
	.D(n12899), 
	.C(n12898), 
	.B(n12897), 
	.A(n12896));
   OAI21XL U10805 (.Y(n12899), 
	.B0(n10007), 
	.A1(n12901), 
	.A0(n12900));
   NAND4X1 U10806 (.Y(n12901), 
	.D(n12905), 
	.C(n12904), 
	.B(n12903), 
	.A(n12902));
   AOI22X1 U10807 (.Y(n12905), 
	.B1(n6342), 
	.B0(\ram[73][14] ), 
	.A1(n6362), 
	.A0(\ram[72][14] ));
   AOI22X1 U10808 (.Y(n12904), 
	.B1(n6381), 
	.B0(\ram[71][14] ), 
	.A1(n6400), 
	.A0(\ram[70][14] ));
   AOI22X1 U10809 (.Y(n12903), 
	.B1(n6419), 
	.B0(\ram[69][14] ), 
	.A1(n6438), 
	.A0(\ram[68][14] ));
   AOI22X1 U10810 (.Y(n12902), 
	.B1(n6457), 
	.B0(\ram[67][14] ), 
	.A1(n6476), 
	.A0(\ram[66][14] ));
   NAND4X1 U10811 (.Y(n12900), 
	.D(n12909), 
	.C(n12908), 
	.B(n12907), 
	.A(n12906));
   AOI22X1 U10812 (.Y(n12909), 
	.B1(n6495), 
	.B0(\ram[65][14] ), 
	.A1(n6514), 
	.A0(\ram[64][14] ));
   AOI22X1 U10813 (.Y(n12908), 
	.B1(n6533), 
	.B0(\ram[79][14] ), 
	.A1(n6553), 
	.A0(\ram[78][14] ));
   AOI22X1 U10814 (.Y(n12907), 
	.B1(n6572), 
	.B0(\ram[77][14] ), 
	.A1(n6591), 
	.A0(\ram[76][14] ));
   AOI22X1 U10815 (.Y(n12906), 
	.B1(n6610), 
	.B0(\ram[75][14] ), 
	.A1(n6629), 
	.A0(\ram[74][14] ));
   OAI21XL U10816 (.Y(n12898), 
	.B0(n10296), 
	.A1(n12911), 
	.A0(n12910));
   NAND4X1 U10817 (.Y(n12911), 
	.D(n12915), 
	.C(n12914), 
	.B(n12913), 
	.A(n12912));
   AOI22X1 U10818 (.Y(n12915), 
	.B1(n6342), 
	.B0(\ram[57][14] ), 
	.A1(n6362), 
	.A0(\ram[56][14] ));
   AOI22X1 U10819 (.Y(n12914), 
	.B1(n6381), 
	.B0(\ram[55][14] ), 
	.A1(n6400), 
	.A0(\ram[54][14] ));
   AOI22X1 U10820 (.Y(n12913), 
	.B1(n6419), 
	.B0(\ram[53][14] ), 
	.A1(n6438), 
	.A0(\ram[52][14] ));
   AOI22X1 U10821 (.Y(n12912), 
	.B1(n6457), 
	.B0(\ram[51][14] ), 
	.A1(n6476), 
	.A0(\ram[50][14] ));
   NAND4X1 U10822 (.Y(n12910), 
	.D(n12919), 
	.C(n12918), 
	.B(n12917), 
	.A(n12916));
   AOI22X1 U10823 (.Y(n12919), 
	.B1(n6495), 
	.B0(\ram[49][14] ), 
	.A1(n6514), 
	.A0(\ram[48][14] ));
   AOI22X1 U10824 (.Y(n12918), 
	.B1(n6533), 
	.B0(\ram[63][14] ), 
	.A1(n6553), 
	.A0(\ram[62][14] ));
   AOI22X1 U10825 (.Y(n12917), 
	.B1(n6572), 
	.B0(\ram[61][14] ), 
	.A1(n6591), 
	.A0(\ram[60][14] ));
   AOI22X1 U10826 (.Y(n12916), 
	.B1(n6610), 
	.B0(\ram[59][14] ), 
	.A1(n6629), 
	.A0(\ram[58][14] ));
   OAI21XL U10827 (.Y(n12897), 
	.B0(n10585), 
	.A1(n12921), 
	.A0(n12920));
   NAND4X1 U10828 (.Y(n12921), 
	.D(n12925), 
	.C(n12924), 
	.B(n12923), 
	.A(n12922));
   AOI22X1 U10829 (.Y(n12925), 
	.B1(n6342), 
	.B0(\ram[41][14] ), 
	.A1(n6362), 
	.A0(\ram[40][14] ));
   AOI22X1 U10830 (.Y(n12924), 
	.B1(n6381), 
	.B0(\ram[39][14] ), 
	.A1(n6400), 
	.A0(\ram[38][14] ));
   AOI22X1 U10831 (.Y(n12923), 
	.B1(n6419), 
	.B0(\ram[37][14] ), 
	.A1(n6438), 
	.A0(\ram[36][14] ));
   AOI22X1 U10832 (.Y(n12922), 
	.B1(n6457), 
	.B0(\ram[35][14] ), 
	.A1(n6476), 
	.A0(\ram[34][14] ));
   NAND4X1 U10833 (.Y(n12920), 
	.D(n12929), 
	.C(n12928), 
	.B(n12927), 
	.A(n12926));
   AOI22X1 U10834 (.Y(n12929), 
	.B1(n6495), 
	.B0(\ram[33][14] ), 
	.A1(n6514), 
	.A0(\ram[32][14] ));
   AOI22X1 U10835 (.Y(n12928), 
	.B1(n6533), 
	.B0(\ram[47][14] ), 
	.A1(n6553), 
	.A0(\ram[46][14] ));
   AOI22X1 U10836 (.Y(n12927), 
	.B1(n6572), 
	.B0(\ram[45][14] ), 
	.A1(n6591), 
	.A0(\ram[44][14] ));
   AOI22X1 U10837 (.Y(n12926), 
	.B1(n6610), 
	.B0(\ram[43][14] ), 
	.A1(n6629), 
	.A0(\ram[42][14] ));
   OAI21XL U10838 (.Y(n12896), 
	.B0(n6343), 
	.A1(n12931), 
	.A0(n12930));
   NAND4X1 U10839 (.Y(n12931), 
	.D(n12935), 
	.C(n12934), 
	.B(n12933), 
	.A(n12932));
   AOI22X1 U10840 (.Y(n12935), 
	.B1(n6342), 
	.B0(\ram[25][14] ), 
	.A1(n6362), 
	.A0(\ram[24][14] ));
   AOI22X1 U10841 (.Y(n12934), 
	.B1(n6381), 
	.B0(\ram[23][14] ), 
	.A1(n6400), 
	.A0(\ram[22][14] ));
   AOI22X1 U10842 (.Y(n12933), 
	.B1(n6419), 
	.B0(\ram[21][14] ), 
	.A1(n6438), 
	.A0(\ram[20][14] ));
   AOI22X1 U10843 (.Y(n12932), 
	.B1(n6457), 
	.B0(\ram[19][14] ), 
	.A1(n6476), 
	.A0(\ram[18][14] ));
   NAND4X1 U10844 (.Y(n12930), 
	.D(n12939), 
	.C(n12938), 
	.B(n12937), 
	.A(n12936));
   AOI22X1 U10845 (.Y(n12939), 
	.B1(n6495), 
	.B0(\ram[17][14] ), 
	.A1(n6514), 
	.A0(\ram[16][14] ));
   AOI22X1 U10846 (.Y(n12938), 
	.B1(n6533), 
	.B0(\ram[31][14] ), 
	.A1(n6553), 
	.A0(\ram[30][14] ));
   AOI22X1 U10847 (.Y(n12937), 
	.B1(n6572), 
	.B0(\ram[29][14] ), 
	.A1(n6591), 
	.A0(\ram[28][14] ));
   AOI22X1 U10848 (.Y(n12936), 
	.B1(n6610), 
	.B0(\ram[27][14] ), 
	.A1(n6629), 
	.A0(\ram[26][14] ));
   OR4X1 U10849 (.Y(mem_read_data[13]), 
	.D(n12943), 
	.C(n12942), 
	.B(n12941), 
	.A(n12940));
   NAND4X1 U10850 (.Y(n12943), 
	.D(n12947), 
	.C(n12946), 
	.B(n12945), 
	.A(n12944));
   OAI21XL U10851 (.Y(n12947), 
	.B0(n6534), 
	.A1(n12949), 
	.A0(n12948));
   NAND4X1 U10852 (.Y(n12949), 
	.D(n12953), 
	.C(n12952), 
	.B(n12951), 
	.A(n12950));
   AOI22X1 U10853 (.Y(n12953), 
	.B1(n6342), 
	.B0(\ram[9][13] ), 
	.A1(n6362), 
	.A0(\ram[8][13] ));
   AOI22X1 U10854 (.Y(n12952), 
	.B1(n6381), 
	.B0(\ram[7][13] ), 
	.A1(n6400), 
	.A0(\ram[6][13] ));
   AOI22X1 U10855 (.Y(n12951), 
	.B1(n6419), 
	.B0(\ram[5][13] ), 
	.A1(n6438), 
	.A0(\ram[4][13] ));
   AOI22X1 U10856 (.Y(n12950), 
	.B1(n6457), 
	.B0(\ram[3][13] ), 
	.A1(n6476), 
	.A0(\ram[2][13] ));
   NAND4X1 U10857 (.Y(n12948), 
	.D(n12957), 
	.C(n12956), 
	.B(n12955), 
	.A(n12954));
   AOI22X1 U10858 (.Y(n12957), 
	.B1(n6495), 
	.B0(\ram[1][13] ), 
	.A1(n6514), 
	.A0(\ram[0][13] ));
   AOI22X1 U10859 (.Y(n12956), 
	.B1(n6533), 
	.B0(\ram[15][13] ), 
	.A1(n6553), 
	.A0(\ram[14][13] ));
   AOI22X1 U10860 (.Y(n12955), 
	.B1(n6572), 
	.B0(\ram[13][13] ), 
	.A1(n6591), 
	.A0(\ram[12][13] ));
   AOI22X1 U10861 (.Y(n12954), 
	.B1(n6610), 
	.B0(\ram[11][13] ), 
	.A1(n6629), 
	.A0(\ram[10][13] ));
   OAI21XL U10862 (.Y(n12946), 
	.B0(n6828), 
	.A1(n12959), 
	.A0(n12958));
   NAND4X1 U10863 (.Y(n12959), 
	.D(n12963), 
	.C(n12962), 
	.B(n12961), 
	.A(n12960));
   AOI22X1 U10864 (.Y(n12963), 
	.B1(n6342), 
	.B0(\ram[249][13] ), 
	.A1(n6362), 
	.A0(\ram[248][13] ));
   AOI22X1 U10865 (.Y(n12962), 
	.B1(n6381), 
	.B0(\ram[247][13] ), 
	.A1(n6400), 
	.A0(\ram[246][13] ));
   AOI22X1 U10866 (.Y(n12961), 
	.B1(n6419), 
	.B0(\ram[245][13] ), 
	.A1(n6438), 
	.A0(\ram[244][13] ));
   AOI22X1 U10867 (.Y(n12960), 
	.B1(n6457), 
	.B0(\ram[243][13] ), 
	.A1(n6476), 
	.A0(\ram[242][13] ));
   NAND4X1 U10868 (.Y(n12958), 
	.D(n12967), 
	.C(n12966), 
	.B(n12965), 
	.A(n12964));
   AOI22X1 U10869 (.Y(n12967), 
	.B1(n6495), 
	.B0(\ram[241][13] ), 
	.A1(n6514), 
	.A0(\ram[240][13] ));
   AOI22X1 U10870 (.Y(n12966), 
	.B1(n6533), 
	.B0(\ram[255][13] ), 
	.A1(n6553), 
	.A0(\ram[254][13] ));
   AOI22X1 U10871 (.Y(n12965), 
	.B1(n6572), 
	.B0(\ram[253][13] ), 
	.A1(n6591), 
	.A0(\ram[252][13] ));
   AOI22X1 U10872 (.Y(n12964), 
	.B1(n6610), 
	.B0(\ram[251][13] ), 
	.A1(n6629), 
	.A0(\ram[250][13] ));
   OAI21XL U10873 (.Y(n12945), 
	.B0(n7117), 
	.A1(n12969), 
	.A0(n12968));
   NAND4X1 U10874 (.Y(n12969), 
	.D(n12973), 
	.C(n12972), 
	.B(n12971), 
	.A(n12970));
   AOI22X1 U10875 (.Y(n12973), 
	.B1(n6342), 
	.B0(\ram[233][13] ), 
	.A1(n6362), 
	.A0(\ram[232][13] ));
   AOI22X1 U10876 (.Y(n12972), 
	.B1(n6381), 
	.B0(\ram[231][13] ), 
	.A1(n6400), 
	.A0(\ram[230][13] ));
   AOI22X1 U10877 (.Y(n12971), 
	.B1(n6419), 
	.B0(\ram[229][13] ), 
	.A1(n6438), 
	.A0(\ram[228][13] ));
   AOI22X1 U10878 (.Y(n12970), 
	.B1(n6457), 
	.B0(\ram[227][13] ), 
	.A1(n6476), 
	.A0(\ram[226][13] ));
   NAND4X1 U10879 (.Y(n12968), 
	.D(n12977), 
	.C(n12976), 
	.B(n12975), 
	.A(n12974));
   AOI22X1 U10880 (.Y(n12977), 
	.B1(n6495), 
	.B0(\ram[225][13] ), 
	.A1(n6514), 
	.A0(\ram[224][13] ));
   AOI22X1 U10881 (.Y(n12976), 
	.B1(n6533), 
	.B0(\ram[239][13] ), 
	.A1(n6553), 
	.A0(\ram[238][13] ));
   AOI22X1 U10882 (.Y(n12975), 
	.B1(n6572), 
	.B0(\ram[237][13] ), 
	.A1(n6591), 
	.A0(\ram[236][13] ));
   AOI22X1 U10883 (.Y(n12974), 
	.B1(n6610), 
	.B0(\ram[235][13] ), 
	.A1(n6629), 
	.A0(\ram[234][13] ));
   OAI21XL U10884 (.Y(n12944), 
	.B0(n7406), 
	.A1(n12979), 
	.A0(n12978));
   NAND4X1 U10885 (.Y(n12979), 
	.D(n12983), 
	.C(n12982), 
	.B(n12981), 
	.A(n12980));
   AOI22X1 U10886 (.Y(n12983), 
	.B1(n6342), 
	.B0(\ram[217][13] ), 
	.A1(n6362), 
	.A0(\ram[216][13] ));
   AOI22X1 U10887 (.Y(n12982), 
	.B1(n6381), 
	.B0(\ram[215][13] ), 
	.A1(n6400), 
	.A0(\ram[214][13] ));
   AOI22X1 U10888 (.Y(n12981), 
	.B1(n6419), 
	.B0(\ram[213][13] ), 
	.A1(n6438), 
	.A0(\ram[212][13] ));
   AOI22X1 U10889 (.Y(n12980), 
	.B1(n6457), 
	.B0(\ram[211][13] ), 
	.A1(n6476), 
	.A0(\ram[210][13] ));
   NAND4X1 U10890 (.Y(n12978), 
	.D(n12987), 
	.C(n12986), 
	.B(n12985), 
	.A(n12984));
   AOI22X1 U10891 (.Y(n12987), 
	.B1(n6495), 
	.B0(\ram[209][13] ), 
	.A1(n6514), 
	.A0(\ram[208][13] ));
   AOI22X1 U10892 (.Y(n12986), 
	.B1(n6533), 
	.B0(\ram[223][13] ), 
	.A1(n6553), 
	.A0(\ram[222][13] ));
   AOI22X1 U10893 (.Y(n12985), 
	.B1(n6572), 
	.B0(\ram[221][13] ), 
	.A1(n6591), 
	.A0(\ram[220][13] ));
   AOI22X1 U10894 (.Y(n12984), 
	.B1(n6610), 
	.B0(\ram[219][13] ), 
	.A1(n6629), 
	.A0(\ram[218][13] ));
   NAND4X1 U10895 (.Y(n12942), 
	.D(n12991), 
	.C(n12990), 
	.B(n12989), 
	.A(n12988));
   OAI21XL U10896 (.Y(n12991), 
	.B0(n7695), 
	.A1(n12993), 
	.A0(n12992));
   NAND4X1 U10897 (.Y(n12993), 
	.D(n12997), 
	.C(n12996), 
	.B(n12995), 
	.A(n12994));
   AOI22X1 U10898 (.Y(n12997), 
	.B1(n6342), 
	.B0(\ram[201][13] ), 
	.A1(n6362), 
	.A0(\ram[200][13] ));
   AOI22X1 U10899 (.Y(n12996), 
	.B1(n6381), 
	.B0(\ram[199][13] ), 
	.A1(n6400), 
	.A0(\ram[198][13] ));
   AOI22X1 U10900 (.Y(n12995), 
	.B1(n6419), 
	.B0(\ram[197][13] ), 
	.A1(n6438), 
	.A0(\ram[196][13] ));
   AOI22X1 U10901 (.Y(n12994), 
	.B1(n6457), 
	.B0(\ram[195][13] ), 
	.A1(n6476), 
	.A0(\ram[194][13] ));
   NAND4X1 U10902 (.Y(n12992), 
	.D(n13001), 
	.C(n13000), 
	.B(n12999), 
	.A(n12998));
   AOI22X1 U10903 (.Y(n13001), 
	.B1(n6495), 
	.B0(\ram[193][13] ), 
	.A1(n6514), 
	.A0(\ram[192][13] ));
   AOI22X1 U10904 (.Y(n13000), 
	.B1(n6533), 
	.B0(\ram[207][13] ), 
	.A1(n6553), 
	.A0(\ram[206][13] ));
   AOI22X1 U10905 (.Y(n12999), 
	.B1(n6572), 
	.B0(\ram[205][13] ), 
	.A1(n6591), 
	.A0(\ram[204][13] ));
   AOI22X1 U10906 (.Y(n12998), 
	.B1(n6610), 
	.B0(\ram[203][13] ), 
	.A1(n6629), 
	.A0(\ram[202][13] ));
   OAI21XL U10907 (.Y(n12990), 
	.B0(n7984), 
	.A1(n13003), 
	.A0(n13002));
   NAND4X1 U10908 (.Y(n13003), 
	.D(n13007), 
	.C(n13006), 
	.B(n13005), 
	.A(n13004));
   AOI22X1 U10909 (.Y(n13007), 
	.B1(n6342), 
	.B0(\ram[185][13] ), 
	.A1(n6362), 
	.A0(\ram[184][13] ));
   AOI22X1 U10910 (.Y(n13006), 
	.B1(n6381), 
	.B0(\ram[183][13] ), 
	.A1(n6400), 
	.A0(\ram[182][13] ));
   AOI22X1 U10911 (.Y(n13005), 
	.B1(n6419), 
	.B0(\ram[181][13] ), 
	.A1(n6438), 
	.A0(\ram[180][13] ));
   AOI22X1 U10912 (.Y(n13004), 
	.B1(n6457), 
	.B0(\ram[179][13] ), 
	.A1(n6476), 
	.A0(\ram[178][13] ));
   NAND4X1 U10913 (.Y(n13002), 
	.D(n13011), 
	.C(n13010), 
	.B(n13009), 
	.A(n13008));
   AOI22X1 U10914 (.Y(n13011), 
	.B1(n6495), 
	.B0(\ram[177][13] ), 
	.A1(n6514), 
	.A0(\ram[176][13] ));
   AOI22X1 U10915 (.Y(n13010), 
	.B1(n6533), 
	.B0(\ram[191][13] ), 
	.A1(n6553), 
	.A0(\ram[190][13] ));
   AOI22X1 U10916 (.Y(n13009), 
	.B1(n6572), 
	.B0(\ram[189][13] ), 
	.A1(n6591), 
	.A0(\ram[188][13] ));
   AOI22X1 U10917 (.Y(n13008), 
	.B1(n6610), 
	.B0(\ram[187][13] ), 
	.A1(n6629), 
	.A0(\ram[186][13] ));
   OAI21XL U10918 (.Y(n12989), 
	.B0(n8273), 
	.A1(n13013), 
	.A0(n13012));
   NAND4X1 U10919 (.Y(n13013), 
	.D(n13017), 
	.C(n13016), 
	.B(n13015), 
	.A(n13014));
   AOI22X1 U10920 (.Y(n13017), 
	.B1(n6342), 
	.B0(\ram[169][13] ), 
	.A1(n6362), 
	.A0(\ram[168][13] ));
   AOI22X1 U10921 (.Y(n13016), 
	.B1(n6381), 
	.B0(\ram[167][13] ), 
	.A1(n6400), 
	.A0(\ram[166][13] ));
   AOI22X1 U10922 (.Y(n13015), 
	.B1(n6419), 
	.B0(\ram[165][13] ), 
	.A1(n6438), 
	.A0(\ram[164][13] ));
   AOI22X1 U10923 (.Y(n13014), 
	.B1(n6457), 
	.B0(\ram[163][13] ), 
	.A1(n6476), 
	.A0(\ram[162][13] ));
   NAND4X1 U10924 (.Y(n13012), 
	.D(n13021), 
	.C(n13020), 
	.B(n13019), 
	.A(n13018));
   AOI22X1 U10925 (.Y(n13021), 
	.B1(n6495), 
	.B0(\ram[161][13] ), 
	.A1(n6514), 
	.A0(\ram[160][13] ));
   AOI22X1 U10926 (.Y(n13020), 
	.B1(n6533), 
	.B0(\ram[175][13] ), 
	.A1(n6553), 
	.A0(\ram[174][13] ));
   AOI22X1 U10927 (.Y(n13019), 
	.B1(n6572), 
	.B0(\ram[173][13] ), 
	.A1(n6591), 
	.A0(\ram[172][13] ));
   AOI22X1 U10928 (.Y(n13018), 
	.B1(n6610), 
	.B0(\ram[171][13] ), 
	.A1(n6629), 
	.A0(\ram[170][13] ));
   OAI21XL U10929 (.Y(n12988), 
	.B0(n8562), 
	.A1(n13023), 
	.A0(n13022));
   NAND4X1 U10930 (.Y(n13023), 
	.D(n13027), 
	.C(n13026), 
	.B(n13025), 
	.A(n13024));
   AOI22X1 U10931 (.Y(n13027), 
	.B1(n6342), 
	.B0(\ram[153][13] ), 
	.A1(n6362), 
	.A0(\ram[152][13] ));
   AOI22X1 U10932 (.Y(n13026), 
	.B1(n6381), 
	.B0(\ram[151][13] ), 
	.A1(n6400), 
	.A0(\ram[150][13] ));
   AOI22X1 U10933 (.Y(n13025), 
	.B1(n6419), 
	.B0(\ram[149][13] ), 
	.A1(n6438), 
	.A0(\ram[148][13] ));
   AOI22X1 U10934 (.Y(n13024), 
	.B1(n6457), 
	.B0(\ram[147][13] ), 
	.A1(n6476), 
	.A0(\ram[146][13] ));
   NAND4X1 U10935 (.Y(n13022), 
	.D(n13031), 
	.C(n13030), 
	.B(n13029), 
	.A(n13028));
   AOI22X1 U10936 (.Y(n13031), 
	.B1(n6495), 
	.B0(\ram[145][13] ), 
	.A1(n6514), 
	.A0(\ram[144][13] ));
   AOI22X1 U10937 (.Y(n13030), 
	.B1(n6533), 
	.B0(\ram[159][13] ), 
	.A1(n6553), 
	.A0(\ram[158][13] ));
   AOI22X1 U10938 (.Y(n13029), 
	.B1(n6572), 
	.B0(\ram[157][13] ), 
	.A1(n6591), 
	.A0(\ram[156][13] ));
   AOI22X1 U10939 (.Y(n13028), 
	.B1(n6610), 
	.B0(\ram[155][13] ), 
	.A1(n6629), 
	.A0(\ram[154][13] ));
   NAND4X1 U10940 (.Y(n12941), 
	.D(n13035), 
	.C(n13034), 
	.B(n13033), 
	.A(n13032));
   OAI21XL U10941 (.Y(n13035), 
	.B0(n8851), 
	.A1(n13037), 
	.A0(n13036));
   NAND4X1 U10942 (.Y(n13037), 
	.D(n13041), 
	.C(n13040), 
	.B(n13039), 
	.A(n13038));
   AOI22X1 U10943 (.Y(n13041), 
	.B1(n6342), 
	.B0(\ram[137][13] ), 
	.A1(n6362), 
	.A0(\ram[136][13] ));
   AOI22X1 U10944 (.Y(n13040), 
	.B1(n6381), 
	.B0(\ram[135][13] ), 
	.A1(n6400), 
	.A0(\ram[134][13] ));
   AOI22X1 U10945 (.Y(n13039), 
	.B1(n6419), 
	.B0(\ram[133][13] ), 
	.A1(n6438), 
	.A0(\ram[132][13] ));
   AOI22X1 U10946 (.Y(n13038), 
	.B1(n6457), 
	.B0(\ram[131][13] ), 
	.A1(n6476), 
	.A0(\ram[130][13] ));
   NAND4X1 U10947 (.Y(n13036), 
	.D(n13045), 
	.C(n13044), 
	.B(n13043), 
	.A(n13042));
   AOI22X1 U10948 (.Y(n13045), 
	.B1(n6495), 
	.B0(\ram[129][13] ), 
	.A1(n6514), 
	.A0(\ram[128][13] ));
   AOI22X1 U10949 (.Y(n13044), 
	.B1(n6533), 
	.B0(\ram[143][13] ), 
	.A1(n6553), 
	.A0(\ram[142][13] ));
   AOI22X1 U10950 (.Y(n13043), 
	.B1(n6572), 
	.B0(\ram[141][13] ), 
	.A1(n6591), 
	.A0(\ram[140][13] ));
   AOI22X1 U10951 (.Y(n13042), 
	.B1(n6610), 
	.B0(\ram[139][13] ), 
	.A1(n6629), 
	.A0(\ram[138][13] ));
   OAI21XL U10952 (.Y(n13034), 
	.B0(n9140), 
	.A1(n13047), 
	.A0(n13046));
   NAND4X1 U10953 (.Y(n13047), 
	.D(n13051), 
	.C(n13050), 
	.B(n13049), 
	.A(n13048));
   AOI22X1 U10954 (.Y(n13051), 
	.B1(n6342), 
	.B0(\ram[121][13] ), 
	.A1(n6362), 
	.A0(\ram[120][13] ));
   AOI22X1 U10955 (.Y(n13050), 
	.B1(n6381), 
	.B0(\ram[119][13] ), 
	.A1(n6400), 
	.A0(\ram[118][13] ));
   AOI22X1 U10956 (.Y(n13049), 
	.B1(n6419), 
	.B0(\ram[117][13] ), 
	.A1(n6438), 
	.A0(\ram[116][13] ));
   AOI22X1 U10957 (.Y(n13048), 
	.B1(n6457), 
	.B0(\ram[115][13] ), 
	.A1(n6476), 
	.A0(\ram[114][13] ));
   NAND4X1 U10958 (.Y(n13046), 
	.D(n13055), 
	.C(n13054), 
	.B(n13053), 
	.A(n13052));
   AOI22X1 U10959 (.Y(n13055), 
	.B1(n6495), 
	.B0(\ram[113][13] ), 
	.A1(n6514), 
	.A0(\ram[112][13] ));
   AOI22X1 U10960 (.Y(n13054), 
	.B1(n6533), 
	.B0(\ram[127][13] ), 
	.A1(n6553), 
	.A0(\ram[126][13] ));
   AOI22X1 U10961 (.Y(n13053), 
	.B1(n6572), 
	.B0(\ram[125][13] ), 
	.A1(n6591), 
	.A0(\ram[124][13] ));
   AOI22X1 U10962 (.Y(n13052), 
	.B1(n6610), 
	.B0(\ram[123][13] ), 
	.A1(n6629), 
	.A0(\ram[122][13] ));
   OAI21XL U10963 (.Y(n13033), 
	.B0(n9429), 
	.A1(n13057), 
	.A0(n13056));
   NAND4X1 U10964 (.Y(n13057), 
	.D(n13061), 
	.C(n13060), 
	.B(n13059), 
	.A(n13058));
   AOI22X1 U10965 (.Y(n13061), 
	.B1(n6342), 
	.B0(\ram[105][13] ), 
	.A1(n6362), 
	.A0(\ram[104][13] ));
   AOI22X1 U10966 (.Y(n13060), 
	.B1(n6381), 
	.B0(\ram[103][13] ), 
	.A1(n6400), 
	.A0(\ram[102][13] ));
   AOI22X1 U10967 (.Y(n13059), 
	.B1(n6419), 
	.B0(\ram[101][13] ), 
	.A1(n6438), 
	.A0(\ram[100][13] ));
   AOI22X1 U10968 (.Y(n13058), 
	.B1(n6457), 
	.B0(\ram[99][13] ), 
	.A1(n6476), 
	.A0(\ram[98][13] ));
   NAND4X1 U10969 (.Y(n13056), 
	.D(n13065), 
	.C(n13064), 
	.B(n13063), 
	.A(n13062));
   AOI22X1 U10970 (.Y(n13065), 
	.B1(n6495), 
	.B0(\ram[97][13] ), 
	.A1(n6514), 
	.A0(\ram[96][13] ));
   AOI22X1 U10971 (.Y(n13064), 
	.B1(n6533), 
	.B0(\ram[111][13] ), 
	.A1(n6553), 
	.A0(\ram[110][13] ));
   AOI22X1 U10972 (.Y(n13063), 
	.B1(n6572), 
	.B0(\ram[109][13] ), 
	.A1(n6591), 
	.A0(\ram[108][13] ));
   AOI22X1 U10973 (.Y(n13062), 
	.B1(n6610), 
	.B0(\ram[107][13] ), 
	.A1(n6629), 
	.A0(\ram[106][13] ));
   OAI21XL U10974 (.Y(n13032), 
	.B0(n9718), 
	.A1(n13067), 
	.A0(n13066));
   NAND4X1 U10975 (.Y(n13067), 
	.D(n13071), 
	.C(n13070), 
	.B(n13069), 
	.A(n13068));
   AOI22X1 U10976 (.Y(n13071), 
	.B1(n6342), 
	.B0(\ram[89][13] ), 
	.A1(n6362), 
	.A0(\ram[88][13] ));
   AOI22X1 U10977 (.Y(n13070), 
	.B1(n6381), 
	.B0(\ram[87][13] ), 
	.A1(n6400), 
	.A0(\ram[86][13] ));
   AOI22X1 U10978 (.Y(n13069), 
	.B1(n6419), 
	.B0(\ram[85][13] ), 
	.A1(n6438), 
	.A0(\ram[84][13] ));
   AOI22X1 U10979 (.Y(n13068), 
	.B1(n6457), 
	.B0(\ram[83][13] ), 
	.A1(n6476), 
	.A0(\ram[82][13] ));
   NAND4X1 U10980 (.Y(n13066), 
	.D(n13075), 
	.C(n13074), 
	.B(n13073), 
	.A(n13072));
   AOI22X1 U10981 (.Y(n13075), 
	.B1(n6495), 
	.B0(\ram[81][13] ), 
	.A1(n6514), 
	.A0(\ram[80][13] ));
   AOI22X1 U10982 (.Y(n13074), 
	.B1(n6533), 
	.B0(\ram[95][13] ), 
	.A1(n6553), 
	.A0(\ram[94][13] ));
   AOI22X1 U10983 (.Y(n13073), 
	.B1(n6572), 
	.B0(\ram[93][13] ), 
	.A1(n6591), 
	.A0(\ram[92][13] ));
   AOI22X1 U10984 (.Y(n13072), 
	.B1(n6610), 
	.B0(\ram[91][13] ), 
	.A1(n6629), 
	.A0(\ram[90][13] ));
   NAND4X1 U10985 (.Y(n12940), 
	.D(n13079), 
	.C(n13078), 
	.B(n13077), 
	.A(n13076));
   OAI21XL U10986 (.Y(n13079), 
	.B0(n10007), 
	.A1(n13081), 
	.A0(n13080));
   NAND4X1 U10987 (.Y(n13081), 
	.D(n13085), 
	.C(n13084), 
	.B(n13083), 
	.A(n13082));
   AOI22X1 U10988 (.Y(n13085), 
	.B1(n6342), 
	.B0(\ram[73][13] ), 
	.A1(n6362), 
	.A0(\ram[72][13] ));
   AOI22X1 U10989 (.Y(n13084), 
	.B1(n6381), 
	.B0(\ram[71][13] ), 
	.A1(n6400), 
	.A0(\ram[70][13] ));
   AOI22X1 U10990 (.Y(n13083), 
	.B1(n6419), 
	.B0(\ram[69][13] ), 
	.A1(n6438), 
	.A0(\ram[68][13] ));
   AOI22X1 U10991 (.Y(n13082), 
	.B1(n6457), 
	.B0(\ram[67][13] ), 
	.A1(n6476), 
	.A0(\ram[66][13] ));
   NAND4X1 U10992 (.Y(n13080), 
	.D(n13089), 
	.C(n13088), 
	.B(n13087), 
	.A(n13086));
   AOI22X1 U10993 (.Y(n13089), 
	.B1(n6495), 
	.B0(\ram[65][13] ), 
	.A1(n6514), 
	.A0(\ram[64][13] ));
   AOI22X1 U10994 (.Y(n13088), 
	.B1(n6533), 
	.B0(\ram[79][13] ), 
	.A1(n6553), 
	.A0(\ram[78][13] ));
   AOI22X1 U10995 (.Y(n13087), 
	.B1(n6572), 
	.B0(\ram[77][13] ), 
	.A1(n6591), 
	.A0(\ram[76][13] ));
   AOI22X1 U10996 (.Y(n13086), 
	.B1(n6610), 
	.B0(\ram[75][13] ), 
	.A1(n6629), 
	.A0(\ram[74][13] ));
   OAI21XL U10997 (.Y(n13078), 
	.B0(n10296), 
	.A1(n13091), 
	.A0(n13090));
   NAND4X1 U10998 (.Y(n13091), 
	.D(n13095), 
	.C(n13094), 
	.B(n13093), 
	.A(n13092));
   AOI22X1 U10999 (.Y(n13095), 
	.B1(n6342), 
	.B0(\ram[57][13] ), 
	.A1(n6362), 
	.A0(\ram[56][13] ));
   AOI22X1 U11000 (.Y(n13094), 
	.B1(n6381), 
	.B0(\ram[55][13] ), 
	.A1(n6400), 
	.A0(\ram[54][13] ));
   AOI22X1 U11001 (.Y(n13093), 
	.B1(n6419), 
	.B0(\ram[53][13] ), 
	.A1(n6438), 
	.A0(\ram[52][13] ));
   AOI22X1 U11002 (.Y(n13092), 
	.B1(n6457), 
	.B0(\ram[51][13] ), 
	.A1(n6476), 
	.A0(\ram[50][13] ));
   NAND4X1 U11003 (.Y(n13090), 
	.D(n13099), 
	.C(n13098), 
	.B(n13097), 
	.A(n13096));
   AOI22X1 U11004 (.Y(n13099), 
	.B1(n6495), 
	.B0(\ram[49][13] ), 
	.A1(n6514), 
	.A0(\ram[48][13] ));
   AOI22X1 U11005 (.Y(n13098), 
	.B1(n6533), 
	.B0(\ram[63][13] ), 
	.A1(n6553), 
	.A0(\ram[62][13] ));
   AOI22X1 U11006 (.Y(n13097), 
	.B1(n6572), 
	.B0(\ram[61][13] ), 
	.A1(n6591), 
	.A0(\ram[60][13] ));
   AOI22X1 U11007 (.Y(n13096), 
	.B1(n6610), 
	.B0(\ram[59][13] ), 
	.A1(n6629), 
	.A0(\ram[58][13] ));
   OAI21XL U11008 (.Y(n13077), 
	.B0(n10585), 
	.A1(n13101), 
	.A0(n13100));
   NAND4X1 U11009 (.Y(n13101), 
	.D(n13105), 
	.C(n13104), 
	.B(n13103), 
	.A(n13102));
   AOI22X1 U11010 (.Y(n13105), 
	.B1(n6342), 
	.B0(\ram[41][13] ), 
	.A1(n6362), 
	.A0(\ram[40][13] ));
   AOI22X1 U11011 (.Y(n13104), 
	.B1(n6381), 
	.B0(\ram[39][13] ), 
	.A1(n6400), 
	.A0(\ram[38][13] ));
   AOI22X1 U11012 (.Y(n13103), 
	.B1(n6419), 
	.B0(\ram[37][13] ), 
	.A1(n6438), 
	.A0(\ram[36][13] ));
   AOI22X1 U11013 (.Y(n13102), 
	.B1(n6457), 
	.B0(\ram[35][13] ), 
	.A1(n6476), 
	.A0(\ram[34][13] ));
   NAND4X1 U11014 (.Y(n13100), 
	.D(n13109), 
	.C(n13108), 
	.B(n13107), 
	.A(n13106));
   AOI22X1 U11015 (.Y(n13109), 
	.B1(n6495), 
	.B0(\ram[33][13] ), 
	.A1(n6514), 
	.A0(\ram[32][13] ));
   AOI22X1 U11016 (.Y(n13108), 
	.B1(n6533), 
	.B0(\ram[47][13] ), 
	.A1(n6553), 
	.A0(\ram[46][13] ));
   AOI22X1 U11017 (.Y(n13107), 
	.B1(n6572), 
	.B0(\ram[45][13] ), 
	.A1(n6591), 
	.A0(\ram[44][13] ));
   AOI22X1 U11018 (.Y(n13106), 
	.B1(n6610), 
	.B0(\ram[43][13] ), 
	.A1(n6629), 
	.A0(\ram[42][13] ));
   OAI21XL U11019 (.Y(n13076), 
	.B0(n6343), 
	.A1(n13111), 
	.A0(n13110));
   NAND4X1 U11020 (.Y(n13111), 
	.D(n13115), 
	.C(n13114), 
	.B(n13113), 
	.A(n13112));
   AOI22X1 U11021 (.Y(n13115), 
	.B1(n6342), 
	.B0(\ram[25][13] ), 
	.A1(n6362), 
	.A0(\ram[24][13] ));
   AOI22X1 U11022 (.Y(n13114), 
	.B1(n6381), 
	.B0(\ram[23][13] ), 
	.A1(n6400), 
	.A0(\ram[22][13] ));
   AOI22X1 U11023 (.Y(n13113), 
	.B1(n6419), 
	.B0(\ram[21][13] ), 
	.A1(n6438), 
	.A0(\ram[20][13] ));
   AOI22X1 U11024 (.Y(n13112), 
	.B1(n6457), 
	.B0(\ram[19][13] ), 
	.A1(n6476), 
	.A0(\ram[18][13] ));
   NAND4X1 U11025 (.Y(n13110), 
	.D(n13119), 
	.C(n13118), 
	.B(n13117), 
	.A(n13116));
   AOI22X1 U11026 (.Y(n13119), 
	.B1(n6495), 
	.B0(\ram[17][13] ), 
	.A1(n6514), 
	.A0(\ram[16][13] ));
   AOI22X1 U11027 (.Y(n13118), 
	.B1(n6533), 
	.B0(\ram[31][13] ), 
	.A1(n6553), 
	.A0(\ram[30][13] ));
   AOI22X1 U11028 (.Y(n13117), 
	.B1(n6572), 
	.B0(\ram[29][13] ), 
	.A1(n6591), 
	.A0(\ram[28][13] ));
   AOI22X1 U11029 (.Y(n13116), 
	.B1(n6610), 
	.B0(\ram[27][13] ), 
	.A1(n6629), 
	.A0(\ram[26][13] ));
   OR4X1 U11030 (.Y(mem_read_data[12]), 
	.D(n13123), 
	.C(n13122), 
	.B(n13121), 
	.A(n13120));
   NAND4X1 U11031 (.Y(n13123), 
	.D(n13127), 
	.C(n13126), 
	.B(n13125), 
	.A(n13124));
   OAI21XL U11032 (.Y(n13127), 
	.B0(n6534), 
	.A1(n13129), 
	.A0(n13128));
   NAND4X1 U11033 (.Y(n13129), 
	.D(n13133), 
	.C(n13132), 
	.B(n13131), 
	.A(n13130));
   AOI22X1 U11034 (.Y(n13133), 
	.B1(n6342), 
	.B0(\ram[9][12] ), 
	.A1(n6362), 
	.A0(\ram[8][12] ));
   AOI22X1 U11035 (.Y(n13132), 
	.B1(n6381), 
	.B0(\ram[7][12] ), 
	.A1(n6400), 
	.A0(\ram[6][12] ));
   AOI22X1 U11036 (.Y(n13131), 
	.B1(n6419), 
	.B0(\ram[5][12] ), 
	.A1(n6438), 
	.A0(\ram[4][12] ));
   AOI22X1 U11037 (.Y(n13130), 
	.B1(n6457), 
	.B0(\ram[3][12] ), 
	.A1(n6476), 
	.A0(\ram[2][12] ));
   NAND4X1 U11038 (.Y(n13128), 
	.D(n13137), 
	.C(n13136), 
	.B(n13135), 
	.A(n13134));
   AOI22X1 U11039 (.Y(n13137), 
	.B1(n6495), 
	.B0(\ram[1][12] ), 
	.A1(n6514), 
	.A0(\ram[0][12] ));
   AOI22X1 U11040 (.Y(n13136), 
	.B1(n6533), 
	.B0(\ram[15][12] ), 
	.A1(n6553), 
	.A0(\ram[14][12] ));
   AOI22X1 U11041 (.Y(n13135), 
	.B1(n6572), 
	.B0(\ram[13][12] ), 
	.A1(n6591), 
	.A0(\ram[12][12] ));
   AOI22X1 U11042 (.Y(n13134), 
	.B1(n6610), 
	.B0(\ram[11][12] ), 
	.A1(n6629), 
	.A0(\ram[10][12] ));
   OAI21XL U11043 (.Y(n13126), 
	.B0(n6828), 
	.A1(n13139), 
	.A0(n13138));
   NAND4X1 U11044 (.Y(n13139), 
	.D(n13143), 
	.C(n13142), 
	.B(n13141), 
	.A(n13140));
   AOI22X1 U11045 (.Y(n13143), 
	.B1(n6342), 
	.B0(\ram[249][12] ), 
	.A1(n6362), 
	.A0(\ram[248][12] ));
   AOI22X1 U11046 (.Y(n13142), 
	.B1(n6381), 
	.B0(\ram[247][12] ), 
	.A1(n6400), 
	.A0(\ram[246][12] ));
   AOI22X1 U11047 (.Y(n13141), 
	.B1(n6419), 
	.B0(\ram[245][12] ), 
	.A1(n6438), 
	.A0(\ram[244][12] ));
   AOI22X1 U11048 (.Y(n13140), 
	.B1(n6457), 
	.B0(\ram[243][12] ), 
	.A1(n6476), 
	.A0(\ram[242][12] ));
   NAND4X1 U11049 (.Y(n13138), 
	.D(n13147), 
	.C(n13146), 
	.B(n13145), 
	.A(n13144));
   AOI22X1 U11050 (.Y(n13147), 
	.B1(n6495), 
	.B0(\ram[241][12] ), 
	.A1(n6514), 
	.A0(\ram[240][12] ));
   AOI22X1 U11051 (.Y(n13146), 
	.B1(n6533), 
	.B0(\ram[255][12] ), 
	.A1(n6553), 
	.A0(\ram[254][12] ));
   AOI22X1 U11052 (.Y(n13145), 
	.B1(n6572), 
	.B0(\ram[253][12] ), 
	.A1(n6591), 
	.A0(\ram[252][12] ));
   AOI22X1 U11053 (.Y(n13144), 
	.B1(n6610), 
	.B0(\ram[251][12] ), 
	.A1(n6629), 
	.A0(\ram[250][12] ));
   OAI21XL U11054 (.Y(n13125), 
	.B0(n7117), 
	.A1(n13149), 
	.A0(n13148));
   NAND4X1 U11055 (.Y(n13149), 
	.D(n13153), 
	.C(n13152), 
	.B(n13151), 
	.A(n13150));
   AOI22X1 U11056 (.Y(n13153), 
	.B1(n6342), 
	.B0(\ram[233][12] ), 
	.A1(n6362), 
	.A0(\ram[232][12] ));
   AOI22X1 U11057 (.Y(n13152), 
	.B1(n6381), 
	.B0(\ram[231][12] ), 
	.A1(n6400), 
	.A0(\ram[230][12] ));
   AOI22X1 U11058 (.Y(n13151), 
	.B1(n6419), 
	.B0(\ram[229][12] ), 
	.A1(n6438), 
	.A0(\ram[228][12] ));
   AOI22X1 U11059 (.Y(n13150), 
	.B1(n6457), 
	.B0(\ram[227][12] ), 
	.A1(n6476), 
	.A0(\ram[226][12] ));
   NAND4X1 U11060 (.Y(n13148), 
	.D(n13157), 
	.C(n13156), 
	.B(n13155), 
	.A(n13154));
   AOI22X1 U11061 (.Y(n13157), 
	.B1(n6495), 
	.B0(\ram[225][12] ), 
	.A1(n6514), 
	.A0(\ram[224][12] ));
   AOI22X1 U11062 (.Y(n13156), 
	.B1(n6533), 
	.B0(\ram[239][12] ), 
	.A1(n6553), 
	.A0(\ram[238][12] ));
   AOI22X1 U11063 (.Y(n13155), 
	.B1(n6572), 
	.B0(\ram[237][12] ), 
	.A1(n6591), 
	.A0(\ram[236][12] ));
   AOI22X1 U11064 (.Y(n13154), 
	.B1(n6610), 
	.B0(\ram[235][12] ), 
	.A1(n6629), 
	.A0(\ram[234][12] ));
   OAI21XL U11065 (.Y(n13124), 
	.B0(n7406), 
	.A1(n13159), 
	.A0(n13158));
   NAND4X1 U11066 (.Y(n13159), 
	.D(n13163), 
	.C(n13162), 
	.B(n13161), 
	.A(n13160));
   AOI22X1 U11067 (.Y(n13163), 
	.B1(n6342), 
	.B0(\ram[217][12] ), 
	.A1(n6362), 
	.A0(\ram[216][12] ));
   AOI22X1 U11068 (.Y(n13162), 
	.B1(n6381), 
	.B0(\ram[215][12] ), 
	.A1(n6400), 
	.A0(\ram[214][12] ));
   AOI22X1 U11069 (.Y(n13161), 
	.B1(n6419), 
	.B0(\ram[213][12] ), 
	.A1(n6438), 
	.A0(\ram[212][12] ));
   AOI22X1 U11070 (.Y(n13160), 
	.B1(n6457), 
	.B0(\ram[211][12] ), 
	.A1(n6476), 
	.A0(\ram[210][12] ));
   NAND4X1 U11071 (.Y(n13158), 
	.D(n13167), 
	.C(n13166), 
	.B(n13165), 
	.A(n13164));
   AOI22X1 U11072 (.Y(n13167), 
	.B1(n6495), 
	.B0(\ram[209][12] ), 
	.A1(n6514), 
	.A0(\ram[208][12] ));
   AOI22X1 U11073 (.Y(n13166), 
	.B1(n6533), 
	.B0(\ram[223][12] ), 
	.A1(n6553), 
	.A0(\ram[222][12] ));
   AOI22X1 U11074 (.Y(n13165), 
	.B1(n6572), 
	.B0(\ram[221][12] ), 
	.A1(n6591), 
	.A0(\ram[220][12] ));
   AOI22X1 U11075 (.Y(n13164), 
	.B1(n6610), 
	.B0(\ram[219][12] ), 
	.A1(n6629), 
	.A0(\ram[218][12] ));
   NAND4X1 U11076 (.Y(n13122), 
	.D(n13171), 
	.C(n13170), 
	.B(n13169), 
	.A(n13168));
   OAI21XL U11077 (.Y(n13171), 
	.B0(n7695), 
	.A1(n13173), 
	.A0(n13172));
   NAND4X1 U11078 (.Y(n13173), 
	.D(n13177), 
	.C(n13176), 
	.B(n13175), 
	.A(n13174));
   AOI22X1 U11079 (.Y(n13177), 
	.B1(n6342), 
	.B0(\ram[201][12] ), 
	.A1(n6362), 
	.A0(\ram[200][12] ));
   AOI22X1 U11080 (.Y(n13176), 
	.B1(n6381), 
	.B0(\ram[199][12] ), 
	.A1(n6400), 
	.A0(\ram[198][12] ));
   AOI22X1 U11081 (.Y(n13175), 
	.B1(n6419), 
	.B0(\ram[197][12] ), 
	.A1(n6438), 
	.A0(\ram[196][12] ));
   AOI22X1 U11082 (.Y(n13174), 
	.B1(n6457), 
	.B0(\ram[195][12] ), 
	.A1(n6476), 
	.A0(\ram[194][12] ));
   NAND4X1 U11083 (.Y(n13172), 
	.D(n13181), 
	.C(n13180), 
	.B(n13179), 
	.A(n13178));
   AOI22X1 U11084 (.Y(n13181), 
	.B1(n6495), 
	.B0(\ram[193][12] ), 
	.A1(n6514), 
	.A0(\ram[192][12] ));
   AOI22X1 U11085 (.Y(n13180), 
	.B1(n6533), 
	.B0(\ram[207][12] ), 
	.A1(n6553), 
	.A0(\ram[206][12] ));
   AOI22X1 U11086 (.Y(n13179), 
	.B1(n6572), 
	.B0(\ram[205][12] ), 
	.A1(n6591), 
	.A0(\ram[204][12] ));
   AOI22X1 U11087 (.Y(n13178), 
	.B1(n6610), 
	.B0(\ram[203][12] ), 
	.A1(n6629), 
	.A0(\ram[202][12] ));
   OAI21XL U11088 (.Y(n13170), 
	.B0(n7984), 
	.A1(n13183), 
	.A0(n13182));
   NAND4X1 U11089 (.Y(n13183), 
	.D(n13187), 
	.C(n13186), 
	.B(n13185), 
	.A(n13184));
   AOI22X1 U11090 (.Y(n13187), 
	.B1(n6342), 
	.B0(\ram[185][12] ), 
	.A1(n6362), 
	.A0(\ram[184][12] ));
   AOI22X1 U11091 (.Y(n13186), 
	.B1(n6381), 
	.B0(\ram[183][12] ), 
	.A1(n6400), 
	.A0(\ram[182][12] ));
   AOI22X1 U11092 (.Y(n13185), 
	.B1(n6419), 
	.B0(\ram[181][12] ), 
	.A1(n6438), 
	.A0(\ram[180][12] ));
   AOI22X1 U11093 (.Y(n13184), 
	.B1(n6457), 
	.B0(\ram[179][12] ), 
	.A1(n6476), 
	.A0(\ram[178][12] ));
   NAND4X1 U11094 (.Y(n13182), 
	.D(n13191), 
	.C(n13190), 
	.B(n13189), 
	.A(n13188));
   AOI22X1 U11095 (.Y(n13191), 
	.B1(n6495), 
	.B0(\ram[177][12] ), 
	.A1(n6514), 
	.A0(\ram[176][12] ));
   AOI22X1 U11096 (.Y(n13190), 
	.B1(n6533), 
	.B0(\ram[191][12] ), 
	.A1(n6553), 
	.A0(\ram[190][12] ));
   AOI22X1 U11097 (.Y(n13189), 
	.B1(n6572), 
	.B0(\ram[189][12] ), 
	.A1(n6591), 
	.A0(\ram[188][12] ));
   AOI22X1 U11098 (.Y(n13188), 
	.B1(n6610), 
	.B0(\ram[187][12] ), 
	.A1(n6629), 
	.A0(\ram[186][12] ));
   OAI21XL U11099 (.Y(n13169), 
	.B0(n8273), 
	.A1(n13193), 
	.A0(n13192));
   NAND4X1 U11100 (.Y(n13193), 
	.D(n13197), 
	.C(n13196), 
	.B(n13195), 
	.A(n13194));
   AOI22X1 U11101 (.Y(n13197), 
	.B1(n6342), 
	.B0(\ram[169][12] ), 
	.A1(n6362), 
	.A0(\ram[168][12] ));
   AOI22X1 U11102 (.Y(n13196), 
	.B1(n6381), 
	.B0(\ram[167][12] ), 
	.A1(n6400), 
	.A0(\ram[166][12] ));
   AOI22X1 U11103 (.Y(n13195), 
	.B1(n6419), 
	.B0(\ram[165][12] ), 
	.A1(n6438), 
	.A0(\ram[164][12] ));
   AOI22X1 U11104 (.Y(n13194), 
	.B1(n6457), 
	.B0(\ram[163][12] ), 
	.A1(n6476), 
	.A0(\ram[162][12] ));
   NAND4X1 U11105 (.Y(n13192), 
	.D(n13201), 
	.C(n13200), 
	.B(n13199), 
	.A(n13198));
   AOI22X1 U11106 (.Y(n13201), 
	.B1(n6495), 
	.B0(\ram[161][12] ), 
	.A1(n6514), 
	.A0(\ram[160][12] ));
   AOI22X1 U11107 (.Y(n13200), 
	.B1(n6533), 
	.B0(\ram[175][12] ), 
	.A1(n6553), 
	.A0(\ram[174][12] ));
   AOI22X1 U11108 (.Y(n13199), 
	.B1(n6572), 
	.B0(\ram[173][12] ), 
	.A1(n6591), 
	.A0(\ram[172][12] ));
   AOI22X1 U11109 (.Y(n13198), 
	.B1(n6610), 
	.B0(\ram[171][12] ), 
	.A1(n6629), 
	.A0(\ram[170][12] ));
   OAI21XL U11110 (.Y(n13168), 
	.B0(n8562), 
	.A1(n13203), 
	.A0(n13202));
   NAND4X1 U11111 (.Y(n13203), 
	.D(n13207), 
	.C(n13206), 
	.B(n13205), 
	.A(n13204));
   AOI22X1 U11112 (.Y(n13207), 
	.B1(n6342), 
	.B0(\ram[153][12] ), 
	.A1(n6362), 
	.A0(\ram[152][12] ));
   AOI22X1 U11113 (.Y(n13206), 
	.B1(n6381), 
	.B0(\ram[151][12] ), 
	.A1(n6400), 
	.A0(\ram[150][12] ));
   AOI22X1 U11114 (.Y(n13205), 
	.B1(n6419), 
	.B0(\ram[149][12] ), 
	.A1(n6438), 
	.A0(\ram[148][12] ));
   AOI22X1 U11115 (.Y(n13204), 
	.B1(n6457), 
	.B0(\ram[147][12] ), 
	.A1(n6476), 
	.A0(\ram[146][12] ));
   NAND4X1 U11116 (.Y(n13202), 
	.D(n13211), 
	.C(n13210), 
	.B(n13209), 
	.A(n13208));
   AOI22X1 U11117 (.Y(n13211), 
	.B1(n6495), 
	.B0(\ram[145][12] ), 
	.A1(n6514), 
	.A0(\ram[144][12] ));
   AOI22X1 U11118 (.Y(n13210), 
	.B1(n6533), 
	.B0(\ram[159][12] ), 
	.A1(n6553), 
	.A0(\ram[158][12] ));
   AOI22X1 U11119 (.Y(n13209), 
	.B1(n6572), 
	.B0(\ram[157][12] ), 
	.A1(n6591), 
	.A0(\ram[156][12] ));
   AOI22X1 U11120 (.Y(n13208), 
	.B1(n6610), 
	.B0(\ram[155][12] ), 
	.A1(n6629), 
	.A0(\ram[154][12] ));
   NAND4X1 U11121 (.Y(n13121), 
	.D(n13215), 
	.C(n13214), 
	.B(n13213), 
	.A(n13212));
   OAI21XL U11122 (.Y(n13215), 
	.B0(n8851), 
	.A1(n13217), 
	.A0(n13216));
   NAND4X1 U11123 (.Y(n13217), 
	.D(n13221), 
	.C(n13220), 
	.B(n13219), 
	.A(n13218));
   AOI22X1 U11124 (.Y(n13221), 
	.B1(n6342), 
	.B0(\ram[137][12] ), 
	.A1(n6362), 
	.A0(\ram[136][12] ));
   AOI22X1 U11125 (.Y(n13220), 
	.B1(n6381), 
	.B0(\ram[135][12] ), 
	.A1(n6400), 
	.A0(\ram[134][12] ));
   AOI22X1 U11126 (.Y(n13219), 
	.B1(n6419), 
	.B0(\ram[133][12] ), 
	.A1(n6438), 
	.A0(\ram[132][12] ));
   AOI22X1 U11127 (.Y(n13218), 
	.B1(n6457), 
	.B0(\ram[131][12] ), 
	.A1(n6476), 
	.A0(\ram[130][12] ));
   NAND4X1 U11128 (.Y(n13216), 
	.D(n13225), 
	.C(n13224), 
	.B(n13223), 
	.A(n13222));
   AOI22X1 U11129 (.Y(n13225), 
	.B1(n6495), 
	.B0(\ram[129][12] ), 
	.A1(n6514), 
	.A0(\ram[128][12] ));
   AOI22X1 U11130 (.Y(n13224), 
	.B1(n6533), 
	.B0(\ram[143][12] ), 
	.A1(n6553), 
	.A0(\ram[142][12] ));
   AOI22X1 U11131 (.Y(n13223), 
	.B1(n6572), 
	.B0(\ram[141][12] ), 
	.A1(n6591), 
	.A0(\ram[140][12] ));
   AOI22X1 U11132 (.Y(n13222), 
	.B1(n6610), 
	.B0(\ram[139][12] ), 
	.A1(n6629), 
	.A0(\ram[138][12] ));
   OAI21XL U11133 (.Y(n13214), 
	.B0(n9140), 
	.A1(n13227), 
	.A0(n13226));
   NAND4X1 U11134 (.Y(n13227), 
	.D(n13231), 
	.C(n13230), 
	.B(n13229), 
	.A(n13228));
   AOI22X1 U11135 (.Y(n13231), 
	.B1(n6342), 
	.B0(\ram[121][12] ), 
	.A1(n6362), 
	.A0(\ram[120][12] ));
   AOI22X1 U11136 (.Y(n13230), 
	.B1(n6381), 
	.B0(\ram[119][12] ), 
	.A1(n6400), 
	.A0(\ram[118][12] ));
   AOI22X1 U11137 (.Y(n13229), 
	.B1(n6419), 
	.B0(\ram[117][12] ), 
	.A1(n6438), 
	.A0(\ram[116][12] ));
   AOI22X1 U11138 (.Y(n13228), 
	.B1(n6457), 
	.B0(\ram[115][12] ), 
	.A1(n6476), 
	.A0(\ram[114][12] ));
   NAND4X1 U11139 (.Y(n13226), 
	.D(n13235), 
	.C(n13234), 
	.B(n13233), 
	.A(n13232));
   AOI22X1 U11140 (.Y(n13235), 
	.B1(n6495), 
	.B0(\ram[113][12] ), 
	.A1(n6514), 
	.A0(\ram[112][12] ));
   AOI22X1 U11141 (.Y(n13234), 
	.B1(n6533), 
	.B0(\ram[127][12] ), 
	.A1(n6553), 
	.A0(\ram[126][12] ));
   AOI22X1 U11142 (.Y(n13233), 
	.B1(n6572), 
	.B0(\ram[125][12] ), 
	.A1(n6591), 
	.A0(\ram[124][12] ));
   AOI22X1 U11143 (.Y(n13232), 
	.B1(n6610), 
	.B0(\ram[123][12] ), 
	.A1(n6629), 
	.A0(\ram[122][12] ));
   OAI21XL U11144 (.Y(n13213), 
	.B0(n9429), 
	.A1(n13237), 
	.A0(n13236));
   NAND4X1 U11145 (.Y(n13237), 
	.D(n13241), 
	.C(n13240), 
	.B(n13239), 
	.A(n13238));
   AOI22X1 U11146 (.Y(n13241), 
	.B1(n6342), 
	.B0(\ram[105][12] ), 
	.A1(n6362), 
	.A0(\ram[104][12] ));
   AOI22X1 U11147 (.Y(n13240), 
	.B1(n6381), 
	.B0(\ram[103][12] ), 
	.A1(n6400), 
	.A0(\ram[102][12] ));
   AOI22X1 U11148 (.Y(n13239), 
	.B1(n6419), 
	.B0(\ram[101][12] ), 
	.A1(n6438), 
	.A0(\ram[100][12] ));
   AOI22X1 U11149 (.Y(n13238), 
	.B1(n6457), 
	.B0(\ram[99][12] ), 
	.A1(n6476), 
	.A0(\ram[98][12] ));
   NAND4X1 U11150 (.Y(n13236), 
	.D(n13245), 
	.C(n13244), 
	.B(n13243), 
	.A(n13242));
   AOI22X1 U11151 (.Y(n13245), 
	.B1(n6495), 
	.B0(\ram[97][12] ), 
	.A1(n6514), 
	.A0(\ram[96][12] ));
   AOI22X1 U11152 (.Y(n13244), 
	.B1(n6533), 
	.B0(\ram[111][12] ), 
	.A1(n6553), 
	.A0(\ram[110][12] ));
   AOI22X1 U11153 (.Y(n13243), 
	.B1(n6572), 
	.B0(\ram[109][12] ), 
	.A1(n6591), 
	.A0(\ram[108][12] ));
   AOI22X1 U11154 (.Y(n13242), 
	.B1(n6610), 
	.B0(\ram[107][12] ), 
	.A1(n6629), 
	.A0(\ram[106][12] ));
   OAI21XL U11155 (.Y(n13212), 
	.B0(n9718), 
	.A1(n13247), 
	.A0(n13246));
   NAND4X1 U11156 (.Y(n13247), 
	.D(n13251), 
	.C(n13250), 
	.B(n13249), 
	.A(n13248));
   AOI22X1 U11157 (.Y(n13251), 
	.B1(n6342), 
	.B0(\ram[89][12] ), 
	.A1(n6362), 
	.A0(\ram[88][12] ));
   AOI22X1 U11158 (.Y(n13250), 
	.B1(n6381), 
	.B0(\ram[87][12] ), 
	.A1(n6400), 
	.A0(\ram[86][12] ));
   AOI22X1 U11159 (.Y(n13249), 
	.B1(n6419), 
	.B0(\ram[85][12] ), 
	.A1(n6438), 
	.A0(\ram[84][12] ));
   AOI22X1 U11160 (.Y(n13248), 
	.B1(n6457), 
	.B0(\ram[83][12] ), 
	.A1(n6476), 
	.A0(\ram[82][12] ));
   NAND4X1 U11161 (.Y(n13246), 
	.D(n13255), 
	.C(n13254), 
	.B(n13253), 
	.A(n13252));
   AOI22X1 U11162 (.Y(n13255), 
	.B1(n6495), 
	.B0(\ram[81][12] ), 
	.A1(n6514), 
	.A0(\ram[80][12] ));
   AOI22X1 U11163 (.Y(n13254), 
	.B1(n6533), 
	.B0(\ram[95][12] ), 
	.A1(n6553), 
	.A0(\ram[94][12] ));
   AOI22X1 U11164 (.Y(n13253), 
	.B1(n6572), 
	.B0(\ram[93][12] ), 
	.A1(n6591), 
	.A0(\ram[92][12] ));
   AOI22X1 U11165 (.Y(n13252), 
	.B1(n6610), 
	.B0(\ram[91][12] ), 
	.A1(n6629), 
	.A0(\ram[90][12] ));
   NAND4X1 U11166 (.Y(n13120), 
	.D(n13259), 
	.C(n13258), 
	.B(n13257), 
	.A(n13256));
   OAI21XL U11167 (.Y(n13259), 
	.B0(n10007), 
	.A1(n13261), 
	.A0(n13260));
   NAND4X1 U11168 (.Y(n13261), 
	.D(n13265), 
	.C(n13264), 
	.B(n13263), 
	.A(n13262));
   AOI22X1 U11169 (.Y(n13265), 
	.B1(n6342), 
	.B0(\ram[73][12] ), 
	.A1(n6362), 
	.A0(\ram[72][12] ));
   AOI22X1 U11170 (.Y(n13264), 
	.B1(n6381), 
	.B0(\ram[71][12] ), 
	.A1(n6400), 
	.A0(\ram[70][12] ));
   AOI22X1 U11171 (.Y(n13263), 
	.B1(n6419), 
	.B0(\ram[69][12] ), 
	.A1(n6438), 
	.A0(\ram[68][12] ));
   AOI22X1 U11172 (.Y(n13262), 
	.B1(n6457), 
	.B0(\ram[67][12] ), 
	.A1(n6476), 
	.A0(\ram[66][12] ));
   NAND4X1 U11173 (.Y(n13260), 
	.D(n13269), 
	.C(n13268), 
	.B(n13267), 
	.A(n13266));
   AOI22X1 U11174 (.Y(n13269), 
	.B1(n6495), 
	.B0(\ram[65][12] ), 
	.A1(n6514), 
	.A0(\ram[64][12] ));
   AOI22X1 U11175 (.Y(n13268), 
	.B1(n6533), 
	.B0(\ram[79][12] ), 
	.A1(n6553), 
	.A0(\ram[78][12] ));
   AOI22X1 U11176 (.Y(n13267), 
	.B1(n6572), 
	.B0(\ram[77][12] ), 
	.A1(n6591), 
	.A0(\ram[76][12] ));
   AOI22X1 U11177 (.Y(n13266), 
	.B1(n6610), 
	.B0(\ram[75][12] ), 
	.A1(n6629), 
	.A0(\ram[74][12] ));
   OAI21XL U11178 (.Y(n13258), 
	.B0(n10296), 
	.A1(n13271), 
	.A0(n13270));
   NAND4X1 U11179 (.Y(n13271), 
	.D(n13275), 
	.C(n13274), 
	.B(n13273), 
	.A(n13272));
   AOI22X1 U11180 (.Y(n13275), 
	.B1(n6342), 
	.B0(\ram[57][12] ), 
	.A1(n6362), 
	.A0(\ram[56][12] ));
   AOI22X1 U11181 (.Y(n13274), 
	.B1(n6381), 
	.B0(\ram[55][12] ), 
	.A1(n6400), 
	.A0(\ram[54][12] ));
   AOI22X1 U11182 (.Y(n13273), 
	.B1(n6419), 
	.B0(\ram[53][12] ), 
	.A1(n6438), 
	.A0(\ram[52][12] ));
   AOI22X1 U11183 (.Y(n13272), 
	.B1(n6457), 
	.B0(\ram[51][12] ), 
	.A1(n6476), 
	.A0(\ram[50][12] ));
   NAND4X1 U11184 (.Y(n13270), 
	.D(n13279), 
	.C(n13278), 
	.B(n13277), 
	.A(n13276));
   AOI22X1 U11185 (.Y(n13279), 
	.B1(n6495), 
	.B0(\ram[49][12] ), 
	.A1(n6514), 
	.A0(\ram[48][12] ));
   AOI22X1 U11186 (.Y(n13278), 
	.B1(n6533), 
	.B0(\ram[63][12] ), 
	.A1(n6553), 
	.A0(\ram[62][12] ));
   AOI22X1 U11187 (.Y(n13277), 
	.B1(n6572), 
	.B0(\ram[61][12] ), 
	.A1(n6591), 
	.A0(\ram[60][12] ));
   AOI22X1 U11188 (.Y(n13276), 
	.B1(n6610), 
	.B0(\ram[59][12] ), 
	.A1(n6629), 
	.A0(\ram[58][12] ));
   OAI21XL U11189 (.Y(n13257), 
	.B0(n10585), 
	.A1(n13281), 
	.A0(n13280));
   NAND4X1 U11190 (.Y(n13281), 
	.D(n13285), 
	.C(n13284), 
	.B(n13283), 
	.A(n13282));
   AOI22X1 U11191 (.Y(n13285), 
	.B1(n6342), 
	.B0(\ram[41][12] ), 
	.A1(n6362), 
	.A0(\ram[40][12] ));
   AOI22X1 U11192 (.Y(n13284), 
	.B1(n6381), 
	.B0(\ram[39][12] ), 
	.A1(n6400), 
	.A0(\ram[38][12] ));
   AOI22X1 U11193 (.Y(n13283), 
	.B1(n6419), 
	.B0(\ram[37][12] ), 
	.A1(n6438), 
	.A0(\ram[36][12] ));
   AOI22X1 U11194 (.Y(n13282), 
	.B1(n6457), 
	.B0(\ram[35][12] ), 
	.A1(n6476), 
	.A0(\ram[34][12] ));
   NAND4X1 U11195 (.Y(n13280), 
	.D(n13289), 
	.C(n13288), 
	.B(n13287), 
	.A(n13286));
   AOI22X1 U11196 (.Y(n13289), 
	.B1(n6495), 
	.B0(\ram[33][12] ), 
	.A1(n6514), 
	.A0(\ram[32][12] ));
   AOI22X1 U11197 (.Y(n13288), 
	.B1(n6533), 
	.B0(\ram[47][12] ), 
	.A1(n6553), 
	.A0(\ram[46][12] ));
   AOI22X1 U11198 (.Y(n13287), 
	.B1(n6572), 
	.B0(\ram[45][12] ), 
	.A1(n6591), 
	.A0(\ram[44][12] ));
   AOI22X1 U11199 (.Y(n13286), 
	.B1(n6610), 
	.B0(\ram[43][12] ), 
	.A1(n6629), 
	.A0(\ram[42][12] ));
   OAI21XL U11200 (.Y(n13256), 
	.B0(n6343), 
	.A1(n13291), 
	.A0(n13290));
   NAND4X1 U11201 (.Y(n13291), 
	.D(n13295), 
	.C(n13294), 
	.B(n13293), 
	.A(n13292));
   AOI22X1 U11202 (.Y(n13295), 
	.B1(n6342), 
	.B0(\ram[25][12] ), 
	.A1(n6362), 
	.A0(\ram[24][12] ));
   AOI22X1 U11203 (.Y(n13294), 
	.B1(n6381), 
	.B0(\ram[23][12] ), 
	.A1(n6400), 
	.A0(\ram[22][12] ));
   AOI22X1 U11204 (.Y(n13293), 
	.B1(n6419), 
	.B0(\ram[21][12] ), 
	.A1(n6438), 
	.A0(\ram[20][12] ));
   AOI22X1 U11205 (.Y(n13292), 
	.B1(n6457), 
	.B0(\ram[19][12] ), 
	.A1(n6476), 
	.A0(\ram[18][12] ));
   NAND4X1 U11206 (.Y(n13290), 
	.D(n13299), 
	.C(n13298), 
	.B(n13297), 
	.A(n13296));
   AOI22X1 U11207 (.Y(n13299), 
	.B1(n6495), 
	.B0(\ram[17][12] ), 
	.A1(n6514), 
	.A0(\ram[16][12] ));
   AOI22X1 U11208 (.Y(n13298), 
	.B1(n6533), 
	.B0(\ram[31][12] ), 
	.A1(n6553), 
	.A0(\ram[30][12] ));
   AOI22X1 U11209 (.Y(n13297), 
	.B1(n6572), 
	.B0(\ram[29][12] ), 
	.A1(n6591), 
	.A0(\ram[28][12] ));
   AOI22X1 U11210 (.Y(n13296), 
	.B1(n6610), 
	.B0(\ram[27][12] ), 
	.A1(n6629), 
	.A0(\ram[26][12] ));
   OR4X1 U11211 (.Y(mem_read_data[11]), 
	.D(n13303), 
	.C(n13302), 
	.B(n13301), 
	.A(n13300));
   NAND4X1 U11212 (.Y(n13303), 
	.D(n13307), 
	.C(n13306), 
	.B(n13305), 
	.A(n13304));
   OAI21XL U11213 (.Y(n13307), 
	.B0(n6534), 
	.A1(n13309), 
	.A0(n13308));
   NAND4X1 U11214 (.Y(n13309), 
	.D(n13313), 
	.C(n13312), 
	.B(n13311), 
	.A(n13310));
   AOI22X1 U11215 (.Y(n13313), 
	.B1(n6342), 
	.B0(\ram[9][11] ), 
	.A1(n6362), 
	.A0(\ram[8][11] ));
   AOI22X1 U11216 (.Y(n13312), 
	.B1(n6381), 
	.B0(\ram[7][11] ), 
	.A1(n6400), 
	.A0(\ram[6][11] ));
   AOI22X1 U11217 (.Y(n13311), 
	.B1(n6419), 
	.B0(\ram[5][11] ), 
	.A1(n6438), 
	.A0(\ram[4][11] ));
   AOI22X1 U11218 (.Y(n13310), 
	.B1(n6457), 
	.B0(\ram[3][11] ), 
	.A1(n6476), 
	.A0(\ram[2][11] ));
   NAND4X1 U11219 (.Y(n13308), 
	.D(n13317), 
	.C(n13316), 
	.B(n13315), 
	.A(n13314));
   AOI22X1 U11220 (.Y(n13317), 
	.B1(n6495), 
	.B0(\ram[1][11] ), 
	.A1(n6514), 
	.A0(\ram[0][11] ));
   AOI22X1 U11221 (.Y(n13316), 
	.B1(n6533), 
	.B0(\ram[15][11] ), 
	.A1(n6553), 
	.A0(\ram[14][11] ));
   AOI22X1 U11222 (.Y(n13315), 
	.B1(n6572), 
	.B0(\ram[13][11] ), 
	.A1(n6591), 
	.A0(\ram[12][11] ));
   AOI22X1 U11223 (.Y(n13314), 
	.B1(n6610), 
	.B0(\ram[11][11] ), 
	.A1(n6629), 
	.A0(\ram[10][11] ));
   OAI21XL U11224 (.Y(n13306), 
	.B0(n6828), 
	.A1(n13319), 
	.A0(n13318));
   NAND4X1 U11225 (.Y(n13319), 
	.D(n13323), 
	.C(n13322), 
	.B(n13321), 
	.A(n13320));
   AOI22X1 U11226 (.Y(n13323), 
	.B1(n6342), 
	.B0(\ram[249][11] ), 
	.A1(n6362), 
	.A0(\ram[248][11] ));
   AOI22X1 U11227 (.Y(n13322), 
	.B1(n6381), 
	.B0(\ram[247][11] ), 
	.A1(n6400), 
	.A0(\ram[246][11] ));
   AOI22X1 U11228 (.Y(n13321), 
	.B1(n6419), 
	.B0(\ram[245][11] ), 
	.A1(n6438), 
	.A0(\ram[244][11] ));
   AOI22X1 U11229 (.Y(n13320), 
	.B1(n6457), 
	.B0(\ram[243][11] ), 
	.A1(n6476), 
	.A0(\ram[242][11] ));
   NAND4X1 U11230 (.Y(n13318), 
	.D(n13327), 
	.C(n13326), 
	.B(n13325), 
	.A(n13324));
   AOI22X1 U11231 (.Y(n13327), 
	.B1(n6495), 
	.B0(\ram[241][11] ), 
	.A1(n6514), 
	.A0(\ram[240][11] ));
   AOI22X1 U11232 (.Y(n13326), 
	.B1(n6533), 
	.B0(\ram[255][11] ), 
	.A1(n6553), 
	.A0(\ram[254][11] ));
   AOI22X1 U11233 (.Y(n13325), 
	.B1(n6572), 
	.B0(\ram[253][11] ), 
	.A1(n6591), 
	.A0(\ram[252][11] ));
   AOI22X1 U11234 (.Y(n13324), 
	.B1(n6610), 
	.B0(\ram[251][11] ), 
	.A1(n6629), 
	.A0(\ram[250][11] ));
   OAI21XL U11235 (.Y(n13305), 
	.B0(n7117), 
	.A1(n13329), 
	.A0(n13328));
   NAND4X1 U11236 (.Y(n13329), 
	.D(n13333), 
	.C(n13332), 
	.B(n13331), 
	.A(n13330));
   AOI22X1 U11237 (.Y(n13333), 
	.B1(n6342), 
	.B0(\ram[233][11] ), 
	.A1(n6362), 
	.A0(\ram[232][11] ));
   AOI22X1 U11238 (.Y(n13332), 
	.B1(n6381), 
	.B0(\ram[231][11] ), 
	.A1(n6400), 
	.A0(\ram[230][11] ));
   AOI22X1 U11239 (.Y(n13331), 
	.B1(n6419), 
	.B0(\ram[229][11] ), 
	.A1(n6438), 
	.A0(\ram[228][11] ));
   AOI22X1 U11240 (.Y(n13330), 
	.B1(n6457), 
	.B0(\ram[227][11] ), 
	.A1(n6476), 
	.A0(\ram[226][11] ));
   NAND4X1 U11241 (.Y(n13328), 
	.D(n13337), 
	.C(n13336), 
	.B(n13335), 
	.A(n13334));
   AOI22X1 U11242 (.Y(n13337), 
	.B1(n6495), 
	.B0(\ram[225][11] ), 
	.A1(n6514), 
	.A0(\ram[224][11] ));
   AOI22X1 U11243 (.Y(n13336), 
	.B1(n6533), 
	.B0(\ram[239][11] ), 
	.A1(n6553), 
	.A0(\ram[238][11] ));
   AOI22X1 U11244 (.Y(n13335), 
	.B1(n6572), 
	.B0(\ram[237][11] ), 
	.A1(n6591), 
	.A0(\ram[236][11] ));
   AOI22X1 U11245 (.Y(n13334), 
	.B1(n6610), 
	.B0(\ram[235][11] ), 
	.A1(n6629), 
	.A0(\ram[234][11] ));
   OAI21XL U11246 (.Y(n13304), 
	.B0(n7406), 
	.A1(n13339), 
	.A0(n13338));
   NAND4X1 U11247 (.Y(n13339), 
	.D(n13343), 
	.C(n13342), 
	.B(n13341), 
	.A(n13340));
   AOI22X1 U11248 (.Y(n13343), 
	.B1(n6342), 
	.B0(\ram[217][11] ), 
	.A1(n6362), 
	.A0(\ram[216][11] ));
   AOI22X1 U11249 (.Y(n13342), 
	.B1(n6381), 
	.B0(\ram[215][11] ), 
	.A1(n6400), 
	.A0(\ram[214][11] ));
   AOI22X1 U11250 (.Y(n13341), 
	.B1(n6419), 
	.B0(\ram[213][11] ), 
	.A1(n6438), 
	.A0(\ram[212][11] ));
   AOI22X1 U11251 (.Y(n13340), 
	.B1(n6457), 
	.B0(\ram[211][11] ), 
	.A1(n6476), 
	.A0(\ram[210][11] ));
   NAND4X1 U11252 (.Y(n13338), 
	.D(n13347), 
	.C(n13346), 
	.B(n13345), 
	.A(n13344));
   AOI22X1 U11253 (.Y(n13347), 
	.B1(n6495), 
	.B0(\ram[209][11] ), 
	.A1(n6514), 
	.A0(\ram[208][11] ));
   AOI22X1 U11254 (.Y(n13346), 
	.B1(n6533), 
	.B0(\ram[223][11] ), 
	.A1(n6553), 
	.A0(\ram[222][11] ));
   AOI22X1 U11255 (.Y(n13345), 
	.B1(n6572), 
	.B0(\ram[221][11] ), 
	.A1(n6591), 
	.A0(\ram[220][11] ));
   AOI22X1 U11256 (.Y(n13344), 
	.B1(n6610), 
	.B0(\ram[219][11] ), 
	.A1(n6629), 
	.A0(\ram[218][11] ));
   NAND4X1 U11257 (.Y(n13302), 
	.D(n13351), 
	.C(n13350), 
	.B(n13349), 
	.A(n13348));
   OAI21XL U11258 (.Y(n13351), 
	.B0(n7695), 
	.A1(n13353), 
	.A0(n13352));
   NAND4X1 U11259 (.Y(n13353), 
	.D(n13357), 
	.C(n13356), 
	.B(n13355), 
	.A(n13354));
   AOI22X1 U11260 (.Y(n13357), 
	.B1(n6342), 
	.B0(\ram[201][11] ), 
	.A1(n6362), 
	.A0(\ram[200][11] ));
   AOI22X1 U11261 (.Y(n13356), 
	.B1(n6381), 
	.B0(\ram[199][11] ), 
	.A1(n6400), 
	.A0(\ram[198][11] ));
   AOI22X1 U11262 (.Y(n13355), 
	.B1(n6419), 
	.B0(\ram[197][11] ), 
	.A1(n6438), 
	.A0(\ram[196][11] ));
   AOI22X1 U11263 (.Y(n13354), 
	.B1(n6457), 
	.B0(\ram[195][11] ), 
	.A1(n6476), 
	.A0(\ram[194][11] ));
   NAND4X1 U11264 (.Y(n13352), 
	.D(n13361), 
	.C(n13360), 
	.B(n13359), 
	.A(n13358));
   AOI22X1 U11265 (.Y(n13361), 
	.B1(n6495), 
	.B0(\ram[193][11] ), 
	.A1(n6514), 
	.A0(\ram[192][11] ));
   AOI22X1 U11266 (.Y(n13360), 
	.B1(n6533), 
	.B0(\ram[207][11] ), 
	.A1(n6553), 
	.A0(\ram[206][11] ));
   AOI22X1 U11267 (.Y(n13359), 
	.B1(n6572), 
	.B0(\ram[205][11] ), 
	.A1(n6591), 
	.A0(\ram[204][11] ));
   AOI22X1 U11268 (.Y(n13358), 
	.B1(n6610), 
	.B0(\ram[203][11] ), 
	.A1(n6629), 
	.A0(\ram[202][11] ));
   OAI21XL U11269 (.Y(n13350), 
	.B0(n7984), 
	.A1(n13363), 
	.A0(n13362));
   NAND4X1 U11270 (.Y(n13363), 
	.D(n13367), 
	.C(n13366), 
	.B(n13365), 
	.A(n13364));
   AOI22X1 U11271 (.Y(n13367), 
	.B1(n6342), 
	.B0(\ram[185][11] ), 
	.A1(n6362), 
	.A0(\ram[184][11] ));
   AOI22X1 U11272 (.Y(n13366), 
	.B1(n6381), 
	.B0(\ram[183][11] ), 
	.A1(n6400), 
	.A0(\ram[182][11] ));
   AOI22X1 U11273 (.Y(n13365), 
	.B1(n6419), 
	.B0(\ram[181][11] ), 
	.A1(n6438), 
	.A0(\ram[180][11] ));
   AOI22X1 U11274 (.Y(n13364), 
	.B1(n6457), 
	.B0(\ram[179][11] ), 
	.A1(n6476), 
	.A0(\ram[178][11] ));
   NAND4X1 U11275 (.Y(n13362), 
	.D(n13371), 
	.C(n13370), 
	.B(n13369), 
	.A(n13368));
   AOI22X1 U11276 (.Y(n13371), 
	.B1(n6495), 
	.B0(\ram[177][11] ), 
	.A1(n6514), 
	.A0(\ram[176][11] ));
   AOI22X1 U11277 (.Y(n13370), 
	.B1(n6533), 
	.B0(\ram[191][11] ), 
	.A1(n6553), 
	.A0(\ram[190][11] ));
   AOI22X1 U11278 (.Y(n13369), 
	.B1(n6572), 
	.B0(\ram[189][11] ), 
	.A1(n6591), 
	.A0(\ram[188][11] ));
   AOI22X1 U11279 (.Y(n13368), 
	.B1(n6610), 
	.B0(\ram[187][11] ), 
	.A1(n6629), 
	.A0(\ram[186][11] ));
   OAI21XL U11280 (.Y(n13349), 
	.B0(n8273), 
	.A1(n13373), 
	.A0(n13372));
   NAND4X1 U11281 (.Y(n13373), 
	.D(n13377), 
	.C(n13376), 
	.B(n13375), 
	.A(n13374));
   AOI22X1 U11282 (.Y(n13377), 
	.B1(n6342), 
	.B0(\ram[169][11] ), 
	.A1(n6362), 
	.A0(\ram[168][11] ));
   AOI22X1 U11283 (.Y(n13376), 
	.B1(n6381), 
	.B0(\ram[167][11] ), 
	.A1(n6400), 
	.A0(\ram[166][11] ));
   AOI22X1 U11284 (.Y(n13375), 
	.B1(n6419), 
	.B0(\ram[165][11] ), 
	.A1(n6438), 
	.A0(\ram[164][11] ));
   AOI22X1 U11285 (.Y(n13374), 
	.B1(n6457), 
	.B0(\ram[163][11] ), 
	.A1(n6476), 
	.A0(\ram[162][11] ));
   NAND4X1 U11286 (.Y(n13372), 
	.D(n13381), 
	.C(n13380), 
	.B(n13379), 
	.A(n13378));
   AOI22X1 U11287 (.Y(n13381), 
	.B1(n6495), 
	.B0(\ram[161][11] ), 
	.A1(n6514), 
	.A0(\ram[160][11] ));
   AOI22X1 U11288 (.Y(n13380), 
	.B1(n6533), 
	.B0(\ram[175][11] ), 
	.A1(n6553), 
	.A0(\ram[174][11] ));
   AOI22X1 U11289 (.Y(n13379), 
	.B1(n6572), 
	.B0(\ram[173][11] ), 
	.A1(n6591), 
	.A0(\ram[172][11] ));
   AOI22X1 U11290 (.Y(n13378), 
	.B1(n6610), 
	.B0(\ram[171][11] ), 
	.A1(n6629), 
	.A0(\ram[170][11] ));
   OAI21XL U11291 (.Y(n13348), 
	.B0(n8562), 
	.A1(n13383), 
	.A0(n13382));
   NAND4X1 U11292 (.Y(n13383), 
	.D(n13387), 
	.C(n13386), 
	.B(n13385), 
	.A(n13384));
   AOI22X1 U11293 (.Y(n13387), 
	.B1(n6342), 
	.B0(\ram[153][11] ), 
	.A1(n6362), 
	.A0(\ram[152][11] ));
   AOI22X1 U11294 (.Y(n13386), 
	.B1(n6381), 
	.B0(\ram[151][11] ), 
	.A1(n6400), 
	.A0(\ram[150][11] ));
   AOI22X1 U11295 (.Y(n13385), 
	.B1(n6419), 
	.B0(\ram[149][11] ), 
	.A1(n6438), 
	.A0(\ram[148][11] ));
   AOI22X1 U11296 (.Y(n13384), 
	.B1(n6457), 
	.B0(\ram[147][11] ), 
	.A1(n6476), 
	.A0(\ram[146][11] ));
   NAND4X1 U11297 (.Y(n13382), 
	.D(n13391), 
	.C(n13390), 
	.B(n13389), 
	.A(n13388));
   AOI22X1 U11298 (.Y(n13391), 
	.B1(n6495), 
	.B0(\ram[145][11] ), 
	.A1(n6514), 
	.A0(\ram[144][11] ));
   AOI22X1 U11299 (.Y(n13390), 
	.B1(n6533), 
	.B0(\ram[159][11] ), 
	.A1(n6553), 
	.A0(\ram[158][11] ));
   AOI22X1 U11300 (.Y(n13389), 
	.B1(n6572), 
	.B0(\ram[157][11] ), 
	.A1(n6591), 
	.A0(\ram[156][11] ));
   AOI22X1 U11301 (.Y(n13388), 
	.B1(n6610), 
	.B0(\ram[155][11] ), 
	.A1(n6629), 
	.A0(\ram[154][11] ));
   NAND4X1 U11302 (.Y(n13301), 
	.D(n13395), 
	.C(n13394), 
	.B(n13393), 
	.A(n13392));
   OAI21XL U11303 (.Y(n13395), 
	.B0(n8851), 
	.A1(n13397), 
	.A0(n13396));
   NAND4X1 U11304 (.Y(n13397), 
	.D(n13401), 
	.C(n13400), 
	.B(n13399), 
	.A(n13398));
   AOI22X1 U11305 (.Y(n13401), 
	.B1(n6342), 
	.B0(\ram[137][11] ), 
	.A1(n6362), 
	.A0(\ram[136][11] ));
   AOI22X1 U11306 (.Y(n13400), 
	.B1(n6381), 
	.B0(\ram[135][11] ), 
	.A1(n6400), 
	.A0(\ram[134][11] ));
   AOI22X1 U11307 (.Y(n13399), 
	.B1(n6419), 
	.B0(\ram[133][11] ), 
	.A1(n6438), 
	.A0(\ram[132][11] ));
   AOI22X1 U11308 (.Y(n13398), 
	.B1(n6457), 
	.B0(\ram[131][11] ), 
	.A1(n6476), 
	.A0(\ram[130][11] ));
   NAND4X1 U11309 (.Y(n13396), 
	.D(n13405), 
	.C(n13404), 
	.B(n13403), 
	.A(n13402));
   AOI22X1 U11310 (.Y(n13405), 
	.B1(n6495), 
	.B0(\ram[129][11] ), 
	.A1(n6514), 
	.A0(\ram[128][11] ));
   AOI22X1 U11311 (.Y(n13404), 
	.B1(n6533), 
	.B0(\ram[143][11] ), 
	.A1(n6553), 
	.A0(\ram[142][11] ));
   AOI22X1 U11312 (.Y(n13403), 
	.B1(n6572), 
	.B0(\ram[141][11] ), 
	.A1(n6591), 
	.A0(\ram[140][11] ));
   AOI22X1 U11313 (.Y(n13402), 
	.B1(n6610), 
	.B0(\ram[139][11] ), 
	.A1(n6629), 
	.A0(\ram[138][11] ));
   OAI21XL U11314 (.Y(n13394), 
	.B0(n9140), 
	.A1(n13407), 
	.A0(n13406));
   NAND4X1 U11315 (.Y(n13407), 
	.D(n13411), 
	.C(n13410), 
	.B(n13409), 
	.A(n13408));
   AOI22X1 U11316 (.Y(n13411), 
	.B1(n6342), 
	.B0(\ram[121][11] ), 
	.A1(n6362), 
	.A0(\ram[120][11] ));
   AOI22X1 U11317 (.Y(n13410), 
	.B1(n6381), 
	.B0(\ram[119][11] ), 
	.A1(n6400), 
	.A0(\ram[118][11] ));
   AOI22X1 U11318 (.Y(n13409), 
	.B1(n6419), 
	.B0(\ram[117][11] ), 
	.A1(n6438), 
	.A0(\ram[116][11] ));
   AOI22X1 U11319 (.Y(n13408), 
	.B1(n6457), 
	.B0(\ram[115][11] ), 
	.A1(n6476), 
	.A0(\ram[114][11] ));
   NAND4X1 U11320 (.Y(n13406), 
	.D(n13415), 
	.C(n13414), 
	.B(n13413), 
	.A(n13412));
   AOI22X1 U11321 (.Y(n13415), 
	.B1(n6495), 
	.B0(\ram[113][11] ), 
	.A1(n6514), 
	.A0(\ram[112][11] ));
   AOI22X1 U11322 (.Y(n13414), 
	.B1(n6533), 
	.B0(\ram[127][11] ), 
	.A1(n6553), 
	.A0(\ram[126][11] ));
   AOI22X1 U11323 (.Y(n13413), 
	.B1(n6572), 
	.B0(\ram[125][11] ), 
	.A1(n6591), 
	.A0(\ram[124][11] ));
   AOI22X1 U11324 (.Y(n13412), 
	.B1(n6610), 
	.B0(\ram[123][11] ), 
	.A1(n6629), 
	.A0(\ram[122][11] ));
   OAI21XL U11325 (.Y(n13393), 
	.B0(n9429), 
	.A1(n13417), 
	.A0(n13416));
   NAND4X1 U11326 (.Y(n13417), 
	.D(n13421), 
	.C(n13420), 
	.B(n13419), 
	.A(n13418));
   AOI22X1 U11327 (.Y(n13421), 
	.B1(n6342), 
	.B0(\ram[105][11] ), 
	.A1(n6362), 
	.A0(\ram[104][11] ));
   AOI22X1 U11328 (.Y(n13420), 
	.B1(n6381), 
	.B0(\ram[103][11] ), 
	.A1(n6400), 
	.A0(\ram[102][11] ));
   AOI22X1 U11329 (.Y(n13419), 
	.B1(n6419), 
	.B0(\ram[101][11] ), 
	.A1(n6438), 
	.A0(\ram[100][11] ));
   AOI22X1 U11330 (.Y(n13418), 
	.B1(n6457), 
	.B0(\ram[99][11] ), 
	.A1(n6476), 
	.A0(\ram[98][11] ));
   NAND4X1 U11331 (.Y(n13416), 
	.D(n13425), 
	.C(n13424), 
	.B(n13423), 
	.A(n13422));
   AOI22X1 U11332 (.Y(n13425), 
	.B1(n6495), 
	.B0(\ram[97][11] ), 
	.A1(n6514), 
	.A0(\ram[96][11] ));
   AOI22X1 U11333 (.Y(n13424), 
	.B1(n6533), 
	.B0(\ram[111][11] ), 
	.A1(n6553), 
	.A0(\ram[110][11] ));
   AOI22X1 U11334 (.Y(n13423), 
	.B1(n6572), 
	.B0(\ram[109][11] ), 
	.A1(n6591), 
	.A0(\ram[108][11] ));
   AOI22X1 U11335 (.Y(n13422), 
	.B1(n6610), 
	.B0(\ram[107][11] ), 
	.A1(n6629), 
	.A0(\ram[106][11] ));
   OAI21XL U11336 (.Y(n13392), 
	.B0(n9718), 
	.A1(n13427), 
	.A0(n13426));
   NAND4X1 U11337 (.Y(n13427), 
	.D(n13431), 
	.C(n13430), 
	.B(n13429), 
	.A(n13428));
   AOI22X1 U11338 (.Y(n13431), 
	.B1(n6342), 
	.B0(\ram[89][11] ), 
	.A1(n6362), 
	.A0(\ram[88][11] ));
   AOI22X1 U11339 (.Y(n13430), 
	.B1(n6381), 
	.B0(\ram[87][11] ), 
	.A1(n6400), 
	.A0(\ram[86][11] ));
   AOI22X1 U11340 (.Y(n13429), 
	.B1(n6419), 
	.B0(\ram[85][11] ), 
	.A1(n6438), 
	.A0(\ram[84][11] ));
   AOI22X1 U11341 (.Y(n13428), 
	.B1(n6457), 
	.B0(\ram[83][11] ), 
	.A1(n6476), 
	.A0(\ram[82][11] ));
   NAND4X1 U11342 (.Y(n13426), 
	.D(n13435), 
	.C(n13434), 
	.B(n13433), 
	.A(n13432));
   AOI22X1 U11343 (.Y(n13435), 
	.B1(n6495), 
	.B0(\ram[81][11] ), 
	.A1(n6514), 
	.A0(\ram[80][11] ));
   AOI22X1 U11344 (.Y(n13434), 
	.B1(n6533), 
	.B0(\ram[95][11] ), 
	.A1(n6553), 
	.A0(\ram[94][11] ));
   AOI22X1 U11345 (.Y(n13433), 
	.B1(n6572), 
	.B0(\ram[93][11] ), 
	.A1(n6591), 
	.A0(\ram[92][11] ));
   AOI22X1 U11346 (.Y(n13432), 
	.B1(n6610), 
	.B0(\ram[91][11] ), 
	.A1(n6629), 
	.A0(\ram[90][11] ));
   NAND4X1 U11347 (.Y(n13300), 
	.D(n13439), 
	.C(n13438), 
	.B(n13437), 
	.A(n13436));
   OAI21XL U11348 (.Y(n13439), 
	.B0(n10007), 
	.A1(n13441), 
	.A0(n13440));
   NAND4X1 U11349 (.Y(n13441), 
	.D(n13445), 
	.C(n13444), 
	.B(n13443), 
	.A(n13442));
   AOI22X1 U11350 (.Y(n13445), 
	.B1(n6342), 
	.B0(\ram[73][11] ), 
	.A1(n6362), 
	.A0(\ram[72][11] ));
   AOI22X1 U11351 (.Y(n13444), 
	.B1(n6381), 
	.B0(\ram[71][11] ), 
	.A1(n6400), 
	.A0(\ram[70][11] ));
   AOI22X1 U11352 (.Y(n13443), 
	.B1(n6419), 
	.B0(\ram[69][11] ), 
	.A1(n6438), 
	.A0(\ram[68][11] ));
   AOI22X1 U11353 (.Y(n13442), 
	.B1(n6457), 
	.B0(\ram[67][11] ), 
	.A1(n6476), 
	.A0(\ram[66][11] ));
   NAND4X1 U11354 (.Y(n13440), 
	.D(n13449), 
	.C(n13448), 
	.B(n13447), 
	.A(n13446));
   AOI22X1 U11355 (.Y(n13449), 
	.B1(n6495), 
	.B0(\ram[65][11] ), 
	.A1(n6514), 
	.A0(\ram[64][11] ));
   AOI22X1 U11356 (.Y(n13448), 
	.B1(n6533), 
	.B0(\ram[79][11] ), 
	.A1(n6553), 
	.A0(\ram[78][11] ));
   AOI22X1 U11357 (.Y(n13447), 
	.B1(n6572), 
	.B0(\ram[77][11] ), 
	.A1(n6591), 
	.A0(\ram[76][11] ));
   AOI22X1 U11358 (.Y(n13446), 
	.B1(n6610), 
	.B0(\ram[75][11] ), 
	.A1(n6629), 
	.A0(\ram[74][11] ));
   OAI21XL U11359 (.Y(n13438), 
	.B0(n10296), 
	.A1(n13451), 
	.A0(n13450));
   NAND4X1 U11360 (.Y(n13451), 
	.D(n13455), 
	.C(n13454), 
	.B(n13453), 
	.A(n13452));
   AOI22X1 U11361 (.Y(n13455), 
	.B1(n6342), 
	.B0(\ram[57][11] ), 
	.A1(n6362), 
	.A0(\ram[56][11] ));
   AOI22X1 U11362 (.Y(n13454), 
	.B1(n6381), 
	.B0(\ram[55][11] ), 
	.A1(n6400), 
	.A0(\ram[54][11] ));
   AOI22X1 U11363 (.Y(n13453), 
	.B1(n6419), 
	.B0(\ram[53][11] ), 
	.A1(n6438), 
	.A0(\ram[52][11] ));
   AOI22X1 U11364 (.Y(n13452), 
	.B1(n6457), 
	.B0(\ram[51][11] ), 
	.A1(n6476), 
	.A0(\ram[50][11] ));
   NAND4X1 U11365 (.Y(n13450), 
	.D(n13459), 
	.C(n13458), 
	.B(n13457), 
	.A(n13456));
   AOI22X1 U11366 (.Y(n13459), 
	.B1(n6495), 
	.B0(\ram[49][11] ), 
	.A1(n6514), 
	.A0(\ram[48][11] ));
   AOI22X1 U11367 (.Y(n13458), 
	.B1(n6533), 
	.B0(\ram[63][11] ), 
	.A1(n6553), 
	.A0(\ram[62][11] ));
   AOI22X1 U11368 (.Y(n13457), 
	.B1(n6572), 
	.B0(\ram[61][11] ), 
	.A1(n6591), 
	.A0(\ram[60][11] ));
   AOI22X1 U11369 (.Y(n13456), 
	.B1(n6610), 
	.B0(\ram[59][11] ), 
	.A1(n6629), 
	.A0(\ram[58][11] ));
   OAI21XL U11370 (.Y(n13437), 
	.B0(n10585), 
	.A1(n13461), 
	.A0(n13460));
   NAND4X1 U11371 (.Y(n13461), 
	.D(n13465), 
	.C(n13464), 
	.B(n13463), 
	.A(n13462));
   AOI22X1 U11372 (.Y(n13465), 
	.B1(n6342), 
	.B0(\ram[41][11] ), 
	.A1(n6362), 
	.A0(\ram[40][11] ));
   AOI22X1 U11373 (.Y(n13464), 
	.B1(n6381), 
	.B0(\ram[39][11] ), 
	.A1(n6400), 
	.A0(\ram[38][11] ));
   AOI22X1 U11374 (.Y(n13463), 
	.B1(n6419), 
	.B0(\ram[37][11] ), 
	.A1(n6438), 
	.A0(\ram[36][11] ));
   AOI22X1 U11375 (.Y(n13462), 
	.B1(n6457), 
	.B0(\ram[35][11] ), 
	.A1(n6476), 
	.A0(\ram[34][11] ));
   NAND4X1 U11376 (.Y(n13460), 
	.D(n13469), 
	.C(n13468), 
	.B(n13467), 
	.A(n13466));
   AOI22X1 U11377 (.Y(n13469), 
	.B1(n6495), 
	.B0(\ram[33][11] ), 
	.A1(n6514), 
	.A0(\ram[32][11] ));
   AOI22X1 U11378 (.Y(n13468), 
	.B1(n6533), 
	.B0(\ram[47][11] ), 
	.A1(n6553), 
	.A0(\ram[46][11] ));
   AOI22X1 U11379 (.Y(n13467), 
	.B1(n6572), 
	.B0(\ram[45][11] ), 
	.A1(n6591), 
	.A0(\ram[44][11] ));
   AOI22X1 U11380 (.Y(n13466), 
	.B1(n6610), 
	.B0(\ram[43][11] ), 
	.A1(n6629), 
	.A0(\ram[42][11] ));
   OAI21XL U11381 (.Y(n13436), 
	.B0(n6343), 
	.A1(n13471), 
	.A0(n13470));
   NAND4X1 U11382 (.Y(n13471), 
	.D(n13475), 
	.C(n13474), 
	.B(n13473), 
	.A(n13472));
   AOI22X1 U11383 (.Y(n13475), 
	.B1(n6342), 
	.B0(\ram[25][11] ), 
	.A1(n6362), 
	.A0(\ram[24][11] ));
   AOI22X1 U11384 (.Y(n13474), 
	.B1(n6381), 
	.B0(\ram[23][11] ), 
	.A1(n6400), 
	.A0(\ram[22][11] ));
   AOI22X1 U11385 (.Y(n13473), 
	.B1(n6419), 
	.B0(\ram[21][11] ), 
	.A1(n6438), 
	.A0(\ram[20][11] ));
   AOI22X1 U11386 (.Y(n13472), 
	.B1(n6457), 
	.B0(\ram[19][11] ), 
	.A1(n6476), 
	.A0(\ram[18][11] ));
   NAND4X1 U11387 (.Y(n13470), 
	.D(n13479), 
	.C(n13478), 
	.B(n13477), 
	.A(n13476));
   AOI22X1 U11388 (.Y(n13479), 
	.B1(n6495), 
	.B0(\ram[17][11] ), 
	.A1(n6514), 
	.A0(\ram[16][11] ));
   AOI22X1 U11389 (.Y(n13478), 
	.B1(n6533), 
	.B0(\ram[31][11] ), 
	.A1(n6553), 
	.A0(\ram[30][11] ));
   AOI22X1 U11390 (.Y(n13477), 
	.B1(n6572), 
	.B0(\ram[29][11] ), 
	.A1(n6591), 
	.A0(\ram[28][11] ));
   AOI22X1 U11391 (.Y(n13476), 
	.B1(n6610), 
	.B0(\ram[27][11] ), 
	.A1(n6629), 
	.A0(\ram[26][11] ));
   OR4X1 U11392 (.Y(mem_read_data[10]), 
	.D(n13483), 
	.C(n13482), 
	.B(n13481), 
	.A(n13480));
   NAND4X1 U11393 (.Y(n13483), 
	.D(n13487), 
	.C(n13486), 
	.B(n13485), 
	.A(n13484));
   OAI21XL U11394 (.Y(n13487), 
	.B0(n6534), 
	.A1(n13489), 
	.A0(n13488));
   NAND4X1 U11395 (.Y(n13489), 
	.D(n13493), 
	.C(n13492), 
	.B(n13491), 
	.A(n13490));
   AOI22X1 U11396 (.Y(n13493), 
	.B1(n6342), 
	.B0(\ram[9][10] ), 
	.A1(n6362), 
	.A0(\ram[8][10] ));
   AOI22X1 U11397 (.Y(n13492), 
	.B1(n6381), 
	.B0(\ram[7][10] ), 
	.A1(n6400), 
	.A0(\ram[6][10] ));
   AOI22X1 U11398 (.Y(n13491), 
	.B1(n6419), 
	.B0(\ram[5][10] ), 
	.A1(n6438), 
	.A0(\ram[4][10] ));
   AOI22X1 U11399 (.Y(n13490), 
	.B1(n6457), 
	.B0(\ram[3][10] ), 
	.A1(n6476), 
	.A0(\ram[2][10] ));
   NAND4X1 U11400 (.Y(n13488), 
	.D(n13497), 
	.C(n13496), 
	.B(n13495), 
	.A(n13494));
   AOI22X1 U11401 (.Y(n13497), 
	.B1(n6495), 
	.B0(\ram[1][10] ), 
	.A1(n6514), 
	.A0(\ram[0][10] ));
   AOI22X1 U11402 (.Y(n13496), 
	.B1(n6533), 
	.B0(\ram[15][10] ), 
	.A1(n6553), 
	.A0(\ram[14][10] ));
   AOI22X1 U11403 (.Y(n13495), 
	.B1(n6572), 
	.B0(\ram[13][10] ), 
	.A1(n6591), 
	.A0(\ram[12][10] ));
   AOI22X1 U11404 (.Y(n13494), 
	.B1(n6610), 
	.B0(\ram[11][10] ), 
	.A1(n6629), 
	.A0(\ram[10][10] ));
   OAI21XL U11405 (.Y(n13486), 
	.B0(n6828), 
	.A1(n13499), 
	.A0(n13498));
   NAND4X1 U11406 (.Y(n13499), 
	.D(n13503), 
	.C(n13502), 
	.B(n13501), 
	.A(n13500));
   AOI22X1 U11407 (.Y(n13503), 
	.B1(n6342), 
	.B0(\ram[249][10] ), 
	.A1(n6362), 
	.A0(\ram[248][10] ));
   AOI22X1 U11408 (.Y(n13502), 
	.B1(n6381), 
	.B0(\ram[247][10] ), 
	.A1(n6400), 
	.A0(\ram[246][10] ));
   AOI22X1 U11409 (.Y(n13501), 
	.B1(n6419), 
	.B0(\ram[245][10] ), 
	.A1(n6438), 
	.A0(\ram[244][10] ));
   AOI22X1 U11410 (.Y(n13500), 
	.B1(n6457), 
	.B0(\ram[243][10] ), 
	.A1(n6476), 
	.A0(\ram[242][10] ));
   NAND4X1 U11411 (.Y(n13498), 
	.D(n13507), 
	.C(n13506), 
	.B(n13505), 
	.A(n13504));
   AOI22X1 U11412 (.Y(n13507), 
	.B1(n6495), 
	.B0(\ram[241][10] ), 
	.A1(n6514), 
	.A0(\ram[240][10] ));
   AOI22X1 U11413 (.Y(n13506), 
	.B1(n6533), 
	.B0(\ram[255][10] ), 
	.A1(n6553), 
	.A0(\ram[254][10] ));
   AOI22X1 U11414 (.Y(n13505), 
	.B1(n6572), 
	.B0(\ram[253][10] ), 
	.A1(n6591), 
	.A0(\ram[252][10] ));
   AOI22X1 U11415 (.Y(n13504), 
	.B1(n6610), 
	.B0(\ram[251][10] ), 
	.A1(n6629), 
	.A0(\ram[250][10] ));
   OAI21XL U11416 (.Y(n13485), 
	.B0(n7117), 
	.A1(n13509), 
	.A0(n13508));
   NAND4X1 U11417 (.Y(n13509), 
	.D(n13513), 
	.C(n13512), 
	.B(n13511), 
	.A(n13510));
   AOI22X1 U11418 (.Y(n13513), 
	.B1(n6342), 
	.B0(\ram[233][10] ), 
	.A1(n6362), 
	.A0(\ram[232][10] ));
   AOI22X1 U11419 (.Y(n13512), 
	.B1(n6381), 
	.B0(\ram[231][10] ), 
	.A1(n6400), 
	.A0(\ram[230][10] ));
   AOI22X1 U11420 (.Y(n13511), 
	.B1(n6419), 
	.B0(\ram[229][10] ), 
	.A1(n6438), 
	.A0(\ram[228][10] ));
   AOI22X1 U11421 (.Y(n13510), 
	.B1(n6457), 
	.B0(\ram[227][10] ), 
	.A1(n6476), 
	.A0(\ram[226][10] ));
   NAND4X1 U11422 (.Y(n13508), 
	.D(n13517), 
	.C(n13516), 
	.B(n13515), 
	.A(n13514));
   AOI22X1 U11423 (.Y(n13517), 
	.B1(n6495), 
	.B0(\ram[225][10] ), 
	.A1(n6514), 
	.A0(\ram[224][10] ));
   AOI22X1 U11424 (.Y(n13516), 
	.B1(n6533), 
	.B0(\ram[239][10] ), 
	.A1(n6553), 
	.A0(\ram[238][10] ));
   AOI22X1 U11425 (.Y(n13515), 
	.B1(n6572), 
	.B0(\ram[237][10] ), 
	.A1(n6591), 
	.A0(\ram[236][10] ));
   AOI22X1 U11426 (.Y(n13514), 
	.B1(n6610), 
	.B0(\ram[235][10] ), 
	.A1(n6629), 
	.A0(\ram[234][10] ));
   OAI21XL U11427 (.Y(n13484), 
	.B0(n7406), 
	.A1(n13519), 
	.A0(n13518));
   NAND4X1 U11428 (.Y(n13519), 
	.D(n13523), 
	.C(n13522), 
	.B(n13521), 
	.A(n13520));
   AOI22X1 U11429 (.Y(n13523), 
	.B1(n6342), 
	.B0(\ram[217][10] ), 
	.A1(n6362), 
	.A0(\ram[216][10] ));
   AOI22X1 U11430 (.Y(n13522), 
	.B1(n6381), 
	.B0(\ram[215][10] ), 
	.A1(n6400), 
	.A0(\ram[214][10] ));
   AOI22X1 U11431 (.Y(n13521), 
	.B1(n6419), 
	.B0(\ram[213][10] ), 
	.A1(n6438), 
	.A0(\ram[212][10] ));
   AOI22X1 U11432 (.Y(n13520), 
	.B1(n6457), 
	.B0(\ram[211][10] ), 
	.A1(n6476), 
	.A0(\ram[210][10] ));
   NAND4X1 U11433 (.Y(n13518), 
	.D(n13527), 
	.C(n13526), 
	.B(n13525), 
	.A(n13524));
   AOI22X1 U11434 (.Y(n13527), 
	.B1(n6495), 
	.B0(\ram[209][10] ), 
	.A1(n6514), 
	.A0(\ram[208][10] ));
   AOI22X1 U11435 (.Y(n13526), 
	.B1(n6533), 
	.B0(\ram[223][10] ), 
	.A1(n6553), 
	.A0(\ram[222][10] ));
   AOI22X1 U11436 (.Y(n13525), 
	.B1(n6572), 
	.B0(\ram[221][10] ), 
	.A1(n6591), 
	.A0(\ram[220][10] ));
   AOI22X1 U11437 (.Y(n13524), 
	.B1(n6610), 
	.B0(\ram[219][10] ), 
	.A1(n6629), 
	.A0(\ram[218][10] ));
   NAND4X1 U11438 (.Y(n13482), 
	.D(n13531), 
	.C(n13530), 
	.B(n13529), 
	.A(n13528));
   OAI21XL U11439 (.Y(n13531), 
	.B0(n7695), 
	.A1(n13533), 
	.A0(n13532));
   NAND4X1 U11440 (.Y(n13533), 
	.D(n13537), 
	.C(n13536), 
	.B(n13535), 
	.A(n13534));
   AOI22X1 U11441 (.Y(n13537), 
	.B1(n6342), 
	.B0(\ram[201][10] ), 
	.A1(n6362), 
	.A0(\ram[200][10] ));
   AOI22X1 U11442 (.Y(n13536), 
	.B1(n6381), 
	.B0(\ram[199][10] ), 
	.A1(n6400), 
	.A0(\ram[198][10] ));
   AOI22X1 U11443 (.Y(n13535), 
	.B1(n6419), 
	.B0(\ram[197][10] ), 
	.A1(n6438), 
	.A0(\ram[196][10] ));
   AOI22X1 U11444 (.Y(n13534), 
	.B1(n6457), 
	.B0(\ram[195][10] ), 
	.A1(n6476), 
	.A0(\ram[194][10] ));
   NAND4X1 U11445 (.Y(n13532), 
	.D(n13541), 
	.C(n13540), 
	.B(n13539), 
	.A(n13538));
   AOI22X1 U11446 (.Y(n13541), 
	.B1(n6495), 
	.B0(\ram[193][10] ), 
	.A1(n6514), 
	.A0(\ram[192][10] ));
   AOI22X1 U11447 (.Y(n13540), 
	.B1(n6533), 
	.B0(\ram[207][10] ), 
	.A1(n6553), 
	.A0(\ram[206][10] ));
   AOI22X1 U11448 (.Y(n13539), 
	.B1(n6572), 
	.B0(\ram[205][10] ), 
	.A1(n6591), 
	.A0(\ram[204][10] ));
   AOI22X1 U11449 (.Y(n13538), 
	.B1(n6610), 
	.B0(\ram[203][10] ), 
	.A1(n6629), 
	.A0(\ram[202][10] ));
   OAI21XL U11450 (.Y(n13530), 
	.B0(n7984), 
	.A1(n13543), 
	.A0(n13542));
   NAND4X1 U11451 (.Y(n13543), 
	.D(n13547), 
	.C(n13546), 
	.B(n13545), 
	.A(n13544));
   AOI22X1 U11452 (.Y(n13547), 
	.B1(n6342), 
	.B0(\ram[185][10] ), 
	.A1(n6362), 
	.A0(\ram[184][10] ));
   AOI22X1 U11453 (.Y(n13546), 
	.B1(n6381), 
	.B0(\ram[183][10] ), 
	.A1(n6400), 
	.A0(\ram[182][10] ));
   AOI22X1 U11454 (.Y(n13545), 
	.B1(n6419), 
	.B0(\ram[181][10] ), 
	.A1(n6438), 
	.A0(\ram[180][10] ));
   AOI22X1 U11455 (.Y(n13544), 
	.B1(n6457), 
	.B0(\ram[179][10] ), 
	.A1(n6476), 
	.A0(\ram[178][10] ));
   NAND4X1 U11456 (.Y(n13542), 
	.D(n13551), 
	.C(n13550), 
	.B(n13549), 
	.A(n13548));
   AOI22X1 U11457 (.Y(n13551), 
	.B1(n6495), 
	.B0(\ram[177][10] ), 
	.A1(n6514), 
	.A0(\ram[176][10] ));
   AOI22X1 U11458 (.Y(n13550), 
	.B1(n6533), 
	.B0(\ram[191][10] ), 
	.A1(n6553), 
	.A0(\ram[190][10] ));
   AOI22X1 U11459 (.Y(n13549), 
	.B1(n6572), 
	.B0(\ram[189][10] ), 
	.A1(n6591), 
	.A0(\ram[188][10] ));
   AOI22X1 U11460 (.Y(n13548), 
	.B1(n6610), 
	.B0(\ram[187][10] ), 
	.A1(n6629), 
	.A0(\ram[186][10] ));
   OAI21XL U11461 (.Y(n13529), 
	.B0(n8273), 
	.A1(n13553), 
	.A0(n13552));
   NAND4X1 U11462 (.Y(n13553), 
	.D(n13557), 
	.C(n13556), 
	.B(n13555), 
	.A(n13554));
   AOI22X1 U11463 (.Y(n13557), 
	.B1(n6342), 
	.B0(\ram[169][10] ), 
	.A1(n6362), 
	.A0(\ram[168][10] ));
   AOI22X1 U11464 (.Y(n13556), 
	.B1(n6381), 
	.B0(\ram[167][10] ), 
	.A1(n6400), 
	.A0(\ram[166][10] ));
   AOI22X1 U11465 (.Y(n13555), 
	.B1(n6419), 
	.B0(\ram[165][10] ), 
	.A1(n6438), 
	.A0(\ram[164][10] ));
   AOI22X1 U11466 (.Y(n13554), 
	.B1(n6457), 
	.B0(\ram[163][10] ), 
	.A1(n6476), 
	.A0(\ram[162][10] ));
   NAND4X1 U11467 (.Y(n13552), 
	.D(n13561), 
	.C(n13560), 
	.B(n13559), 
	.A(n13558));
   AOI22X1 U11468 (.Y(n13561), 
	.B1(n6495), 
	.B0(\ram[161][10] ), 
	.A1(n6514), 
	.A0(\ram[160][10] ));
   AOI22X1 U11469 (.Y(n13560), 
	.B1(n6533), 
	.B0(\ram[175][10] ), 
	.A1(n6553), 
	.A0(\ram[174][10] ));
   AOI22X1 U11470 (.Y(n13559), 
	.B1(n6572), 
	.B0(\ram[173][10] ), 
	.A1(n6591), 
	.A0(\ram[172][10] ));
   AOI22X1 U11471 (.Y(n13558), 
	.B1(n6610), 
	.B0(\ram[171][10] ), 
	.A1(n6629), 
	.A0(\ram[170][10] ));
   OAI21XL U11472 (.Y(n13528), 
	.B0(n8562), 
	.A1(n13563), 
	.A0(n13562));
   NAND4X1 U11473 (.Y(n13563), 
	.D(n13567), 
	.C(n13566), 
	.B(n13565), 
	.A(n13564));
   AOI22X1 U11474 (.Y(n13567), 
	.B1(n6342), 
	.B0(\ram[153][10] ), 
	.A1(n6362), 
	.A0(\ram[152][10] ));
   AOI22X1 U11475 (.Y(n13566), 
	.B1(n6381), 
	.B0(\ram[151][10] ), 
	.A1(n6400), 
	.A0(\ram[150][10] ));
   AOI22X1 U11476 (.Y(n13565), 
	.B1(n6419), 
	.B0(\ram[149][10] ), 
	.A1(n6438), 
	.A0(\ram[148][10] ));
   AOI22X1 U11477 (.Y(n13564), 
	.B1(n6457), 
	.B0(\ram[147][10] ), 
	.A1(n6476), 
	.A0(\ram[146][10] ));
   NAND4X1 U11478 (.Y(n13562), 
	.D(n13571), 
	.C(n13570), 
	.B(n13569), 
	.A(n13568));
   AOI22X1 U11479 (.Y(n13571), 
	.B1(n6495), 
	.B0(\ram[145][10] ), 
	.A1(n6514), 
	.A0(\ram[144][10] ));
   AOI22X1 U11480 (.Y(n13570), 
	.B1(n6533), 
	.B0(\ram[159][10] ), 
	.A1(n6553), 
	.A0(\ram[158][10] ));
   AOI22X1 U11481 (.Y(n13569), 
	.B1(n6572), 
	.B0(\ram[157][10] ), 
	.A1(n6591), 
	.A0(\ram[156][10] ));
   AOI22X1 U11482 (.Y(n13568), 
	.B1(n6610), 
	.B0(\ram[155][10] ), 
	.A1(n6629), 
	.A0(\ram[154][10] ));
   NAND4X1 U11483 (.Y(n13481), 
	.D(n13575), 
	.C(n13574), 
	.B(n13573), 
	.A(n13572));
   OAI21XL U11484 (.Y(n13575), 
	.B0(n8851), 
	.A1(n13577), 
	.A0(n13576));
   NAND4X1 U11485 (.Y(n13577), 
	.D(n13581), 
	.C(n13580), 
	.B(n13579), 
	.A(n13578));
   AOI22X1 U11486 (.Y(n13581), 
	.B1(n6342), 
	.B0(\ram[137][10] ), 
	.A1(n6362), 
	.A0(\ram[136][10] ));
   AOI22X1 U11487 (.Y(n13580), 
	.B1(n6381), 
	.B0(\ram[135][10] ), 
	.A1(n6400), 
	.A0(\ram[134][10] ));
   AOI22X1 U11488 (.Y(n13579), 
	.B1(n6419), 
	.B0(\ram[133][10] ), 
	.A1(n6438), 
	.A0(\ram[132][10] ));
   AOI22X1 U11489 (.Y(n13578), 
	.B1(n6457), 
	.B0(\ram[131][10] ), 
	.A1(n6476), 
	.A0(\ram[130][10] ));
   NAND4X1 U11490 (.Y(n13576), 
	.D(n13585), 
	.C(n13584), 
	.B(n13583), 
	.A(n13582));
   AOI22X1 U11491 (.Y(n13585), 
	.B1(n6495), 
	.B0(\ram[129][10] ), 
	.A1(n6514), 
	.A0(\ram[128][10] ));
   AOI22X1 U11492 (.Y(n13584), 
	.B1(n6533), 
	.B0(\ram[143][10] ), 
	.A1(n6553), 
	.A0(\ram[142][10] ));
   AOI22X1 U11493 (.Y(n13583), 
	.B1(n6572), 
	.B0(\ram[141][10] ), 
	.A1(n6591), 
	.A0(\ram[140][10] ));
   AOI22X1 U11494 (.Y(n13582), 
	.B1(n6610), 
	.B0(\ram[139][10] ), 
	.A1(n6629), 
	.A0(\ram[138][10] ));
   OAI21XL U11495 (.Y(n13574), 
	.B0(n9140), 
	.A1(n13587), 
	.A0(n13586));
   NAND4X1 U11496 (.Y(n13587), 
	.D(n13591), 
	.C(n13590), 
	.B(n13589), 
	.A(n13588));
   AOI22X1 U11497 (.Y(n13591), 
	.B1(n6342), 
	.B0(\ram[121][10] ), 
	.A1(n6362), 
	.A0(\ram[120][10] ));
   AOI22X1 U11498 (.Y(n13590), 
	.B1(n6381), 
	.B0(\ram[119][10] ), 
	.A1(n6400), 
	.A0(\ram[118][10] ));
   AOI22X1 U11499 (.Y(n13589), 
	.B1(n6419), 
	.B0(\ram[117][10] ), 
	.A1(n6438), 
	.A0(\ram[116][10] ));
   AOI22X1 U11500 (.Y(n13588), 
	.B1(n6457), 
	.B0(\ram[115][10] ), 
	.A1(n6476), 
	.A0(\ram[114][10] ));
   NAND4X1 U11501 (.Y(n13586), 
	.D(n13595), 
	.C(n13594), 
	.B(n13593), 
	.A(n13592));
   AOI22X1 U11502 (.Y(n13595), 
	.B1(n6495), 
	.B0(\ram[113][10] ), 
	.A1(n6514), 
	.A0(\ram[112][10] ));
   AOI22X1 U11503 (.Y(n13594), 
	.B1(n6533), 
	.B0(\ram[127][10] ), 
	.A1(n6553), 
	.A0(\ram[126][10] ));
   AOI22X1 U11504 (.Y(n13593), 
	.B1(n6572), 
	.B0(\ram[125][10] ), 
	.A1(n6591), 
	.A0(\ram[124][10] ));
   AOI22X1 U11505 (.Y(n13592), 
	.B1(n6610), 
	.B0(\ram[123][10] ), 
	.A1(n6629), 
	.A0(\ram[122][10] ));
   OAI21XL U11506 (.Y(n13573), 
	.B0(n9429), 
	.A1(n13597), 
	.A0(n13596));
   NAND4X1 U11507 (.Y(n13597), 
	.D(n13601), 
	.C(n13600), 
	.B(n13599), 
	.A(n13598));
   AOI22X1 U11508 (.Y(n13601), 
	.B1(n6342), 
	.B0(\ram[105][10] ), 
	.A1(n6362), 
	.A0(\ram[104][10] ));
   AOI22X1 U11509 (.Y(n13600), 
	.B1(n6381), 
	.B0(\ram[103][10] ), 
	.A1(n6400), 
	.A0(\ram[102][10] ));
   AOI22X1 U11510 (.Y(n13599), 
	.B1(n6419), 
	.B0(\ram[101][10] ), 
	.A1(n6438), 
	.A0(\ram[100][10] ));
   AOI22X1 U11511 (.Y(n13598), 
	.B1(n6457), 
	.B0(\ram[99][10] ), 
	.A1(n6476), 
	.A0(\ram[98][10] ));
   NAND4X1 U11512 (.Y(n13596), 
	.D(n13605), 
	.C(n13604), 
	.B(n13603), 
	.A(n13602));
   AOI22X1 U11513 (.Y(n13605), 
	.B1(n6495), 
	.B0(\ram[97][10] ), 
	.A1(n6514), 
	.A0(\ram[96][10] ));
   AOI22X1 U11514 (.Y(n13604), 
	.B1(n6533), 
	.B0(\ram[111][10] ), 
	.A1(n6553), 
	.A0(\ram[110][10] ));
   AOI22X1 U11515 (.Y(n13603), 
	.B1(n6572), 
	.B0(\ram[109][10] ), 
	.A1(n6591), 
	.A0(\ram[108][10] ));
   AOI22X1 U11516 (.Y(n13602), 
	.B1(n6610), 
	.B0(\ram[107][10] ), 
	.A1(n6629), 
	.A0(\ram[106][10] ));
   OAI21XL U11517 (.Y(n13572), 
	.B0(n9718), 
	.A1(n13607), 
	.A0(n13606));
   NAND4X1 U11518 (.Y(n13607), 
	.D(n13611), 
	.C(n13610), 
	.B(n13609), 
	.A(n13608));
   AOI22X1 U11519 (.Y(n13611), 
	.B1(n6342), 
	.B0(\ram[89][10] ), 
	.A1(n6362), 
	.A0(\ram[88][10] ));
   AOI22X1 U11520 (.Y(n13610), 
	.B1(n6381), 
	.B0(\ram[87][10] ), 
	.A1(n6400), 
	.A0(\ram[86][10] ));
   AOI22X1 U11521 (.Y(n13609), 
	.B1(n6419), 
	.B0(\ram[85][10] ), 
	.A1(n6438), 
	.A0(\ram[84][10] ));
   AOI22X1 U11522 (.Y(n13608), 
	.B1(n6457), 
	.B0(\ram[83][10] ), 
	.A1(n6476), 
	.A0(\ram[82][10] ));
   NAND4X1 U11523 (.Y(n13606), 
	.D(n13615), 
	.C(n13614), 
	.B(n13613), 
	.A(n13612));
   AOI22X1 U11524 (.Y(n13615), 
	.B1(n6495), 
	.B0(\ram[81][10] ), 
	.A1(n6514), 
	.A0(\ram[80][10] ));
   AOI22X1 U11525 (.Y(n13614), 
	.B1(n6533), 
	.B0(\ram[95][10] ), 
	.A1(n6553), 
	.A0(\ram[94][10] ));
   AOI22X1 U11526 (.Y(n13613), 
	.B1(n6572), 
	.B0(\ram[93][10] ), 
	.A1(n6591), 
	.A0(\ram[92][10] ));
   AOI22X1 U11527 (.Y(n13612), 
	.B1(n6610), 
	.B0(\ram[91][10] ), 
	.A1(n6629), 
	.A0(\ram[90][10] ));
   NAND4X1 U11528 (.Y(n13480), 
	.D(n13619), 
	.C(n13618), 
	.B(n13617), 
	.A(n13616));
   OAI21XL U11529 (.Y(n13619), 
	.B0(n10007), 
	.A1(n13621), 
	.A0(n13620));
   NAND4X1 U11530 (.Y(n13621), 
	.D(n13625), 
	.C(n13624), 
	.B(n13623), 
	.A(n13622));
   AOI22X1 U11531 (.Y(n13625), 
	.B1(n6342), 
	.B0(\ram[73][10] ), 
	.A1(n6362), 
	.A0(\ram[72][10] ));
   AOI22X1 U11532 (.Y(n13624), 
	.B1(n6381), 
	.B0(\ram[71][10] ), 
	.A1(n6400), 
	.A0(\ram[70][10] ));
   AOI22X1 U11533 (.Y(n13623), 
	.B1(n6419), 
	.B0(\ram[69][10] ), 
	.A1(n6438), 
	.A0(\ram[68][10] ));
   AOI22X1 U11534 (.Y(n13622), 
	.B1(n6457), 
	.B0(\ram[67][10] ), 
	.A1(n6476), 
	.A0(\ram[66][10] ));
   NAND4X1 U11535 (.Y(n13620), 
	.D(n13629), 
	.C(n13628), 
	.B(n13627), 
	.A(n13626));
   AOI22X1 U11536 (.Y(n13629), 
	.B1(n6495), 
	.B0(\ram[65][10] ), 
	.A1(n6514), 
	.A0(\ram[64][10] ));
   AOI22X1 U11537 (.Y(n13628), 
	.B1(n6533), 
	.B0(\ram[79][10] ), 
	.A1(n6553), 
	.A0(\ram[78][10] ));
   AOI22X1 U11538 (.Y(n13627), 
	.B1(n6572), 
	.B0(\ram[77][10] ), 
	.A1(n6591), 
	.A0(\ram[76][10] ));
   AOI22X1 U11539 (.Y(n13626), 
	.B1(n6610), 
	.B0(\ram[75][10] ), 
	.A1(n6629), 
	.A0(\ram[74][10] ));
   OAI21XL U11540 (.Y(n13618), 
	.B0(n10296), 
	.A1(n13631), 
	.A0(n13630));
   NAND4X1 U11541 (.Y(n13631), 
	.D(n13635), 
	.C(n13634), 
	.B(n13633), 
	.A(n13632));
   AOI22X1 U11542 (.Y(n13635), 
	.B1(n6342), 
	.B0(\ram[57][10] ), 
	.A1(n6362), 
	.A0(\ram[56][10] ));
   AOI22X1 U11543 (.Y(n13634), 
	.B1(n6381), 
	.B0(\ram[55][10] ), 
	.A1(n6400), 
	.A0(\ram[54][10] ));
   AOI22X1 U11544 (.Y(n13633), 
	.B1(n6419), 
	.B0(\ram[53][10] ), 
	.A1(n6438), 
	.A0(\ram[52][10] ));
   AOI22X1 U11545 (.Y(n13632), 
	.B1(n6457), 
	.B0(\ram[51][10] ), 
	.A1(n6476), 
	.A0(\ram[50][10] ));
   NAND4X1 U11546 (.Y(n13630), 
	.D(n13639), 
	.C(n13638), 
	.B(n13637), 
	.A(n13636));
   AOI22X1 U11547 (.Y(n13639), 
	.B1(n6495), 
	.B0(\ram[49][10] ), 
	.A1(n6514), 
	.A0(\ram[48][10] ));
   AOI22X1 U11548 (.Y(n13638), 
	.B1(n6533), 
	.B0(\ram[63][10] ), 
	.A1(n6553), 
	.A0(\ram[62][10] ));
   AOI22X1 U11549 (.Y(n13637), 
	.B1(n6572), 
	.B0(\ram[61][10] ), 
	.A1(n6591), 
	.A0(\ram[60][10] ));
   AOI22X1 U11550 (.Y(n13636), 
	.B1(n6610), 
	.B0(\ram[59][10] ), 
	.A1(n6629), 
	.A0(\ram[58][10] ));
   OAI21XL U11551 (.Y(n13617), 
	.B0(n10585), 
	.A1(n13641), 
	.A0(n13640));
   NAND4X1 U11552 (.Y(n13641), 
	.D(n13645), 
	.C(n13644), 
	.B(n13643), 
	.A(n13642));
   AOI22X1 U11553 (.Y(n13645), 
	.B1(n6342), 
	.B0(\ram[41][10] ), 
	.A1(n6362), 
	.A0(\ram[40][10] ));
   AOI22X1 U11554 (.Y(n13644), 
	.B1(n6381), 
	.B0(\ram[39][10] ), 
	.A1(n6400), 
	.A0(\ram[38][10] ));
   AOI22X1 U11555 (.Y(n13643), 
	.B1(n6419), 
	.B0(\ram[37][10] ), 
	.A1(n6438), 
	.A0(\ram[36][10] ));
   AOI22X1 U11556 (.Y(n13642), 
	.B1(n6457), 
	.B0(\ram[35][10] ), 
	.A1(n6476), 
	.A0(\ram[34][10] ));
   NAND4X1 U11557 (.Y(n13640), 
	.D(n13649), 
	.C(n13648), 
	.B(n13647), 
	.A(n13646));
   AOI22X1 U11558 (.Y(n13649), 
	.B1(n6495), 
	.B0(\ram[33][10] ), 
	.A1(n6514), 
	.A0(\ram[32][10] ));
   AOI22X1 U11559 (.Y(n13648), 
	.B1(n6533), 
	.B0(\ram[47][10] ), 
	.A1(n6553), 
	.A0(\ram[46][10] ));
   AOI22X1 U11560 (.Y(n13647), 
	.B1(n6572), 
	.B0(\ram[45][10] ), 
	.A1(n6591), 
	.A0(\ram[44][10] ));
   AOI22X1 U11561 (.Y(n13646), 
	.B1(n6610), 
	.B0(\ram[43][10] ), 
	.A1(n6629), 
	.A0(\ram[42][10] ));
   OAI21XL U11562 (.Y(n13616), 
	.B0(n6343), 
	.A1(n13651), 
	.A0(n13650));
   NAND4X1 U11563 (.Y(n13651), 
	.D(n13655), 
	.C(n13654), 
	.B(n13653), 
	.A(n13652));
   AOI22X1 U11564 (.Y(n13655), 
	.B1(n6342), 
	.B0(\ram[25][10] ), 
	.A1(n6362), 
	.A0(\ram[24][10] ));
   AOI22X1 U11565 (.Y(n13654), 
	.B1(n6381), 
	.B0(\ram[23][10] ), 
	.A1(n6400), 
	.A0(\ram[22][10] ));
   AOI22X1 U11566 (.Y(n13653), 
	.B1(n6419), 
	.B0(\ram[21][10] ), 
	.A1(n6438), 
	.A0(\ram[20][10] ));
   AOI22X1 U11567 (.Y(n13652), 
	.B1(n6457), 
	.B0(\ram[19][10] ), 
	.A1(n6476), 
	.A0(\ram[18][10] ));
   NAND4X1 U11568 (.Y(n13650), 
	.D(n13659), 
	.C(n13658), 
	.B(n13657), 
	.A(n13656));
   AOI22X1 U11569 (.Y(n13659), 
	.B1(n6495), 
	.B0(\ram[17][10] ), 
	.A1(n6514), 
	.A0(\ram[16][10] ));
   AOI22X1 U11570 (.Y(n13658), 
	.B1(n6533), 
	.B0(\ram[31][10] ), 
	.A1(n6553), 
	.A0(\ram[30][10] ));
   AOI22X1 U11571 (.Y(n13657), 
	.B1(n6572), 
	.B0(\ram[29][10] ), 
	.A1(n6591), 
	.A0(\ram[28][10] ));
   AOI22X1 U11572 (.Y(n13656), 
	.B1(n6610), 
	.B0(\ram[27][10] ), 
	.A1(n6629), 
	.A0(\ram[26][10] ));
   OR4X1 U11573 (.Y(mem_read_data[0]), 
	.D(n13663), 
	.C(n13662), 
	.B(n13661), 
	.A(n13660));
   NAND4X1 U11574 (.Y(n13663), 
	.D(n13667), 
	.C(n13666), 
	.B(n13665), 
	.A(n13664));
   OAI21XL U11575 (.Y(n13667), 
	.B0(n6534), 
	.A1(n13669), 
	.A0(n13668));
   AND2X1 U11576 (.Y(n6534), 
	.B(n13671), 
	.A(n13670));
   NAND4X1 U11577 (.Y(n13669), 
	.D(n13675), 
	.C(n13674), 
	.B(n13673), 
	.A(n13672));
   AOI22X1 U11578 (.Y(n13675), 
	.B1(n6342), 
	.B0(\ram[9][0] ), 
	.A1(n6362), 
	.A0(\ram[8][0] ));
   AOI22X1 U11579 (.Y(n13674), 
	.B1(n6381), 
	.B0(\ram[7][0] ), 
	.A1(n6400), 
	.A0(\ram[6][0] ));
   AOI22X1 U11580 (.Y(n13673), 
	.B1(n6419), 
	.B0(\ram[5][0] ), 
	.A1(n6438), 
	.A0(\ram[4][0] ));
   AOI22X1 U11581 (.Y(n13672), 
	.B1(n6457), 
	.B0(\ram[3][0] ), 
	.A1(n6476), 
	.A0(\ram[2][0] ));
   NAND4X1 U11582 (.Y(n13668), 
	.D(n13679), 
	.C(n13678), 
	.B(n13677), 
	.A(n13676));
   AOI22X1 U11583 (.Y(n13679), 
	.B1(n6495), 
	.B0(\ram[1][0] ), 
	.A1(n6514), 
	.A0(\ram[0][0] ));
   AOI22X1 U11584 (.Y(n13678), 
	.B1(n6533), 
	.B0(\ram[15][0] ), 
	.A1(n6553), 
	.A0(\ram[14][0] ));
   AOI22X1 U11585 (.Y(n13677), 
	.B1(n6572), 
	.B0(\ram[13][0] ), 
	.A1(n6591), 
	.A0(\ram[12][0] ));
   AOI22X1 U11586 (.Y(n13676), 
	.B1(n6610), 
	.B0(\ram[11][0] ), 
	.A1(n6629), 
	.A0(\ram[10][0] ));
   OAI21XL U11587 (.Y(n13666), 
	.B0(n6828), 
	.A1(n13681), 
	.A0(n13680));
   AND2X1 U11588 (.Y(n6828), 
	.B(n13683), 
	.A(n13682));
   NAND4X1 U11589 (.Y(n13681), 
	.D(n13687), 
	.C(n13686), 
	.B(n13685), 
	.A(n13684));
   AOI22X1 U11590 (.Y(n13687), 
	.B1(n6342), 
	.B0(\ram[249][0] ), 
	.A1(n6362), 
	.A0(\ram[248][0] ));
   AOI22X1 U11591 (.Y(n13686), 
	.B1(n6381), 
	.B0(\ram[247][0] ), 
	.A1(n6400), 
	.A0(\ram[246][0] ));
   AOI22X1 U11592 (.Y(n13685), 
	.B1(n6419), 
	.B0(\ram[245][0] ), 
	.A1(n6438), 
	.A0(\ram[244][0] ));
   AOI22X1 U11593 (.Y(n13684), 
	.B1(n6457), 
	.B0(\ram[243][0] ), 
	.A1(n6476), 
	.A0(\ram[242][0] ));
   NAND4X1 U11594 (.Y(n13680), 
	.D(n13691), 
	.C(n13690), 
	.B(n13689), 
	.A(n13688));
   AOI22X1 U11595 (.Y(n13691), 
	.B1(n6495), 
	.B0(\ram[241][0] ), 
	.A1(n6514), 
	.A0(\ram[240][0] ));
   AOI22X1 U11596 (.Y(n13690), 
	.B1(n6533), 
	.B0(\ram[255][0] ), 
	.A1(n6553), 
	.A0(\ram[254][0] ));
   AOI22X1 U11597 (.Y(n13689), 
	.B1(n6572), 
	.B0(\ram[253][0] ), 
	.A1(n6591), 
	.A0(\ram[252][0] ));
   AOI22X1 U11598 (.Y(n13688), 
	.B1(n6610), 
	.B0(\ram[251][0] ), 
	.A1(n6629), 
	.A0(\ram[250][0] ));
   OAI21XL U11599 (.Y(n13665), 
	.B0(n7117), 
	.A1(n13693), 
	.A0(n13692));
   AND2X1 U11600 (.Y(n7117), 
	.B(n13682), 
	.A(n13694));
   NAND4X1 U11601 (.Y(n13693), 
	.D(n13698), 
	.C(n13697), 
	.B(n13696), 
	.A(n13695));
   AOI22X1 U11602 (.Y(n13698), 
	.B1(n6342), 
	.B0(\ram[233][0] ), 
	.A1(n6362), 
	.A0(\ram[232][0] ));
   AOI22X1 U11603 (.Y(n13697), 
	.B1(n6381), 
	.B0(\ram[231][0] ), 
	.A1(n6400), 
	.A0(\ram[230][0] ));
   AOI22X1 U11604 (.Y(n13696), 
	.B1(n6419), 
	.B0(\ram[229][0] ), 
	.A1(n6438), 
	.A0(\ram[228][0] ));
   AOI22X1 U11605 (.Y(n13695), 
	.B1(n6457), 
	.B0(\ram[227][0] ), 
	.A1(n6476), 
	.A0(\ram[226][0] ));
   NAND4X1 U11606 (.Y(n13692), 
	.D(n13702), 
	.C(n13701), 
	.B(n13700), 
	.A(n13699));
   AOI22X1 U11607 (.Y(n13702), 
	.B1(n6495), 
	.B0(\ram[225][0] ), 
	.A1(n6514), 
	.A0(\ram[224][0] ));
   AOI22X1 U11608 (.Y(n13701), 
	.B1(n6533), 
	.B0(\ram[239][0] ), 
	.A1(n6553), 
	.A0(\ram[238][0] ));
   AOI22X1 U11609 (.Y(n13700), 
	.B1(n6572), 
	.B0(\ram[237][0] ), 
	.A1(n6591), 
	.A0(\ram[236][0] ));
   AOI22X1 U11610 (.Y(n13699), 
	.B1(n6610), 
	.B0(\ram[235][0] ), 
	.A1(n6629), 
	.A0(\ram[234][0] ));
   OAI21XL U11611 (.Y(n13664), 
	.B0(n7406), 
	.A1(n13704), 
	.A0(n13703));
   AND2X1 U11612 (.Y(n7406), 
	.B(n13705), 
	.A(n13682));
   NAND4X1 U11613 (.Y(n13704), 
	.D(n13709), 
	.C(n13708), 
	.B(n13707), 
	.A(n13706));
   AOI22X1 U11614 (.Y(n13709), 
	.B1(n6342), 
	.B0(\ram[217][0] ), 
	.A1(n6362), 
	.A0(\ram[216][0] ));
   AOI22X1 U11615 (.Y(n13708), 
	.B1(n6381), 
	.B0(\ram[215][0] ), 
	.A1(n6400), 
	.A0(\ram[214][0] ));
   AOI22X1 U11616 (.Y(n13707), 
	.B1(n6419), 
	.B0(\ram[213][0] ), 
	.A1(n6438), 
	.A0(\ram[212][0] ));
   AOI22X1 U11617 (.Y(n13706), 
	.B1(n6457), 
	.B0(\ram[211][0] ), 
	.A1(n6476), 
	.A0(\ram[210][0] ));
   NAND4X1 U11618 (.Y(n13703), 
	.D(n13713), 
	.C(n13712), 
	.B(n13711), 
	.A(n13710));
   AOI22X1 U11619 (.Y(n13713), 
	.B1(n6495), 
	.B0(\ram[209][0] ), 
	.A1(n6514), 
	.A0(\ram[208][0] ));
   AOI22X1 U11620 (.Y(n13712), 
	.B1(n6533), 
	.B0(\ram[223][0] ), 
	.A1(n6553), 
	.A0(\ram[222][0] ));
   AOI22X1 U11621 (.Y(n13711), 
	.B1(n6572), 
	.B0(\ram[221][0] ), 
	.A1(n6591), 
	.A0(\ram[220][0] ));
   AOI22X1 U11622 (.Y(n13710), 
	.B1(n6610), 
	.B0(\ram[219][0] ), 
	.A1(n6629), 
	.A0(\ram[218][0] ));
   NAND4X1 U11623 (.Y(n13662), 
	.D(n13717), 
	.C(n13716), 
	.B(n13715), 
	.A(n13714));
   OAI21XL U11624 (.Y(n13717), 
	.B0(n7695), 
	.A1(n13719), 
	.A0(n13718));
   AND2X1 U11625 (.Y(n7695), 
	.B(n13670), 
	.A(n13682));
   NOR2X1 U11626 (.Y(n13682), 
	.B(n13721), 
	.A(n13720));
   NAND4X1 U11627 (.Y(n13719), 
	.D(n13725), 
	.C(n13724), 
	.B(n13723), 
	.A(n13722));
   AOI22X1 U11628 (.Y(n13725), 
	.B1(n6342), 
	.B0(\ram[201][0] ), 
	.A1(n6362), 
	.A0(\ram[200][0] ));
   AOI22X1 U11629 (.Y(n13724), 
	.B1(n6381), 
	.B0(\ram[199][0] ), 
	.A1(n6400), 
	.A0(\ram[198][0] ));
   AOI22X1 U11630 (.Y(n13723), 
	.B1(n6419), 
	.B0(\ram[197][0] ), 
	.A1(n6438), 
	.A0(\ram[196][0] ));
   AOI22X1 U11631 (.Y(n13722), 
	.B1(n6457), 
	.B0(\ram[195][0] ), 
	.A1(n6476), 
	.A0(\ram[194][0] ));
   NAND4X1 U11632 (.Y(n13718), 
	.D(n13729), 
	.C(n13728), 
	.B(n13727), 
	.A(n13726));
   AOI22X1 U11633 (.Y(n13729), 
	.B1(n6495), 
	.B0(\ram[193][0] ), 
	.A1(n6514), 
	.A0(\ram[192][0] ));
   AOI22X1 U11634 (.Y(n13728), 
	.B1(n6533), 
	.B0(\ram[207][0] ), 
	.A1(n6553), 
	.A0(\ram[206][0] ));
   AOI22X1 U11635 (.Y(n13727), 
	.B1(n6572), 
	.B0(\ram[205][0] ), 
	.A1(n6591), 
	.A0(\ram[204][0] ));
   AOI22X1 U11636 (.Y(n13726), 
	.B1(n6610), 
	.B0(\ram[203][0] ), 
	.A1(n6629), 
	.A0(\ram[202][0] ));
   OAI21XL U11637 (.Y(n13716), 
	.B0(n7984), 
	.A1(n13731), 
	.A0(n13730));
   AND2X1 U11638 (.Y(n7984), 
	.B(n13683), 
	.A(n13732));
   NAND4X1 U11639 (.Y(n13731), 
	.D(n13736), 
	.C(n13735), 
	.B(n13734), 
	.A(n13733));
   AOI22X1 U11640 (.Y(n13736), 
	.B1(n6342), 
	.B0(\ram[185][0] ), 
	.A1(n6362), 
	.A0(\ram[184][0] ));
   AOI22X1 U11641 (.Y(n13735), 
	.B1(n6381), 
	.B0(\ram[183][0] ), 
	.A1(n6400), 
	.A0(\ram[182][0] ));
   AOI22X1 U11642 (.Y(n13734), 
	.B1(n6419), 
	.B0(\ram[181][0] ), 
	.A1(n6438), 
	.A0(\ram[180][0] ));
   AOI22X1 U11643 (.Y(n13733), 
	.B1(n6457), 
	.B0(\ram[179][0] ), 
	.A1(n6476), 
	.A0(\ram[178][0] ));
   NAND4X1 U11644 (.Y(n13730), 
	.D(n13740), 
	.C(n13739), 
	.B(n13738), 
	.A(n13737));
   AOI22X1 U11645 (.Y(n13740), 
	.B1(n6495), 
	.B0(\ram[177][0] ), 
	.A1(n6514), 
	.A0(\ram[176][0] ));
   AOI22X1 U11646 (.Y(n13739), 
	.B1(n6533), 
	.B0(\ram[191][0] ), 
	.A1(n6553), 
	.A0(\ram[190][0] ));
   AOI22X1 U11647 (.Y(n13738), 
	.B1(n6572), 
	.B0(\ram[189][0] ), 
	.A1(n6591), 
	.A0(\ram[188][0] ));
   AOI22X1 U11648 (.Y(n13737), 
	.B1(n6610), 
	.B0(\ram[187][0] ), 
	.A1(n6629), 
	.A0(\ram[186][0] ));
   OAI21XL U11649 (.Y(n13715), 
	.B0(n8273), 
	.A1(n13742), 
	.A0(n13741));
   AND2X1 U11650 (.Y(n8273), 
	.B(n13694), 
	.A(n13732));
   NAND4X1 U11651 (.Y(n13742), 
	.D(n13746), 
	.C(n13745), 
	.B(n13744), 
	.A(n13743));
   AOI22X1 U11652 (.Y(n13746), 
	.B1(n6342), 
	.B0(\ram[169][0] ), 
	.A1(n6362), 
	.A0(\ram[168][0] ));
   AOI22X1 U11653 (.Y(n13745), 
	.B1(n6381), 
	.B0(\ram[167][0] ), 
	.A1(n6400), 
	.A0(\ram[166][0] ));
   AOI22X1 U11654 (.Y(n13744), 
	.B1(n6419), 
	.B0(\ram[165][0] ), 
	.A1(n6438), 
	.A0(\ram[164][0] ));
   AOI22X1 U11655 (.Y(n13743), 
	.B1(n6457), 
	.B0(\ram[163][0] ), 
	.A1(n6476), 
	.A0(\ram[162][0] ));
   NAND4X1 U11656 (.Y(n13741), 
	.D(n13750), 
	.C(n13749), 
	.B(n13748), 
	.A(n13747));
   AOI22X1 U11657 (.Y(n13750), 
	.B1(n6495), 
	.B0(\ram[161][0] ), 
	.A1(n6514), 
	.A0(\ram[160][0] ));
   AOI22X1 U11658 (.Y(n13749), 
	.B1(n6533), 
	.B0(\ram[175][0] ), 
	.A1(n6553), 
	.A0(\ram[174][0] ));
   AOI22X1 U11659 (.Y(n13748), 
	.B1(n6572), 
	.B0(\ram[173][0] ), 
	.A1(n6591), 
	.A0(\ram[172][0] ));
   AOI22X1 U11660 (.Y(n13747), 
	.B1(n6610), 
	.B0(\ram[171][0] ), 
	.A1(n6629), 
	.A0(\ram[170][0] ));
   OAI21XL U11661 (.Y(n13714), 
	.B0(n8562), 
	.A1(n13752), 
	.A0(n13751));
   AND2X1 U11662 (.Y(n8562), 
	.B(n13705), 
	.A(n13732));
   NAND4X1 U11663 (.Y(n13752), 
	.D(n13756), 
	.C(n13755), 
	.B(n13754), 
	.A(n13753));
   AOI22X1 U11664 (.Y(n13756), 
	.B1(n6342), 
	.B0(\ram[153][0] ), 
	.A1(n6362), 
	.A0(\ram[152][0] ));
   AOI22X1 U11665 (.Y(n13755), 
	.B1(n6381), 
	.B0(\ram[151][0] ), 
	.A1(n6400), 
	.A0(\ram[150][0] ));
   AOI22X1 U11666 (.Y(n13754), 
	.B1(n6419), 
	.B0(\ram[149][0] ), 
	.A1(n6438), 
	.A0(\ram[148][0] ));
   AOI22X1 U11667 (.Y(n13753), 
	.B1(n6457), 
	.B0(\ram[147][0] ), 
	.A1(n6476), 
	.A0(\ram[146][0] ));
   NAND4X1 U11668 (.Y(n13751), 
	.D(n13760), 
	.C(n13759), 
	.B(n13758), 
	.A(n13757));
   AOI22X1 U11669 (.Y(n13760), 
	.B1(n6495), 
	.B0(\ram[145][0] ), 
	.A1(n6514), 
	.A0(\ram[144][0] ));
   AOI22X1 U11670 (.Y(n13759), 
	.B1(n6533), 
	.B0(\ram[159][0] ), 
	.A1(n6553), 
	.A0(\ram[158][0] ));
   AOI22X1 U11671 (.Y(n13758), 
	.B1(n6572), 
	.B0(\ram[157][0] ), 
	.A1(n6591), 
	.A0(\ram[156][0] ));
   AOI22X1 U11672 (.Y(n13757), 
	.B1(n6610), 
	.B0(\ram[155][0] ), 
	.A1(n6629), 
	.A0(\ram[154][0] ));
   NAND4X1 U11673 (.Y(n13661), 
	.D(n13764), 
	.C(n13763), 
	.B(n13762), 
	.A(n13761));
   OAI21XL U11674 (.Y(n13764), 
	.B0(n8851), 
	.A1(n13766), 
	.A0(n13765));
   AND2X1 U11675 (.Y(n8851), 
	.B(n13670), 
	.A(n13732));
   NOR2X1 U11676 (.Y(n13732), 
	.B(N24), 
	.A(n13720));
   INVX1 U11677 (.Y(n13720), 
	.A(N25));
   NAND4X1 U11678 (.Y(n13766), 
	.D(n13770), 
	.C(n13769), 
	.B(n13768), 
	.A(n13767));
   AOI22X1 U11679 (.Y(n13770), 
	.B1(n6342), 
	.B0(\ram[137][0] ), 
	.A1(n6362), 
	.A0(\ram[136][0] ));
   AOI22X1 U11680 (.Y(n13769), 
	.B1(n6381), 
	.B0(\ram[135][0] ), 
	.A1(n6400), 
	.A0(\ram[134][0] ));
   AOI22X1 U11681 (.Y(n13768), 
	.B1(n6419), 
	.B0(\ram[133][0] ), 
	.A1(n6438), 
	.A0(\ram[132][0] ));
   AOI22X1 U11682 (.Y(n13767), 
	.B1(n6457), 
	.B0(\ram[131][0] ), 
	.A1(n6476), 
	.A0(\ram[130][0] ));
   NAND4X1 U11683 (.Y(n13765), 
	.D(n13774), 
	.C(n13773), 
	.B(n13772), 
	.A(n13771));
   AOI22X1 U11684 (.Y(n13774), 
	.B1(n6495), 
	.B0(\ram[129][0] ), 
	.A1(n6514), 
	.A0(\ram[128][0] ));
   AOI22X1 U11685 (.Y(n13773), 
	.B1(n6533), 
	.B0(\ram[143][0] ), 
	.A1(n6553), 
	.A0(\ram[142][0] ));
   AOI22X1 U11686 (.Y(n13772), 
	.B1(n6572), 
	.B0(\ram[141][0] ), 
	.A1(n6591), 
	.A0(\ram[140][0] ));
   AOI22X1 U11687 (.Y(n13771), 
	.B1(n6610), 
	.B0(\ram[139][0] ), 
	.A1(n6629), 
	.A0(\ram[138][0] ));
   OAI21XL U11688 (.Y(n13763), 
	.B0(n9140), 
	.A1(n13776), 
	.A0(n13775));
   AND2X1 U11689 (.Y(n9140), 
	.B(n13683), 
	.A(n13777));
   NAND4X1 U11690 (.Y(n13776), 
	.D(n13781), 
	.C(n13780), 
	.B(n13779), 
	.A(n13778));
   AOI22X1 U11691 (.Y(n13781), 
	.B1(n6342), 
	.B0(\ram[121][0] ), 
	.A1(n6362), 
	.A0(\ram[120][0] ));
   AOI22X1 U11692 (.Y(n13780), 
	.B1(n6381), 
	.B0(\ram[119][0] ), 
	.A1(n6400), 
	.A0(\ram[118][0] ));
   AOI22X1 U11693 (.Y(n13779), 
	.B1(n6419), 
	.B0(\ram[117][0] ), 
	.A1(n6438), 
	.A0(\ram[116][0] ));
   AOI22X1 U11694 (.Y(n13778), 
	.B1(n6457), 
	.B0(\ram[115][0] ), 
	.A1(n6476), 
	.A0(\ram[114][0] ));
   NAND4X1 U11695 (.Y(n13775), 
	.D(n13785), 
	.C(n13784), 
	.B(n13783), 
	.A(n13782));
   AOI22X1 U11696 (.Y(n13785), 
	.B1(n6495), 
	.B0(\ram[113][0] ), 
	.A1(n6514), 
	.A0(\ram[112][0] ));
   AOI22X1 U11697 (.Y(n13784), 
	.B1(n6533), 
	.B0(\ram[127][0] ), 
	.A1(n6553), 
	.A0(\ram[126][0] ));
   AOI22X1 U11698 (.Y(n13783), 
	.B1(n6572), 
	.B0(\ram[125][0] ), 
	.A1(n6591), 
	.A0(\ram[124][0] ));
   AOI22X1 U11699 (.Y(n13782), 
	.B1(n6610), 
	.B0(\ram[123][0] ), 
	.A1(n6629), 
	.A0(\ram[122][0] ));
   OAI21XL U11700 (.Y(n13762), 
	.B0(n9429), 
	.A1(n13787), 
	.A0(n13786));
   AND2X1 U11701 (.Y(n9429), 
	.B(n13694), 
	.A(n13777));
   NAND4X1 U11702 (.Y(n13787), 
	.D(n13791), 
	.C(n13790), 
	.B(n13789), 
	.A(n13788));
   AOI22X1 U11703 (.Y(n13791), 
	.B1(n6342), 
	.B0(\ram[105][0] ), 
	.A1(n6362), 
	.A0(\ram[104][0] ));
   AOI22X1 U11704 (.Y(n13790), 
	.B1(n6381), 
	.B0(\ram[103][0] ), 
	.A1(n6400), 
	.A0(\ram[102][0] ));
   AOI22X1 U11705 (.Y(n13789), 
	.B1(n6419), 
	.B0(\ram[101][0] ), 
	.A1(n6438), 
	.A0(\ram[100][0] ));
   AOI22X1 U11706 (.Y(n13788), 
	.B1(n6457), 
	.B0(\ram[99][0] ), 
	.A1(n6476), 
	.A0(\ram[98][0] ));
   NAND4X1 U11707 (.Y(n13786), 
	.D(n13795), 
	.C(n13794), 
	.B(n13793), 
	.A(n13792));
   AOI22X1 U11708 (.Y(n13795), 
	.B1(n6495), 
	.B0(\ram[97][0] ), 
	.A1(n6514), 
	.A0(\ram[96][0] ));
   AOI22X1 U11709 (.Y(n13794), 
	.B1(n6533), 
	.B0(\ram[111][0] ), 
	.A1(n6553), 
	.A0(\ram[110][0] ));
   AOI22X1 U11710 (.Y(n13793), 
	.B1(n6572), 
	.B0(\ram[109][0] ), 
	.A1(n6591), 
	.A0(\ram[108][0] ));
   AOI22X1 U11711 (.Y(n13792), 
	.B1(n6610), 
	.B0(\ram[107][0] ), 
	.A1(n6629), 
	.A0(\ram[106][0] ));
   OAI21XL U11712 (.Y(n13761), 
	.B0(n9718), 
	.A1(n13797), 
	.A0(n13796));
   AND2X1 U11713 (.Y(n9718), 
	.B(n13705), 
	.A(n13777));
   NAND4X1 U11714 (.Y(n13797), 
	.D(n13801), 
	.C(n13800), 
	.B(n13799), 
	.A(n13798));
   AOI22X1 U11715 (.Y(n13801), 
	.B1(n6342), 
	.B0(\ram[89][0] ), 
	.A1(n6362), 
	.A0(\ram[88][0] ));
   AOI22X1 U11716 (.Y(n13800), 
	.B1(n6381), 
	.B0(\ram[87][0] ), 
	.A1(n6400), 
	.A0(\ram[86][0] ));
   AOI22X1 U11717 (.Y(n13799), 
	.B1(n6419), 
	.B0(\ram[85][0] ), 
	.A1(n6438), 
	.A0(\ram[84][0] ));
   AOI22X1 U11718 (.Y(n13798), 
	.B1(n6457), 
	.B0(\ram[83][0] ), 
	.A1(n6476), 
	.A0(\ram[82][0] ));
   NAND4X1 U11719 (.Y(n13796), 
	.D(n13805), 
	.C(n13804), 
	.B(n13803), 
	.A(n13802));
   AOI22X1 U11720 (.Y(n13805), 
	.B1(n6495), 
	.B0(\ram[81][0] ), 
	.A1(n6514), 
	.A0(\ram[80][0] ));
   AOI22X1 U11721 (.Y(n13804), 
	.B1(n6533), 
	.B0(\ram[95][0] ), 
	.A1(n6553), 
	.A0(\ram[94][0] ));
   AOI22X1 U11722 (.Y(n13803), 
	.B1(n6572), 
	.B0(\ram[93][0] ), 
	.A1(n6591), 
	.A0(\ram[92][0] ));
   AOI22X1 U11723 (.Y(n13802), 
	.B1(n6610), 
	.B0(\ram[91][0] ), 
	.A1(n6629), 
	.A0(\ram[90][0] ));
   NAND4X1 U11724 (.Y(n13660), 
	.D(n13809), 
	.C(n13808), 
	.B(n13807), 
	.A(n13806));
   OAI21XL U11725 (.Y(n13809), 
	.B0(n10007), 
	.A1(n13811), 
	.A0(n13810));
   AND2X1 U11726 (.Y(n10007), 
	.B(n13670), 
	.A(n13777));
   NOR2X1 U11727 (.Y(n13670), 
	.B(N23), 
	.A(N22));
   NOR2X1 U11728 (.Y(n13777), 
	.B(N25), 
	.A(n13721));
   INVX1 U11729 (.Y(n13721), 
	.A(N24));
   NAND4X1 U11730 (.Y(n13811), 
	.D(n13815), 
	.C(n13814), 
	.B(n13813), 
	.A(n13812));
   AOI22X1 U11731 (.Y(n13815), 
	.B1(n6342), 
	.B0(\ram[73][0] ), 
	.A1(n6362), 
	.A0(\ram[72][0] ));
   AOI22X1 U11732 (.Y(n13814), 
	.B1(n6381), 
	.B0(\ram[71][0] ), 
	.A1(n6400), 
	.A0(\ram[70][0] ));
   AOI22X1 U11733 (.Y(n13813), 
	.B1(n6419), 
	.B0(\ram[69][0] ), 
	.A1(n6438), 
	.A0(\ram[68][0] ));
   AOI22X1 U11734 (.Y(n13812), 
	.B1(n6457), 
	.B0(\ram[67][0] ), 
	.A1(n6476), 
	.A0(\ram[66][0] ));
   NAND4X1 U11735 (.Y(n13810), 
	.D(n13819), 
	.C(n13818), 
	.B(n13817), 
	.A(n13816));
   AOI22X1 U11736 (.Y(n13819), 
	.B1(n6495), 
	.B0(\ram[65][0] ), 
	.A1(n6514), 
	.A0(\ram[64][0] ));
   AOI22X1 U11737 (.Y(n13818), 
	.B1(n6533), 
	.B0(\ram[79][0] ), 
	.A1(n6553), 
	.A0(\ram[78][0] ));
   AOI22X1 U11738 (.Y(n13817), 
	.B1(n6572), 
	.B0(\ram[77][0] ), 
	.A1(n6591), 
	.A0(\ram[76][0] ));
   AOI22X1 U11739 (.Y(n13816), 
	.B1(n6610), 
	.B0(\ram[75][0] ), 
	.A1(n6629), 
	.A0(\ram[74][0] ));
   OAI21XL U11740 (.Y(n13808), 
	.B0(n10296), 
	.A1(n13821), 
	.A0(n13820));
   AND2X1 U11741 (.Y(n10296), 
	.B(n13671), 
	.A(n13683));
   AND2X1 U11742 (.Y(n13683), 
	.B(N22), 
	.A(N23));
   NAND4X1 U11743 (.Y(n13821), 
	.D(n13825), 
	.C(n13824), 
	.B(n13823), 
	.A(n13822));
   AOI22X1 U11744 (.Y(n13825), 
	.B1(n6342), 
	.B0(\ram[57][0] ), 
	.A1(n6362), 
	.A0(\ram[56][0] ));
   AOI22X1 U11745 (.Y(n13824), 
	.B1(n6381), 
	.B0(\ram[55][0] ), 
	.A1(n6400), 
	.A0(\ram[54][0] ));
   AOI22X1 U11746 (.Y(n13823), 
	.B1(n6419), 
	.B0(\ram[53][0] ), 
	.A1(n6438), 
	.A0(\ram[52][0] ));
   AOI22X1 U11747 (.Y(n13822), 
	.B1(n6457), 
	.B0(\ram[51][0] ), 
	.A1(n6476), 
	.A0(\ram[50][0] ));
   NAND4X1 U11748 (.Y(n13820), 
	.D(n13829), 
	.C(n13828), 
	.B(n13827), 
	.A(n13826));
   AOI22X1 U11749 (.Y(n13829), 
	.B1(n6495), 
	.B0(\ram[49][0] ), 
	.A1(n6514), 
	.A0(\ram[48][0] ));
   AOI22X1 U11750 (.Y(n13828), 
	.B1(n6533), 
	.B0(\ram[63][0] ), 
	.A1(n6553), 
	.A0(\ram[62][0] ));
   AOI22X1 U11751 (.Y(n13827), 
	.B1(n6572), 
	.B0(\ram[61][0] ), 
	.A1(n6591), 
	.A0(\ram[60][0] ));
   AOI22X1 U11752 (.Y(n13826), 
	.B1(n6610), 
	.B0(\ram[59][0] ), 
	.A1(n6629), 
	.A0(\ram[58][0] ));
   OAI21XL U11753 (.Y(n13807), 
	.B0(n10585), 
	.A1(n13831), 
	.A0(n13830));
   AND2X1 U11754 (.Y(n10585), 
	.B(n13671), 
	.A(n13694));
   AND2X1 U11755 (.Y(n13694), 
	.B(n13832), 
	.A(N23));
   NAND4X1 U11756 (.Y(n13831), 
	.D(n13836), 
	.C(n13835), 
	.B(n13834), 
	.A(n13833));
   AOI22X1 U11757 (.Y(n13836), 
	.B1(n6342), 
	.B0(\ram[41][0] ), 
	.A1(n6362), 
	.A0(\ram[40][0] ));
   AOI22X1 U11758 (.Y(n13835), 
	.B1(n6381), 
	.B0(\ram[39][0] ), 
	.A1(n6400), 
	.A0(\ram[38][0] ));
   AOI22X1 U11759 (.Y(n13834), 
	.B1(n6419), 
	.B0(\ram[37][0] ), 
	.A1(n6438), 
	.A0(\ram[36][0] ));
   AOI22X1 U11760 (.Y(n13833), 
	.B1(n6457), 
	.B0(\ram[35][0] ), 
	.A1(n6476), 
	.A0(\ram[34][0] ));
   NAND4X1 U11761 (.Y(n13830), 
	.D(n13840), 
	.C(n13839), 
	.B(n13838), 
	.A(n13837));
   AOI22X1 U11762 (.Y(n13840), 
	.B1(n6495), 
	.B0(\ram[33][0] ), 
	.A1(n6514), 
	.A0(\ram[32][0] ));
   AOI22X1 U11763 (.Y(n13839), 
	.B1(n6533), 
	.B0(\ram[47][0] ), 
	.A1(n6553), 
	.A0(\ram[46][0] ));
   AOI22X1 U11764 (.Y(n13838), 
	.B1(n6572), 
	.B0(\ram[45][0] ), 
	.A1(n6591), 
	.A0(\ram[44][0] ));
   AOI22X1 U11765 (.Y(n13837), 
	.B1(n6610), 
	.B0(\ram[43][0] ), 
	.A1(n6629), 
	.A0(\ram[42][0] ));
   OAI21XL U11766 (.Y(n13806), 
	.B0(n6343), 
	.A1(n13842), 
	.A0(n13841));
   AND2X1 U11767 (.Y(n6343), 
	.B(n13705), 
	.A(n13671));
   NOR2X1 U11768 (.Y(n13705), 
	.B(N23), 
	.A(n13832));
   INVX1 U11769 (.Y(n13832), 
	.A(N22));
   NOR2X1 U11770 (.Y(n13671), 
	.B(N25), 
	.A(N24));
   NAND4X1 U11771 (.Y(n13842), 
	.D(n13846), 
	.C(n13845), 
	.B(n13844), 
	.A(n13843));
   AOI22X1 U11772 (.Y(n13846), 
	.B1(n6342), 
	.B0(\ram[25][0] ), 
	.A1(n6362), 
	.A0(\ram[24][0] ));
   AND2X1 U11773 (.Y(n6342), 
	.B(n13848), 
	.A(n13847));
   AND2X1 U11774 (.Y(n6362), 
	.B(n13848), 
	.A(n13849));
   AOI22X1 U11775 (.Y(n13845), 
	.B1(n6381), 
	.B0(\ram[23][0] ), 
	.A1(n6400), 
	.A0(\ram[22][0] ));
   AND2X1 U11776 (.Y(n6381), 
	.B(n13851), 
	.A(n13850));
   AND2X1 U11777 (.Y(n6400), 
	.B(n13852), 
	.A(n13850));
   AOI22X1 U11778 (.Y(n13844), 
	.B1(n6419), 
	.B0(\ram[21][0] ), 
	.A1(n6438), 
	.A0(\ram[20][0] ));
   AND2X1 U11779 (.Y(n6419), 
	.B(n13847), 
	.A(n13850));
   AND2X1 U11780 (.Y(n6438), 
	.B(n13849), 
	.A(n13850));
   NOR2X1 U11781 (.Y(n13850), 
	.B(N21), 
	.A(n13853));
   AOI22X1 U11782 (.Y(n13843), 
	.B1(n6457), 
	.B0(\ram[19][0] ), 
	.A1(n6476), 
	.A0(\ram[18][0] ));
   AND2X1 U11783 (.Y(n6457), 
	.B(n13851), 
	.A(n13854));
   AND2X1 U11784 (.Y(n6476), 
	.B(n13852), 
	.A(n13854));
   NAND4X1 U11785 (.Y(n13841), 
	.D(n13858), 
	.C(n13857), 
	.B(n13856), 
	.A(n13855));
   AOI22X1 U11786 (.Y(n13858), 
	.B1(n6495), 
	.B0(\ram[17][0] ), 
	.A1(n6514), 
	.A0(\ram[16][0] ));
   AND2X1 U11787 (.Y(n6495), 
	.B(n13847), 
	.A(n13854));
   AND2X1 U11788 (.Y(n6514), 
	.B(n13849), 
	.A(n13854));
   NOR2X1 U11789 (.Y(n13854), 
	.B(N21), 
	.A(N20));
   AOI22X1 U11790 (.Y(n13857), 
	.B1(n6533), 
	.B0(\ram[31][0] ), 
	.A1(n6553), 
	.A0(\ram[30][0] ));
   AND2X1 U11791 (.Y(n6533), 
	.B(n13851), 
	.A(n13859));
   AND2X1 U11792 (.Y(n6553), 
	.B(n13852), 
	.A(n13859));
   AOI22X1 U11793 (.Y(n13856), 
	.B1(n6572), 
	.B0(\ram[29][0] ), 
	.A1(n6591), 
	.A0(\ram[28][0] ));
   AND2X1 U11794 (.Y(n6572), 
	.B(n13847), 
	.A(n13859));
   NOR2X1 U11795 (.Y(n13847), 
	.B(N19), 
	.A(n13860));
   AND2X1 U11796 (.Y(n6591), 
	.B(n13849), 
	.A(n13859));
   NOR2X1 U11797 (.Y(n13849), 
	.B(N19), 
	.A(N18));
   NOR2X1 U11798 (.Y(n13859), 
	.B(n13861), 
	.A(n13853));
   INVX1 U11799 (.Y(n13853), 
	.A(N20));
   AOI22X1 U11800 (.Y(n13855), 
	.B1(n6610), 
	.B0(\ram[27][0] ), 
	.A1(n6629), 
	.A0(\ram[26][0] ));
   AND2X1 U11801 (.Y(n6610), 
	.B(n13848), 
	.A(n13851));
   NOR2X1 U11802 (.Y(n13851), 
	.B(n13862), 
	.A(n13860));
   INVX1 U11803 (.Y(n13860), 
	.A(N18));
   AND2X1 U11804 (.Y(n6629), 
	.B(n13852), 
	.A(n13848));
   NOR2X1 U11805 (.Y(n13852), 
	.B(N18), 
	.A(n13862));
   INVX1 U11806 (.Y(n13862), 
	.A(N19));
   NOR2X1 U11807 (.Y(n13848), 
	.B(N20), 
	.A(n13861));
   INVX1 U11808 (.Y(n13861), 
	.A(N21));
endmodule

module MEM_stage (
	clk, 
	rst, 
	pipeline_reg_in, 
	pipeline_reg_out, 
	mem_op_dest);
   input clk;
   input rst;
   input [37:0] pipeline_reg_in;
   output [36:0] pipeline_reg_out;
   output [2:0] mem_op_dest;

   // Internal wires
   wire pipeline_reg_in_0;
   wire \pipeline_reg_in[3] ;
   wire \pipeline_reg_in[2] ;
   wire \pipeline_reg_in[1] ;
   wire n76;
   wire [15:0] mem_read_data;

   assign pipeline_reg_in_0 = pipeline_reg_in[0] ;
   assign mem_op_dest[2] = \pipeline_reg_in[3]  ;
   assign \pipeline_reg_in[3]  = pipeline_reg_in[3] ;
   assign mem_op_dest[1] = \pipeline_reg_in[2]  ;
   assign \pipeline_reg_in[2]  = pipeline_reg_in[2] ;
   assign mem_op_dest[0] = \pipeline_reg_in[1]  ;
   assign \pipeline_reg_in[1]  = pipeline_reg_in[1] ;

   data_mem dmem (.clk(clk), 
	.mem_access_addr({ pipeline_reg_in[37],
		pipeline_reg_in[36],
		pipeline_reg_in[35],
		pipeline_reg_in[34],
		pipeline_reg_in[33],
		pipeline_reg_in[32],
		pipeline_reg_in[31],
		pipeline_reg_in[30],
		pipeline_reg_in[29],
		pipeline_reg_in[28],
		pipeline_reg_in[27],
		pipeline_reg_in[26],
		pipeline_reg_in[25],
		pipeline_reg_in[24],
		pipeline_reg_in[23],
		pipeline_reg_in[22] }), 
	.mem_write_data({ pipeline_reg_in[20],
		pipeline_reg_in[19],
		pipeline_reg_in[18],
		pipeline_reg_in[17],
		pipeline_reg_in[16],
		pipeline_reg_in[15],
		pipeline_reg_in[14],
		pipeline_reg_in[13],
		pipeline_reg_in[12],
		pipeline_reg_in[11],
		pipeline_reg_in[10],
		pipeline_reg_in[9],
		pipeline_reg_in[8],
		pipeline_reg_in[7],
		pipeline_reg_in[6],
		pipeline_reg_in[5] }), 
	.mem_write_en(pipeline_reg_in[21]), 
	.mem_read_data({ mem_read_data[15],
		mem_read_data[14],
		mem_read_data[13],
		mem_read_data[12],
		mem_read_data[11],
		mem_read_data[10],
		mem_read_data[9],
		mem_read_data[8],
		mem_read_data[7],
		mem_read_data[6],
		mem_read_data[5],
		mem_read_data[4],
		mem_read_data[3],
		mem_read_data[2],
		mem_read_data[1],
		mem_read_data[0] }));
   DFFTRX1 \pipeline_reg_out_reg[20]  (.RN(n76), 
	.Q(pipeline_reg_out[20]), 
	.D(mem_read_data[15]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[19]  (.RN(n76), 
	.Q(pipeline_reg_out[19]), 
	.D(mem_read_data[14]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[18]  (.RN(n76), 
	.Q(pipeline_reg_out[18]), 
	.D(mem_read_data[13]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[17]  (.RN(n76), 
	.Q(pipeline_reg_out[17]), 
	.D(mem_read_data[12]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[16]  (.RN(n76), 
	.Q(pipeline_reg_out[16]), 
	.D(mem_read_data[11]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[15]  (.RN(n76), 
	.Q(pipeline_reg_out[15]), 
	.D(mem_read_data[10]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[14]  (.RN(n76), 
	.Q(pipeline_reg_out[14]), 
	.D(mem_read_data[9]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[13]  (.RN(n76), 
	.Q(pipeline_reg_out[13]), 
	.D(mem_read_data[8]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[12]  (.RN(n76), 
	.Q(pipeline_reg_out[12]), 
	.D(mem_read_data[7]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[11]  (.RN(n76), 
	.Q(pipeline_reg_out[11]), 
	.D(mem_read_data[6]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[10]  (.RN(n76), 
	.Q(pipeline_reg_out[10]), 
	.D(mem_read_data[5]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[9]  (.RN(n76), 
	.Q(pipeline_reg_out[9]), 
	.D(mem_read_data[4]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[8]  (.RN(n76), 
	.Q(pipeline_reg_out[8]), 
	.D(mem_read_data[3]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[7]  (.RN(n76), 
	.Q(pipeline_reg_out[7]), 
	.D(mem_read_data[2]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[6]  (.RN(n76), 
	.Q(pipeline_reg_out[6]), 
	.D(mem_read_data[1]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[5]  (.RN(n76), 
	.Q(pipeline_reg_out[5]), 
	.D(mem_read_data[0]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[36]  (.RN(n76), 
	.Q(pipeline_reg_out[36]), 
	.D(pipeline_reg_in[37]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[35]  (.RN(n76), 
	.Q(pipeline_reg_out[35]), 
	.D(pipeline_reg_in[36]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[34]  (.RN(n76), 
	.Q(pipeline_reg_out[34]), 
	.D(pipeline_reg_in[35]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[33]  (.RN(n76), 
	.Q(pipeline_reg_out[33]), 
	.D(pipeline_reg_in[34]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[32]  (.RN(n76), 
	.Q(pipeline_reg_out[32]), 
	.D(pipeline_reg_in[33]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[31]  (.RN(n76), 
	.Q(pipeline_reg_out[31]), 
	.D(pipeline_reg_in[32]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[30]  (.RN(n76), 
	.Q(pipeline_reg_out[30]), 
	.D(pipeline_reg_in[31]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[29]  (.RN(n76), 
	.Q(pipeline_reg_out[29]), 
	.D(pipeline_reg_in[30]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[28]  (.RN(n76), 
	.Q(pipeline_reg_out[28]), 
	.D(pipeline_reg_in[29]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[27]  (.RN(n76), 
	.Q(pipeline_reg_out[27]), 
	.D(pipeline_reg_in[28]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[26]  (.RN(n76), 
	.Q(pipeline_reg_out[26]), 
	.D(pipeline_reg_in[27]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[25]  (.RN(n76), 
	.Q(pipeline_reg_out[25]), 
	.D(pipeline_reg_in[26]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[24]  (.RN(n76), 
	.Q(pipeline_reg_out[24]), 
	.D(pipeline_reg_in[25]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[23]  (.RN(n76), 
	.Q(pipeline_reg_out[23]), 
	.D(pipeline_reg_in[24]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[22]  (.RN(n76), 
	.Q(pipeline_reg_out[22]), 
	.D(pipeline_reg_in[23]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[21]  (.RN(n76), 
	.Q(pipeline_reg_out[21]), 
	.D(pipeline_reg_in[22]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[4]  (.RN(n76), 
	.Q(pipeline_reg_out[4]), 
	.D(pipeline_reg_in[4]), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[2]  (.RN(n76), 
	.Q(pipeline_reg_out[2]), 
	.D(\pipeline_reg_in[2] ), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[3]  (.RN(n76), 
	.Q(pipeline_reg_out[3]), 
	.D(\pipeline_reg_in[3] ), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[1]  (.RN(n76), 
	.Q(pipeline_reg_out[1]), 
	.D(\pipeline_reg_in[1] ), 
	.CK(clk));
   DFFTRX1 \pipeline_reg_out_reg[0]  (.RN(n76), 
	.Q(pipeline_reg_out[0]), 
	.D(pipeline_reg_in_0), 
	.CK(clk));
   INVX1 U3 (.Y(n76), 
	.A(rst));
endmodule

module WB_stage (
	pipeline_reg_in, 
	reg_write_en, 
	reg_write_dest, 
	reg_write_data, 
	wb_op_dest);
   input [36:0] pipeline_reg_in;
   output reg_write_en;
   output [2:0] reg_write_dest;
   output [15:0] reg_write_data;
   output [2:0] wb_op_dest;

   // Internal wires
   wire pipeline_reg_in_0;
   wire \pipeline_reg_in[3] ;
   wire \pipeline_reg_in[2] ;
   wire \pipeline_reg_in[1] ;

   assign reg_write_en = pipeline_reg_in[4] ;
   assign pipeline_reg_in_0 = pipeline_reg_in[0] ;
   assign wb_op_dest[2] = \pipeline_reg_in[3]  ;
   assign reg_write_dest[2] = \pipeline_reg_in[3]  ;
   assign \pipeline_reg_in[3]  = pipeline_reg_in[3] ;
   assign wb_op_dest[1] = \pipeline_reg_in[2]  ;
   assign reg_write_dest[1] = \pipeline_reg_in[2]  ;
   assign \pipeline_reg_in[2]  = pipeline_reg_in[2] ;
   assign wb_op_dest[0] = \pipeline_reg_in[1]  ;
   assign reg_write_dest[0] = \pipeline_reg_in[1]  ;
   assign \pipeline_reg_in[1]  = pipeline_reg_in[1] ;

   MX2X1 U1 (.Y(reg_write_data[15]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[20]), 
	.A(pipeline_reg_in[36]));
   MX2X1 U2 (.Y(reg_write_data[14]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[19]), 
	.A(pipeline_reg_in[35]));
   MX2X1 U3 (.Y(reg_write_data[13]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[18]), 
	.A(pipeline_reg_in[34]));
   MX2X1 U4 (.Y(reg_write_data[12]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[17]), 
	.A(pipeline_reg_in[33]));
   MX2X1 U5 (.Y(reg_write_data[11]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[16]), 
	.A(pipeline_reg_in[32]));
   MX2X1 U6 (.Y(reg_write_data[10]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[15]), 
	.A(pipeline_reg_in[31]));
   MX2X1 U7 (.Y(reg_write_data[9]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[14]), 
	.A(pipeline_reg_in[30]));
   MX2X1 U8 (.Y(reg_write_data[8]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[13]), 
	.A(pipeline_reg_in[29]));
   MX2X1 U9 (.Y(reg_write_data[7]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[12]), 
	.A(pipeline_reg_in[28]));
   MX2X1 U10 (.Y(reg_write_data[6]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[11]), 
	.A(pipeline_reg_in[27]));
   MX2X1 U11 (.Y(reg_write_data[5]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[10]), 
	.A(pipeline_reg_in[26]));
   MX2X1 U12 (.Y(reg_write_data[4]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[9]), 
	.A(pipeline_reg_in[25]));
   MX2X1 U13 (.Y(reg_write_data[3]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[8]), 
	.A(pipeline_reg_in[24]));
   MX2X1 U14 (.Y(reg_write_data[2]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[7]), 
	.A(pipeline_reg_in[23]));
   MX2X1 U15 (.Y(reg_write_data[1]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[6]), 
	.A(pipeline_reg_in[22]));
   MX2X1 U16 (.Y(reg_write_data[0]), 
	.S0(pipeline_reg_in_0), 
	.B(pipeline_reg_in[5]), 
	.A(pipeline_reg_in[21]));
endmodule

module register_file (
	clk, 
	rst, 
	reg_write_en, 
	reg_write_dest, 
	reg_write_data, 
	reg_read_addr_1, 
	reg_read_data_1, 
	reg_read_addr_2, 
	reg_read_data_2);
   input clk;
   input rst;
   input reg_write_en;
   input [2:0] reg_write_dest;
   input [15:0] reg_write_data;
   input [2:0] reg_read_addr_1;
   output [15:0] reg_read_data_1;
   input [2:0] reg_read_addr_2;
   output [15:0] reg_read_data_2;

   // Internal wires
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire \reg_array[7][15] ;
   wire \reg_array[7][14] ;
   wire \reg_array[7][13] ;
   wire \reg_array[7][12] ;
   wire \reg_array[7][11] ;
   wire \reg_array[7][10] ;
   wire \reg_array[7][9] ;
   wire \reg_array[7][8] ;
   wire \reg_array[7][7] ;
   wire \reg_array[7][6] ;
   wire \reg_array[7][5] ;
   wire \reg_array[7][4] ;
   wire \reg_array[7][3] ;
   wire \reg_array[7][2] ;
   wire \reg_array[7][1] ;
   wire \reg_array[7][0] ;
   wire \reg_array[6][15] ;
   wire \reg_array[6][14] ;
   wire \reg_array[6][13] ;
   wire \reg_array[6][12] ;
   wire \reg_array[6][11] ;
   wire \reg_array[6][10] ;
   wire \reg_array[6][9] ;
   wire \reg_array[6][8] ;
   wire \reg_array[6][7] ;
   wire \reg_array[6][6] ;
   wire \reg_array[6][5] ;
   wire \reg_array[6][4] ;
   wire \reg_array[6][3] ;
   wire \reg_array[6][2] ;
   wire \reg_array[6][1] ;
   wire \reg_array[6][0] ;
   wire \reg_array[5][15] ;
   wire \reg_array[5][14] ;
   wire \reg_array[5][13] ;
   wire \reg_array[5][12] ;
   wire \reg_array[5][11] ;
   wire \reg_array[5][10] ;
   wire \reg_array[5][9] ;
   wire \reg_array[5][8] ;
   wire \reg_array[5][7] ;
   wire \reg_array[5][6] ;
   wire \reg_array[5][5] ;
   wire \reg_array[5][4] ;
   wire \reg_array[5][3] ;
   wire \reg_array[5][2] ;
   wire \reg_array[5][1] ;
   wire \reg_array[5][0] ;
   wire \reg_array[4][15] ;
   wire \reg_array[4][14] ;
   wire \reg_array[4][13] ;
   wire \reg_array[4][12] ;
   wire \reg_array[4][11] ;
   wire \reg_array[4][10] ;
   wire \reg_array[4][9] ;
   wire \reg_array[4][8] ;
   wire \reg_array[4][7] ;
   wire \reg_array[4][6] ;
   wire \reg_array[4][5] ;
   wire \reg_array[4][4] ;
   wire \reg_array[4][3] ;
   wire \reg_array[4][2] ;
   wire \reg_array[4][1] ;
   wire \reg_array[4][0] ;
   wire \reg_array[3][15] ;
   wire \reg_array[3][14] ;
   wire \reg_array[3][13] ;
   wire \reg_array[3][12] ;
   wire \reg_array[3][11] ;
   wire \reg_array[3][10] ;
   wire \reg_array[3][9] ;
   wire \reg_array[3][8] ;
   wire \reg_array[3][7] ;
   wire \reg_array[3][6] ;
   wire \reg_array[3][5] ;
   wire \reg_array[3][4] ;
   wire \reg_array[3][3] ;
   wire \reg_array[3][2] ;
   wire \reg_array[3][1] ;
   wire \reg_array[3][0] ;
   wire \reg_array[2][15] ;
   wire \reg_array[2][14] ;
   wire \reg_array[2][13] ;
   wire \reg_array[2][12] ;
   wire \reg_array[2][11] ;
   wire \reg_array[2][10] ;
   wire \reg_array[2][9] ;
   wire \reg_array[2][8] ;
   wire \reg_array[2][7] ;
   wire \reg_array[2][6] ;
   wire \reg_array[2][5] ;
   wire \reg_array[2][4] ;
   wire \reg_array[2][3] ;
   wire \reg_array[2][2] ;
   wire \reg_array[2][1] ;
   wire \reg_array[2][0] ;
   wire \reg_array[1][15] ;
   wire \reg_array[1][14] ;
   wire \reg_array[1][13] ;
   wire \reg_array[1][12] ;
   wire \reg_array[1][11] ;
   wire \reg_array[1][10] ;
   wire \reg_array[1][9] ;
   wire \reg_array[1][8] ;
   wire \reg_array[1][7] ;
   wire \reg_array[1][6] ;
   wire \reg_array[1][5] ;
   wire \reg_array[1][4] ;
   wire \reg_array[1][3] ;
   wire \reg_array[1][2] ;
   wire \reg_array[1][1] ;
   wire \reg_array[1][0] ;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;

   assign N18 = reg_read_addr_1[0] ;
   assign N19 = reg_read_addr_1[1] ;
   assign N20 = reg_read_addr_1[2] ;
   assign N21 = reg_read_addr_2[0] ;
   assign N22 = reg_read_addr_2[1] ;
   assign N23 = reg_read_addr_2[2] ;

   DFFRHQXL \reg_array_reg[5][15]  (.RN(n452), 
	.Q(\reg_array[5][15] ), 
	.D(n340), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][14]  (.RN(n452), 
	.Q(\reg_array[5][14] ), 
	.D(n341), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][13]  (.RN(n452), 
	.Q(\reg_array[5][13] ), 
	.D(n342), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][12]  (.RN(n452), 
	.Q(\reg_array[5][12] ), 
	.D(n343), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][11]  (.RN(n452), 
	.Q(\reg_array[5][11] ), 
	.D(n344), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][10]  (.RN(n452), 
	.Q(\reg_array[5][10] ), 
	.D(n345), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][9]  (.RN(n452), 
	.Q(\reg_array[5][9] ), 
	.D(n346), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][8]  (.RN(n452), 
	.Q(\reg_array[5][8] ), 
	.D(n347), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][7]  (.RN(n452), 
	.Q(\reg_array[5][7] ), 
	.D(n348), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][6]  (.RN(n452), 
	.Q(\reg_array[5][6] ), 
	.D(n349), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][5]  (.RN(n452), 
	.Q(\reg_array[5][5] ), 
	.D(n350), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][4]  (.RN(n452), 
	.Q(\reg_array[5][4] ), 
	.D(n351), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][3]  (.RN(n452), 
	.Q(\reg_array[5][3] ), 
	.D(n352), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][2]  (.RN(n452), 
	.Q(\reg_array[5][2] ), 
	.D(n353), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][1]  (.RN(n452), 
	.Q(\reg_array[5][1] ), 
	.D(n354), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[5][0]  (.RN(n452), 
	.Q(\reg_array[5][0] ), 
	.D(n355), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][15]  (.RN(n452), 
	.Q(\reg_array[4][15] ), 
	.D(n404), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][14]  (.RN(n452), 
	.Q(\reg_array[4][14] ), 
	.D(n405), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][13]  (.RN(n452), 
	.Q(\reg_array[4][13] ), 
	.D(n406), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][12]  (.RN(n452), 
	.Q(\reg_array[4][12] ), 
	.D(n407), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][11]  (.RN(n452), 
	.Q(\reg_array[4][11] ), 
	.D(n408), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][10]  (.RN(n452), 
	.Q(\reg_array[4][10] ), 
	.D(n409), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][9]  (.RN(n452), 
	.Q(\reg_array[4][9] ), 
	.D(n410), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][8]  (.RN(n452), 
	.Q(\reg_array[4][8] ), 
	.D(n411), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][7]  (.RN(n452), 
	.Q(\reg_array[4][7] ), 
	.D(n412), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][6]  (.RN(n452), 
	.Q(\reg_array[4][6] ), 
	.D(n413), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][5]  (.RN(n452), 
	.Q(\reg_array[4][5] ), 
	.D(n414), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][4]  (.RN(n452), 
	.Q(\reg_array[4][4] ), 
	.D(n415), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][3]  (.RN(n452), 
	.Q(\reg_array[4][3] ), 
	.D(n416), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][2]  (.RN(n452), 
	.Q(\reg_array[4][2] ), 
	.D(n417), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][1]  (.RN(n452), 
	.Q(\reg_array[4][1] ), 
	.D(n418), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[4][0]  (.RN(n452), 
	.Q(\reg_array[4][0] ), 
	.D(n419), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][15]  (.RN(n452), 
	.Q(\reg_array[1][15] ), 
	.D(n356), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][14]  (.RN(n452), 
	.Q(\reg_array[1][14] ), 
	.D(n357), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][13]  (.RN(n452), 
	.Q(\reg_array[1][13] ), 
	.D(n358), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][12]  (.RN(n452), 
	.Q(\reg_array[1][12] ), 
	.D(n359), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][11]  (.RN(n452), 
	.Q(\reg_array[1][11] ), 
	.D(n360), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][10]  (.RN(n452), 
	.Q(\reg_array[1][10] ), 
	.D(n361), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][9]  (.RN(n452), 
	.Q(\reg_array[1][9] ), 
	.D(n362), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][8]  (.RN(n452), 
	.Q(\reg_array[1][8] ), 
	.D(n363), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][7]  (.RN(n452), 
	.Q(\reg_array[1][7] ), 
	.D(n364), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][6]  (.RN(n452), 
	.Q(\reg_array[1][6] ), 
	.D(n365), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][5]  (.RN(n452), 
	.Q(\reg_array[1][5] ), 
	.D(n366), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][4]  (.RN(n452), 
	.Q(\reg_array[1][4] ), 
	.D(n367), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][3]  (.RN(n452), 
	.Q(\reg_array[1][3] ), 
	.D(n368), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][2]  (.RN(n452), 
	.Q(\reg_array[1][2] ), 
	.D(n369), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][1]  (.RN(n452), 
	.Q(\reg_array[1][1] ), 
	.D(n370), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[1][0]  (.RN(n452), 
	.Q(\reg_array[1][0] ), 
	.D(n371), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][15]  (.RN(n452), 
	.Q(\reg_array[7][15] ), 
	.D(n372), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][14]  (.RN(n452), 
	.Q(\reg_array[7][14] ), 
	.D(n373), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][13]  (.RN(n452), 
	.Q(\reg_array[7][13] ), 
	.D(n374), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][12]  (.RN(n452), 
	.Q(\reg_array[7][12] ), 
	.D(n375), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][11]  (.RN(n452), 
	.Q(\reg_array[7][11] ), 
	.D(n376), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][10]  (.RN(n452), 
	.Q(\reg_array[7][10] ), 
	.D(n377), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][9]  (.RN(n452), 
	.Q(\reg_array[7][9] ), 
	.D(n378), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][8]  (.RN(n452), 
	.Q(\reg_array[7][8] ), 
	.D(n379), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][7]  (.RN(n452), 
	.Q(\reg_array[7][7] ), 
	.D(n380), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][6]  (.RN(n452), 
	.Q(\reg_array[7][6] ), 
	.D(n381), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][5]  (.RN(n452), 
	.Q(\reg_array[7][5] ), 
	.D(n382), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][4]  (.RN(n452), 
	.Q(\reg_array[7][4] ), 
	.D(n383), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][3]  (.RN(n452), 
	.Q(\reg_array[7][3] ), 
	.D(n384), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][2]  (.RN(n452), 
	.Q(\reg_array[7][2] ), 
	.D(n385), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][1]  (.RN(n452), 
	.Q(\reg_array[7][1] ), 
	.D(n386), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[7][0]  (.RN(n452), 
	.Q(\reg_array[7][0] ), 
	.D(n387), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][15]  (.RN(n452), 
	.Q(\reg_array[3][15] ), 
	.D(n388), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][14]  (.RN(n452), 
	.Q(\reg_array[3][14] ), 
	.D(n389), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][13]  (.RN(n452), 
	.Q(\reg_array[3][13] ), 
	.D(n390), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][12]  (.RN(n452), 
	.Q(\reg_array[3][12] ), 
	.D(n391), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][11]  (.RN(n452), 
	.Q(\reg_array[3][11] ), 
	.D(n392), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][10]  (.RN(n452), 
	.Q(\reg_array[3][10] ), 
	.D(n393), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][9]  (.RN(n452), 
	.Q(\reg_array[3][9] ), 
	.D(n394), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][8]  (.RN(n452), 
	.Q(\reg_array[3][8] ), 
	.D(n395), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][7]  (.RN(n452), 
	.Q(\reg_array[3][7] ), 
	.D(n396), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][6]  (.RN(n452), 
	.Q(\reg_array[3][6] ), 
	.D(n397), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][5]  (.RN(n452), 
	.Q(\reg_array[3][5] ), 
	.D(n398), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][4]  (.RN(n452), 
	.Q(\reg_array[3][4] ), 
	.D(n399), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][3]  (.RN(n452), 
	.Q(\reg_array[3][3] ), 
	.D(n400), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][2]  (.RN(n452), 
	.Q(\reg_array[3][2] ), 
	.D(n401), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][1]  (.RN(n452), 
	.Q(\reg_array[3][1] ), 
	.D(n402), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[3][0]  (.RN(n452), 
	.Q(\reg_array[3][0] ), 
	.D(n403), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][15]  (.RN(n452), 
	.Q(\reg_array[2][15] ), 
	.D(n436), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][14]  (.RN(n452), 
	.Q(\reg_array[2][14] ), 
	.D(n437), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][13]  (.RN(n452), 
	.Q(\reg_array[2][13] ), 
	.D(n438), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][12]  (.RN(n452), 
	.Q(\reg_array[2][12] ), 
	.D(n439), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][11]  (.RN(n452), 
	.Q(\reg_array[2][11] ), 
	.D(n440), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][10]  (.RN(n452), 
	.Q(\reg_array[2][10] ), 
	.D(n441), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][9]  (.RN(n452), 
	.Q(\reg_array[2][9] ), 
	.D(n442), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][8]  (.RN(n452), 
	.Q(\reg_array[2][8] ), 
	.D(n443), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][7]  (.RN(n452), 
	.Q(\reg_array[2][7] ), 
	.D(n444), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][6]  (.RN(n452), 
	.Q(\reg_array[2][6] ), 
	.D(n445), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][5]  (.RN(n452), 
	.Q(\reg_array[2][5] ), 
	.D(n446), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][4]  (.RN(n452), 
	.Q(\reg_array[2][4] ), 
	.D(n447), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][3]  (.RN(n452), 
	.Q(\reg_array[2][3] ), 
	.D(n448), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][2]  (.RN(n452), 
	.Q(\reg_array[2][2] ), 
	.D(n449), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][1]  (.RN(n452), 
	.Q(\reg_array[2][1] ), 
	.D(n450), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[2][0]  (.RN(n452), 
	.Q(\reg_array[2][0] ), 
	.D(n451), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][15]  (.RN(n452), 
	.Q(\reg_array[6][15] ), 
	.D(n420), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][14]  (.RN(n452), 
	.Q(\reg_array[6][14] ), 
	.D(n421), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][13]  (.RN(n452), 
	.Q(\reg_array[6][13] ), 
	.D(n422), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][12]  (.RN(n452), 
	.Q(\reg_array[6][12] ), 
	.D(n423), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][11]  (.RN(n452), 
	.Q(\reg_array[6][11] ), 
	.D(n424), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][10]  (.RN(n452), 
	.Q(\reg_array[6][10] ), 
	.D(n425), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][9]  (.RN(n452), 
	.Q(\reg_array[6][9] ), 
	.D(n426), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][8]  (.RN(n452), 
	.Q(\reg_array[6][8] ), 
	.D(n427), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][7]  (.RN(n452), 
	.Q(\reg_array[6][7] ), 
	.D(n428), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][6]  (.RN(n452), 
	.Q(\reg_array[6][6] ), 
	.D(n429), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][5]  (.RN(n452), 
	.Q(\reg_array[6][5] ), 
	.D(n430), 
	.CK(clk));
   DFFRHQXL \reg_array_reg[6][4]  (.RN(n452), 
	.Q(\reg_array[6][4] ), 
	.D(n431), 
	.CK(clk));
   DFFRHQX1 \reg_array_reg[6][3]  (.RN(n452), 
	.Q(\reg_array[6][3] ), 
	.D(n432), 
	.CK(clk));
   DFFRHQX1 \reg_array_reg[6][2]  (.RN(n452), 
	.Q(\reg_array[6][2] ), 
	.D(n433), 
	.CK(clk));
   DFFRHQX1 \reg_array_reg[6][1]  (.RN(n452), 
	.Q(\reg_array[6][1] ), 
	.D(n434), 
	.CK(clk));
   DFFRHQX1 \reg_array_reg[6][0]  (.RN(n452), 
	.Q(\reg_array[6][0] ), 
	.D(n435), 
	.CK(clk));
   NAND3X1 U2 (.Y(reg_read_data_2[9]), 
	.C(n211), 
	.B(n210), 
	.A(n209));
   AOI222X1 U3 (.Y(n211), 
	.C1(n214), 
	.C0(\reg_array[3][9] ), 
	.B1(n213), 
	.B0(\reg_array[2][9] ), 
	.A1(n212), 
	.A0(\reg_array[6][9] ));
   AOI22X1 U4 (.Y(n210), 
	.B1(n216), 
	.B0(\reg_array[5][9] ), 
	.A1(n215), 
	.A0(\reg_array[7][9] ));
   AOI22X1 U5 (.Y(n209), 
	.B1(n218), 
	.B0(\reg_array[4][9] ), 
	.A1(n217), 
	.A0(\reg_array[1][9] ));
   NAND3X1 U6 (.Y(reg_read_data_2[8]), 
	.C(n221), 
	.B(n220), 
	.A(n219));
   AOI222X1 U7 (.Y(n221), 
	.C1(n214), 
	.C0(\reg_array[3][8] ), 
	.B1(n213), 
	.B0(\reg_array[2][8] ), 
	.A1(n212), 
	.A0(\reg_array[6][8] ));
   AOI22X1 U8 (.Y(n220), 
	.B1(n216), 
	.B0(\reg_array[5][8] ), 
	.A1(n215), 
	.A0(\reg_array[7][8] ));
   AOI22X1 U9 (.Y(n219), 
	.B1(n218), 
	.B0(\reg_array[4][8] ), 
	.A1(n217), 
	.A0(\reg_array[1][8] ));
   NAND3X1 U10 (.Y(reg_read_data_2[7]), 
	.C(n224), 
	.B(n223), 
	.A(n222));
   AOI222X1 U11 (.Y(n224), 
	.C1(n214), 
	.C0(\reg_array[3][7] ), 
	.B1(n213), 
	.B0(\reg_array[2][7] ), 
	.A1(n212), 
	.A0(\reg_array[6][7] ));
   AOI22X1 U12 (.Y(n223), 
	.B1(n216), 
	.B0(\reg_array[5][7] ), 
	.A1(n215), 
	.A0(\reg_array[7][7] ));
   AOI22X1 U13 (.Y(n222), 
	.B1(n218), 
	.B0(\reg_array[4][7] ), 
	.A1(n217), 
	.A0(\reg_array[1][7] ));
   NAND3X1 U14 (.Y(reg_read_data_2[6]), 
	.C(n227), 
	.B(n226), 
	.A(n225));
   AOI222X1 U15 (.Y(n227), 
	.C1(n214), 
	.C0(\reg_array[3][6] ), 
	.B1(n213), 
	.B0(\reg_array[2][6] ), 
	.A1(n212), 
	.A0(\reg_array[6][6] ));
   AOI22X1 U16 (.Y(n226), 
	.B1(n216), 
	.B0(\reg_array[5][6] ), 
	.A1(n215), 
	.A0(\reg_array[7][6] ));
   AOI22X1 U17 (.Y(n225), 
	.B1(n218), 
	.B0(\reg_array[4][6] ), 
	.A1(n217), 
	.A0(\reg_array[1][6] ));
   NAND3X1 U18 (.Y(reg_read_data_2[5]), 
	.C(n230), 
	.B(n229), 
	.A(n228));
   AOI222X1 U19 (.Y(n230), 
	.C1(n214), 
	.C0(\reg_array[3][5] ), 
	.B1(n213), 
	.B0(\reg_array[2][5] ), 
	.A1(n212), 
	.A0(\reg_array[6][5] ));
   AOI22X1 U20 (.Y(n229), 
	.B1(n216), 
	.B0(\reg_array[5][5] ), 
	.A1(n215), 
	.A0(\reg_array[7][5] ));
   AOI22X1 U21 (.Y(n228), 
	.B1(n218), 
	.B0(\reg_array[4][5] ), 
	.A1(n217), 
	.A0(\reg_array[1][5] ));
   NAND3X1 U22 (.Y(reg_read_data_2[4]), 
	.C(n233), 
	.B(n232), 
	.A(n231));
   AOI222X1 U23 (.Y(n233), 
	.C1(n214), 
	.C0(\reg_array[3][4] ), 
	.B1(n213), 
	.B0(\reg_array[2][4] ), 
	.A1(n212), 
	.A0(\reg_array[6][4] ));
   AOI22X1 U24 (.Y(n232), 
	.B1(n216), 
	.B0(\reg_array[5][4] ), 
	.A1(n215), 
	.A0(\reg_array[7][4] ));
   AOI22X1 U25 (.Y(n231), 
	.B1(n218), 
	.B0(\reg_array[4][4] ), 
	.A1(n217), 
	.A0(\reg_array[1][4] ));
   NAND3X1 U26 (.Y(reg_read_data_2[3]), 
	.C(n236), 
	.B(n235), 
	.A(n234));
   AOI222X1 U27 (.Y(n236), 
	.C1(n214), 
	.C0(\reg_array[3][3] ), 
	.B1(n213), 
	.B0(\reg_array[2][3] ), 
	.A1(n212), 
	.A0(\reg_array[6][3] ));
   AOI22X1 U28 (.Y(n235), 
	.B1(n216), 
	.B0(\reg_array[5][3] ), 
	.A1(n215), 
	.A0(\reg_array[7][3] ));
   AOI22X1 U29 (.Y(n234), 
	.B1(n218), 
	.B0(\reg_array[4][3] ), 
	.A1(n217), 
	.A0(\reg_array[1][3] ));
   NAND3X1 U30 (.Y(reg_read_data_2[2]), 
	.C(n239), 
	.B(n238), 
	.A(n237));
   AOI222X1 U31 (.Y(n239), 
	.C1(n214), 
	.C0(\reg_array[3][2] ), 
	.B1(n213), 
	.B0(\reg_array[2][2] ), 
	.A1(n212), 
	.A0(\reg_array[6][2] ));
   AOI22X1 U32 (.Y(n238), 
	.B1(n216), 
	.B0(\reg_array[5][2] ), 
	.A1(n215), 
	.A0(\reg_array[7][2] ));
   AOI22X1 U33 (.Y(n237), 
	.B1(n218), 
	.B0(\reg_array[4][2] ), 
	.A1(n217), 
	.A0(\reg_array[1][2] ));
   NAND3X1 U34 (.Y(reg_read_data_2[1]), 
	.C(n242), 
	.B(n241), 
	.A(n240));
   AOI222X1 U35 (.Y(n242), 
	.C1(n214), 
	.C0(\reg_array[3][1] ), 
	.B1(n213), 
	.B0(\reg_array[2][1] ), 
	.A1(n212), 
	.A0(\reg_array[6][1] ));
   AOI22X1 U36 (.Y(n241), 
	.B1(n216), 
	.B0(\reg_array[5][1] ), 
	.A1(n215), 
	.A0(\reg_array[7][1] ));
   AOI22X1 U37 (.Y(n240), 
	.B1(n218), 
	.B0(\reg_array[4][1] ), 
	.A1(n217), 
	.A0(\reg_array[1][1] ));
   NAND3X1 U38 (.Y(reg_read_data_2[15]), 
	.C(n245), 
	.B(n244), 
	.A(n243));
   AOI222X1 U39 (.Y(n245), 
	.C1(n214), 
	.C0(\reg_array[3][15] ), 
	.B1(n213), 
	.B0(\reg_array[2][15] ), 
	.A1(n212), 
	.A0(\reg_array[6][15] ));
   AOI22X1 U40 (.Y(n244), 
	.B1(n216), 
	.B0(\reg_array[5][15] ), 
	.A1(n215), 
	.A0(\reg_array[7][15] ));
   AOI22X1 U41 (.Y(n243), 
	.B1(n218), 
	.B0(\reg_array[4][15] ), 
	.A1(n217), 
	.A0(\reg_array[1][15] ));
   NAND3X1 U42 (.Y(reg_read_data_2[14]), 
	.C(n248), 
	.B(n247), 
	.A(n246));
   AOI222X1 U43 (.Y(n248), 
	.C1(n214), 
	.C0(\reg_array[3][14] ), 
	.B1(n213), 
	.B0(\reg_array[2][14] ), 
	.A1(n212), 
	.A0(\reg_array[6][14] ));
   AOI22X1 U44 (.Y(n247), 
	.B1(n216), 
	.B0(\reg_array[5][14] ), 
	.A1(n215), 
	.A0(\reg_array[7][14] ));
   AOI22X1 U45 (.Y(n246), 
	.B1(n218), 
	.B0(\reg_array[4][14] ), 
	.A1(n217), 
	.A0(\reg_array[1][14] ));
   NAND3X1 U46 (.Y(reg_read_data_2[13]), 
	.C(n251), 
	.B(n250), 
	.A(n249));
   AOI222X1 U47 (.Y(n251), 
	.C1(n214), 
	.C0(\reg_array[3][13] ), 
	.B1(n213), 
	.B0(\reg_array[2][13] ), 
	.A1(n212), 
	.A0(\reg_array[6][13] ));
   AOI22X1 U48 (.Y(n250), 
	.B1(n216), 
	.B0(\reg_array[5][13] ), 
	.A1(n215), 
	.A0(\reg_array[7][13] ));
   AOI22X1 U49 (.Y(n249), 
	.B1(n218), 
	.B0(\reg_array[4][13] ), 
	.A1(n217), 
	.A0(\reg_array[1][13] ));
   NAND3X1 U50 (.Y(reg_read_data_2[12]), 
	.C(n254), 
	.B(n253), 
	.A(n252));
   AOI222X1 U51 (.Y(n254), 
	.C1(n214), 
	.C0(\reg_array[3][12] ), 
	.B1(n213), 
	.B0(\reg_array[2][12] ), 
	.A1(n212), 
	.A0(\reg_array[6][12] ));
   AOI22X1 U52 (.Y(n253), 
	.B1(n216), 
	.B0(\reg_array[5][12] ), 
	.A1(n215), 
	.A0(\reg_array[7][12] ));
   AOI22X1 U53 (.Y(n252), 
	.B1(n218), 
	.B0(\reg_array[4][12] ), 
	.A1(n217), 
	.A0(\reg_array[1][12] ));
   NAND3X1 U54 (.Y(reg_read_data_2[11]), 
	.C(n257), 
	.B(n256), 
	.A(n255));
   AOI222X1 U55 (.Y(n257), 
	.C1(n214), 
	.C0(\reg_array[3][11] ), 
	.B1(n213), 
	.B0(\reg_array[2][11] ), 
	.A1(n212), 
	.A0(\reg_array[6][11] ));
   AOI22X1 U56 (.Y(n256), 
	.B1(n216), 
	.B0(\reg_array[5][11] ), 
	.A1(n215), 
	.A0(\reg_array[7][11] ));
   AOI22X1 U57 (.Y(n255), 
	.B1(n218), 
	.B0(\reg_array[4][11] ), 
	.A1(n217), 
	.A0(\reg_array[1][11] ));
   NAND3X1 U58 (.Y(reg_read_data_2[10]), 
	.C(n260), 
	.B(n259), 
	.A(n258));
   AOI222X1 U59 (.Y(n260), 
	.C1(n214), 
	.C0(\reg_array[3][10] ), 
	.B1(n213), 
	.B0(\reg_array[2][10] ), 
	.A1(n212), 
	.A0(\reg_array[6][10] ));
   AOI22X1 U60 (.Y(n259), 
	.B1(n216), 
	.B0(\reg_array[5][10] ), 
	.A1(n215), 
	.A0(\reg_array[7][10] ));
   AOI22X1 U61 (.Y(n258), 
	.B1(n218), 
	.B0(\reg_array[4][10] ), 
	.A1(n217), 
	.A0(\reg_array[1][10] ));
   NAND3X1 U62 (.Y(reg_read_data_2[0]), 
	.C(n263), 
	.B(n262), 
	.A(n261));
   AOI222X1 U63 (.Y(n263), 
	.C1(n214), 
	.C0(\reg_array[3][0] ), 
	.B1(n213), 
	.B0(\reg_array[2][0] ), 
	.A1(n212), 
	.A0(\reg_array[6][0] ));
   NOR3X1 U64 (.Y(n214), 
	.C(n265), 
	.B(N23), 
	.A(n264));
   NOR3X1 U65 (.Y(n213), 
	.C(n264), 
	.B(N23), 
	.A(N21));
   NOR3X1 U66 (.Y(n212), 
	.C(n266), 
	.B(N21), 
	.A(n264));
   AOI22X1 U67 (.Y(n262), 
	.B1(n216), 
	.B0(\reg_array[5][0] ), 
	.A1(n215), 
	.A0(\reg_array[7][0] ));
   NOR3X1 U68 (.Y(n216), 
	.C(n266), 
	.B(N22), 
	.A(n265));
   NOR3X1 U69 (.Y(n215), 
	.C(n266), 
	.B(n264), 
	.A(n265));
   INVX1 U70 (.Y(n266), 
	.A(N23));
   AOI22X1 U71 (.Y(n261), 
	.B1(n218), 
	.B0(\reg_array[4][0] ), 
	.A1(n217), 
	.A0(\reg_array[1][0] ));
   AND3X1 U72 (.Y(n218), 
	.C(n267), 
	.B(n264), 
	.A(n265));
   INVX1 U73 (.Y(n264), 
	.A(N22));
   AND2X1 U74 (.Y(n217), 
	.B(n267), 
	.A(n268));
   NAND2X1 U75 (.Y(n267), 
	.B(n265), 
	.A(n268));
   INVX1 U76 (.Y(n265), 
	.A(N21));
   NOR2X1 U77 (.Y(n268), 
	.B(N23), 
	.A(N22));
   NAND3X1 U78 (.Y(reg_read_data_1[9]), 
	.C(n271), 
	.B(n270), 
	.A(n269));
   AOI222X1 U79 (.Y(n271), 
	.C1(\reg_array[3][9] ), 
	.C0(n274), 
	.B1(\reg_array[2][9] ), 
	.B0(n273), 
	.A1(\reg_array[6][9] ), 
	.A0(n272));
   AOI22X1 U80 (.Y(n270), 
	.B1(\reg_array[5][9] ), 
	.B0(n276), 
	.A1(\reg_array[7][9] ), 
	.A0(n275));
   AOI22X1 U81 (.Y(n269), 
	.B1(\reg_array[4][9] ), 
	.B0(n278), 
	.A1(\reg_array[1][9] ), 
	.A0(n277));
   NAND3X1 U82 (.Y(reg_read_data_1[8]), 
	.C(n281), 
	.B(n280), 
	.A(n279));
   AOI222X1 U83 (.Y(n281), 
	.C1(\reg_array[3][8] ), 
	.C0(n274), 
	.B1(\reg_array[2][8] ), 
	.B0(n273), 
	.A1(\reg_array[6][8] ), 
	.A0(n272));
   AOI22X1 U84 (.Y(n280), 
	.B1(\reg_array[5][8] ), 
	.B0(n276), 
	.A1(\reg_array[7][8] ), 
	.A0(n275));
   AOI22X1 U85 (.Y(n279), 
	.B1(\reg_array[4][8] ), 
	.B0(n278), 
	.A1(\reg_array[1][8] ), 
	.A0(n277));
   NAND3X1 U86 (.Y(reg_read_data_1[7]), 
	.C(n284), 
	.B(n283), 
	.A(n282));
   AOI222X1 U87 (.Y(n284), 
	.C1(\reg_array[3][7] ), 
	.C0(n274), 
	.B1(\reg_array[2][7] ), 
	.B0(n273), 
	.A1(\reg_array[6][7] ), 
	.A0(n272));
   AOI22X1 U88 (.Y(n283), 
	.B1(\reg_array[5][7] ), 
	.B0(n276), 
	.A1(\reg_array[7][7] ), 
	.A0(n275));
   AOI22X1 U89 (.Y(n282), 
	.B1(\reg_array[4][7] ), 
	.B0(n278), 
	.A1(\reg_array[1][7] ), 
	.A0(n277));
   NAND3X1 U90 (.Y(reg_read_data_1[6]), 
	.C(n287), 
	.B(n286), 
	.A(n285));
   AOI222X1 U91 (.Y(n287), 
	.C1(\reg_array[3][6] ), 
	.C0(n274), 
	.B1(\reg_array[2][6] ), 
	.B0(n273), 
	.A1(\reg_array[6][6] ), 
	.A0(n272));
   AOI22X1 U92 (.Y(n286), 
	.B1(\reg_array[5][6] ), 
	.B0(n276), 
	.A1(\reg_array[7][6] ), 
	.A0(n275));
   AOI22X1 U93 (.Y(n285), 
	.B1(\reg_array[4][6] ), 
	.B0(n278), 
	.A1(\reg_array[1][6] ), 
	.A0(n277));
   NAND3X1 U94 (.Y(reg_read_data_1[5]), 
	.C(n290), 
	.B(n289), 
	.A(n288));
   AOI222X1 U95 (.Y(n290), 
	.C1(\reg_array[3][5] ), 
	.C0(n274), 
	.B1(\reg_array[2][5] ), 
	.B0(n273), 
	.A1(\reg_array[6][5] ), 
	.A0(n272));
   AOI22X1 U96 (.Y(n289), 
	.B1(\reg_array[5][5] ), 
	.B0(n276), 
	.A1(\reg_array[7][5] ), 
	.A0(n275));
   AOI22X1 U97 (.Y(n288), 
	.B1(\reg_array[4][5] ), 
	.B0(n278), 
	.A1(\reg_array[1][5] ), 
	.A0(n277));
   NAND3X1 U98 (.Y(reg_read_data_1[4]), 
	.C(n293), 
	.B(n292), 
	.A(n291));
   AOI222X1 U99 (.Y(n293), 
	.C1(\reg_array[3][4] ), 
	.C0(n274), 
	.B1(\reg_array[2][4] ), 
	.B0(n273), 
	.A1(\reg_array[6][4] ), 
	.A0(n272));
   AOI22X1 U100 (.Y(n292), 
	.B1(\reg_array[5][4] ), 
	.B0(n276), 
	.A1(\reg_array[7][4] ), 
	.A0(n275));
   AOI22X1 U101 (.Y(n291), 
	.B1(\reg_array[4][4] ), 
	.B0(n278), 
	.A1(\reg_array[1][4] ), 
	.A0(n277));
   NAND3X1 U102 (.Y(reg_read_data_1[3]), 
	.C(n296), 
	.B(n295), 
	.A(n294));
   AOI222X1 U103 (.Y(n296), 
	.C1(\reg_array[3][3] ), 
	.C0(n274), 
	.B1(\reg_array[2][3] ), 
	.B0(n273), 
	.A1(\reg_array[6][3] ), 
	.A0(n272));
   AOI22X1 U104 (.Y(n295), 
	.B1(\reg_array[5][3] ), 
	.B0(n276), 
	.A1(\reg_array[7][3] ), 
	.A0(n275));
   AOI22X1 U105 (.Y(n294), 
	.B1(\reg_array[4][3] ), 
	.B0(n278), 
	.A1(\reg_array[1][3] ), 
	.A0(n277));
   NAND3X1 U106 (.Y(reg_read_data_1[2]), 
	.C(n299), 
	.B(n298), 
	.A(n297));
   AOI222X1 U107 (.Y(n299), 
	.C1(\reg_array[3][2] ), 
	.C0(n274), 
	.B1(\reg_array[2][2] ), 
	.B0(n273), 
	.A1(\reg_array[6][2] ), 
	.A0(n272));
   AOI22X1 U108 (.Y(n298), 
	.B1(\reg_array[5][2] ), 
	.B0(n276), 
	.A1(\reg_array[7][2] ), 
	.A0(n275));
   AOI22X1 U109 (.Y(n297), 
	.B1(\reg_array[4][2] ), 
	.B0(n278), 
	.A1(\reg_array[1][2] ), 
	.A0(n277));
   NAND3X1 U110 (.Y(reg_read_data_1[1]), 
	.C(n302), 
	.B(n301), 
	.A(n300));
   AOI222X1 U111 (.Y(n302), 
	.C1(\reg_array[3][1] ), 
	.C0(n274), 
	.B1(\reg_array[2][1] ), 
	.B0(n273), 
	.A1(\reg_array[6][1] ), 
	.A0(n272));
   AOI22X1 U112 (.Y(n301), 
	.B1(\reg_array[5][1] ), 
	.B0(n276), 
	.A1(\reg_array[7][1] ), 
	.A0(n275));
   AOI22X1 U113 (.Y(n300), 
	.B1(\reg_array[4][1] ), 
	.B0(n278), 
	.A1(\reg_array[1][1] ), 
	.A0(n277));
   NAND3X1 U114 (.Y(reg_read_data_1[15]), 
	.C(n305), 
	.B(n304), 
	.A(n303));
   AOI222X1 U115 (.Y(n305), 
	.C1(\reg_array[3][15] ), 
	.C0(n274), 
	.B1(\reg_array[2][15] ), 
	.B0(n273), 
	.A1(\reg_array[6][15] ), 
	.A0(n272));
   AOI22X1 U116 (.Y(n304), 
	.B1(\reg_array[5][15] ), 
	.B0(n276), 
	.A1(\reg_array[7][15] ), 
	.A0(n275));
   AOI22X1 U117 (.Y(n303), 
	.B1(\reg_array[4][15] ), 
	.B0(n278), 
	.A1(\reg_array[1][15] ), 
	.A0(n277));
   NAND3X1 U118 (.Y(reg_read_data_1[14]), 
	.C(n308), 
	.B(n307), 
	.A(n306));
   AOI222X1 U119 (.Y(n308), 
	.C1(\reg_array[3][14] ), 
	.C0(n274), 
	.B1(\reg_array[2][14] ), 
	.B0(n273), 
	.A1(\reg_array[6][14] ), 
	.A0(n272));
   AOI22X1 U120 (.Y(n307), 
	.B1(\reg_array[5][14] ), 
	.B0(n276), 
	.A1(\reg_array[7][14] ), 
	.A0(n275));
   AOI22X1 U121 (.Y(n306), 
	.B1(\reg_array[4][14] ), 
	.B0(n278), 
	.A1(\reg_array[1][14] ), 
	.A0(n277));
   NAND3X1 U122 (.Y(reg_read_data_1[13]), 
	.C(n311), 
	.B(n310), 
	.A(n309));
   AOI222X1 U123 (.Y(n311), 
	.C1(\reg_array[3][13] ), 
	.C0(n274), 
	.B1(\reg_array[2][13] ), 
	.B0(n273), 
	.A1(\reg_array[6][13] ), 
	.A0(n272));
   AOI22X1 U124 (.Y(n310), 
	.B1(\reg_array[5][13] ), 
	.B0(n276), 
	.A1(\reg_array[7][13] ), 
	.A0(n275));
   AOI22X1 U125 (.Y(n309), 
	.B1(\reg_array[4][13] ), 
	.B0(n278), 
	.A1(\reg_array[1][13] ), 
	.A0(n277));
   NAND3X1 U126 (.Y(reg_read_data_1[12]), 
	.C(n314), 
	.B(n313), 
	.A(n312));
   AOI222X1 U127 (.Y(n314), 
	.C1(\reg_array[3][12] ), 
	.C0(n274), 
	.B1(\reg_array[2][12] ), 
	.B0(n273), 
	.A1(\reg_array[6][12] ), 
	.A0(n272));
   AOI22X1 U128 (.Y(n313), 
	.B1(\reg_array[5][12] ), 
	.B0(n276), 
	.A1(\reg_array[7][12] ), 
	.A0(n275));
   AOI22X1 U129 (.Y(n312), 
	.B1(\reg_array[4][12] ), 
	.B0(n278), 
	.A1(\reg_array[1][12] ), 
	.A0(n277));
   NAND3X1 U130 (.Y(reg_read_data_1[11]), 
	.C(n317), 
	.B(n316), 
	.A(n315));
   AOI222X1 U131 (.Y(n317), 
	.C1(\reg_array[3][11] ), 
	.C0(n274), 
	.B1(\reg_array[2][11] ), 
	.B0(n273), 
	.A1(\reg_array[6][11] ), 
	.A0(n272));
   AOI22X1 U132 (.Y(n316), 
	.B1(\reg_array[5][11] ), 
	.B0(n276), 
	.A1(\reg_array[7][11] ), 
	.A0(n275));
   AOI22X1 U133 (.Y(n315), 
	.B1(\reg_array[4][11] ), 
	.B0(n278), 
	.A1(\reg_array[1][11] ), 
	.A0(n277));
   NAND3X1 U134 (.Y(reg_read_data_1[10]), 
	.C(n320), 
	.B(n319), 
	.A(n318));
   AOI222X1 U135 (.Y(n320), 
	.C1(\reg_array[3][10] ), 
	.C0(n274), 
	.B1(\reg_array[2][10] ), 
	.B0(n273), 
	.A1(\reg_array[6][10] ), 
	.A0(n272));
   AOI22X1 U136 (.Y(n319), 
	.B1(\reg_array[5][10] ), 
	.B0(n276), 
	.A1(\reg_array[7][10] ), 
	.A0(n275));
   AOI22X1 U137 (.Y(n318), 
	.B1(\reg_array[4][10] ), 
	.B0(n278), 
	.A1(\reg_array[1][10] ), 
	.A0(n277));
   NAND3X1 U138 (.Y(reg_read_data_1[0]), 
	.C(n323), 
	.B(n322), 
	.A(n321));
   AOI222X1 U139 (.Y(n323), 
	.C1(\reg_array[3][0] ), 
	.C0(n274), 
	.B1(\reg_array[2][0] ), 
	.B0(n273), 
	.A1(\reg_array[6][0] ), 
	.A0(n272));
   NOR3X1 U140 (.Y(n274), 
	.C(n325), 
	.B(N20), 
	.A(n324));
   NOR3X1 U141 (.Y(n273), 
	.C(n324), 
	.B(N20), 
	.A(N18));
   NOR3X1 U142 (.Y(n272), 
	.C(n326), 
	.B(N18), 
	.A(n324));
   AOI22X1 U143 (.Y(n322), 
	.B1(\reg_array[5][0] ), 
	.B0(n276), 
	.A1(\reg_array[7][0] ), 
	.A0(n275));
   NOR3X1 U144 (.Y(n276), 
	.C(n326), 
	.B(N19), 
	.A(n325));
   NOR3X1 U145 (.Y(n275), 
	.C(n326), 
	.B(n324), 
	.A(n325));
   INVX1 U146 (.Y(n326), 
	.A(N20));
   AOI22X1 U147 (.Y(n321), 
	.B1(\reg_array[4][0] ), 
	.B0(n278), 
	.A1(\reg_array[1][0] ), 
	.A0(n277));
   AND3X1 U148 (.Y(n278), 
	.C(n327), 
	.B(n324), 
	.A(n325));
   INVX1 U149 (.Y(n324), 
	.A(N19));
   AND2X1 U150 (.Y(n277), 
	.B(n327), 
	.A(n328));
   NAND2X1 U151 (.Y(n327), 
	.B(n325), 
	.A(n328));
   INVX1 U152 (.Y(n325), 
	.A(N18));
   NOR2X1 U153 (.Y(n328), 
	.B(N20), 
	.A(N19));
   MX2X1 U154 (.Y(n340), 
	.S0(n329), 
	.B(reg_write_data[15]), 
	.A(\reg_array[5][15] ));
   MX2X1 U155 (.Y(n341), 
	.S0(n329), 
	.B(reg_write_data[14]), 
	.A(\reg_array[5][14] ));
   MX2X1 U156 (.Y(n342), 
	.S0(n329), 
	.B(reg_write_data[13]), 
	.A(\reg_array[5][13] ));
   MX2X1 U157 (.Y(n343), 
	.S0(n329), 
	.B(reg_write_data[12]), 
	.A(\reg_array[5][12] ));
   MX2X1 U158 (.Y(n344), 
	.S0(n329), 
	.B(reg_write_data[11]), 
	.A(\reg_array[5][11] ));
   MX2X1 U159 (.Y(n345), 
	.S0(n329), 
	.B(reg_write_data[10]), 
	.A(\reg_array[5][10] ));
   MX2X1 U160 (.Y(n346), 
	.S0(n329), 
	.B(reg_write_data[9]), 
	.A(\reg_array[5][9] ));
   MX2X1 U161 (.Y(n347), 
	.S0(n329), 
	.B(reg_write_data[8]), 
	.A(\reg_array[5][8] ));
   MX2X1 U162 (.Y(n348), 
	.S0(n329), 
	.B(reg_write_data[7]), 
	.A(\reg_array[5][7] ));
   MX2X1 U163 (.Y(n349), 
	.S0(n329), 
	.B(reg_write_data[6]), 
	.A(\reg_array[5][6] ));
   MX2X1 U164 (.Y(n350), 
	.S0(n329), 
	.B(reg_write_data[5]), 
	.A(\reg_array[5][5] ));
   MX2X1 U165 (.Y(n351), 
	.S0(n329), 
	.B(reg_write_data[4]), 
	.A(\reg_array[5][4] ));
   MX2X1 U166 (.Y(n352), 
	.S0(n329), 
	.B(reg_write_data[3]), 
	.A(\reg_array[5][3] ));
   MX2X1 U167 (.Y(n353), 
	.S0(n329), 
	.B(reg_write_data[2]), 
	.A(\reg_array[5][2] ));
   MX2X1 U168 (.Y(n354), 
	.S0(n329), 
	.B(reg_write_data[1]), 
	.A(\reg_array[5][1] ));
   MX2X1 U169 (.Y(n355), 
	.S0(n329), 
	.B(reg_write_data[0]), 
	.A(\reg_array[5][0] ));
   AND3X1 U170 (.Y(n329), 
	.C(reg_write_dest[2]), 
	.B(n330), 
	.A(reg_write_dest[0]));
   MX2X1 U171 (.Y(n356), 
	.S0(n331), 
	.B(reg_write_data[15]), 
	.A(\reg_array[1][15] ));
   MX2X1 U172 (.Y(n357), 
	.S0(n331), 
	.B(reg_write_data[14]), 
	.A(\reg_array[1][14] ));
   MX2X1 U173 (.Y(n358), 
	.S0(n331), 
	.B(reg_write_data[13]), 
	.A(\reg_array[1][13] ));
   MX2X1 U174 (.Y(n359), 
	.S0(n331), 
	.B(reg_write_data[12]), 
	.A(\reg_array[1][12] ));
   MX2X1 U175 (.Y(n360), 
	.S0(n331), 
	.B(reg_write_data[11]), 
	.A(\reg_array[1][11] ));
   MX2X1 U176 (.Y(n361), 
	.S0(n331), 
	.B(reg_write_data[10]), 
	.A(\reg_array[1][10] ));
   MX2X1 U177 (.Y(n362), 
	.S0(n331), 
	.B(reg_write_data[9]), 
	.A(\reg_array[1][9] ));
   MX2X1 U178 (.Y(n363), 
	.S0(n331), 
	.B(reg_write_data[8]), 
	.A(\reg_array[1][8] ));
   MX2X1 U179 (.Y(n364), 
	.S0(n331), 
	.B(reg_write_data[7]), 
	.A(\reg_array[1][7] ));
   MX2X1 U180 (.Y(n365), 
	.S0(n331), 
	.B(reg_write_data[6]), 
	.A(\reg_array[1][6] ));
   MX2X1 U181 (.Y(n366), 
	.S0(n331), 
	.B(reg_write_data[5]), 
	.A(\reg_array[1][5] ));
   MX2X1 U182 (.Y(n367), 
	.S0(n331), 
	.B(reg_write_data[4]), 
	.A(\reg_array[1][4] ));
   MX2X1 U183 (.Y(n368), 
	.S0(n331), 
	.B(reg_write_data[3]), 
	.A(\reg_array[1][3] ));
   MX2X1 U184 (.Y(n369), 
	.S0(n331), 
	.B(reg_write_data[2]), 
	.A(\reg_array[1][2] ));
   MX2X1 U185 (.Y(n370), 
	.S0(n331), 
	.B(reg_write_data[1]), 
	.A(\reg_array[1][1] ));
   MX2X1 U186 (.Y(n371), 
	.S0(n331), 
	.B(reg_write_data[0]), 
	.A(\reg_array[1][0] ));
   AND3X1 U187 (.Y(n331), 
	.C(reg_write_dest[0]), 
	.B(n332), 
	.A(n330));
   MX2X1 U188 (.Y(n372), 
	.S0(n333), 
	.B(reg_write_data[15]), 
	.A(\reg_array[7][15] ));
   MX2X1 U189 (.Y(n373), 
	.S0(n333), 
	.B(reg_write_data[14]), 
	.A(\reg_array[7][14] ));
   MX2X1 U190 (.Y(n374), 
	.S0(n333), 
	.B(reg_write_data[13]), 
	.A(\reg_array[7][13] ));
   MX2X1 U191 (.Y(n375), 
	.S0(n333), 
	.B(reg_write_data[12]), 
	.A(\reg_array[7][12] ));
   MX2X1 U192 (.Y(n376), 
	.S0(n333), 
	.B(reg_write_data[11]), 
	.A(\reg_array[7][11] ));
   MX2X1 U193 (.Y(n377), 
	.S0(n333), 
	.B(reg_write_data[10]), 
	.A(\reg_array[7][10] ));
   MX2X1 U194 (.Y(n378), 
	.S0(n333), 
	.B(reg_write_data[9]), 
	.A(\reg_array[7][9] ));
   MX2X1 U195 (.Y(n379), 
	.S0(n333), 
	.B(reg_write_data[8]), 
	.A(\reg_array[7][8] ));
   MX2X1 U196 (.Y(n380), 
	.S0(n333), 
	.B(reg_write_data[7]), 
	.A(\reg_array[7][7] ));
   MX2X1 U197 (.Y(n381), 
	.S0(n333), 
	.B(reg_write_data[6]), 
	.A(\reg_array[7][6] ));
   MX2X1 U198 (.Y(n382), 
	.S0(n333), 
	.B(reg_write_data[5]), 
	.A(\reg_array[7][5] ));
   MX2X1 U199 (.Y(n383), 
	.S0(n333), 
	.B(reg_write_data[4]), 
	.A(\reg_array[7][4] ));
   MX2X1 U200 (.Y(n384), 
	.S0(n333), 
	.B(reg_write_data[3]), 
	.A(\reg_array[7][3] ));
   MX2X1 U201 (.Y(n385), 
	.S0(n333), 
	.B(reg_write_data[2]), 
	.A(\reg_array[7][2] ));
   MX2X1 U202 (.Y(n386), 
	.S0(n333), 
	.B(reg_write_data[1]), 
	.A(\reg_array[7][1] ));
   MX2X1 U203 (.Y(n387), 
	.S0(n333), 
	.B(reg_write_data[0]), 
	.A(\reg_array[7][0] ));
   AND3X1 U204 (.Y(n333), 
	.C(n334), 
	.B(reg_write_dest[0]), 
	.A(reg_write_dest[2]));
   MX2X1 U205 (.Y(n388), 
	.S0(n335), 
	.B(reg_write_data[15]), 
	.A(\reg_array[3][15] ));
   MX2X1 U206 (.Y(n389), 
	.S0(n335), 
	.B(reg_write_data[14]), 
	.A(\reg_array[3][14] ));
   MX2X1 U207 (.Y(n390), 
	.S0(n335), 
	.B(reg_write_data[13]), 
	.A(\reg_array[3][13] ));
   MX2X1 U208 (.Y(n391), 
	.S0(n335), 
	.B(reg_write_data[12]), 
	.A(\reg_array[3][12] ));
   MX2X1 U209 (.Y(n392), 
	.S0(n335), 
	.B(reg_write_data[11]), 
	.A(\reg_array[3][11] ));
   MX2X1 U210 (.Y(n393), 
	.S0(n335), 
	.B(reg_write_data[10]), 
	.A(\reg_array[3][10] ));
   MX2X1 U211 (.Y(n394), 
	.S0(n335), 
	.B(reg_write_data[9]), 
	.A(\reg_array[3][9] ));
   MX2X1 U212 (.Y(n395), 
	.S0(n335), 
	.B(reg_write_data[8]), 
	.A(\reg_array[3][8] ));
   MX2X1 U213 (.Y(n396), 
	.S0(n335), 
	.B(reg_write_data[7]), 
	.A(\reg_array[3][7] ));
   MX2X1 U214 (.Y(n397), 
	.S0(n335), 
	.B(reg_write_data[6]), 
	.A(\reg_array[3][6] ));
   MX2X1 U215 (.Y(n398), 
	.S0(n335), 
	.B(reg_write_data[5]), 
	.A(\reg_array[3][5] ));
   MX2X1 U216 (.Y(n399), 
	.S0(n335), 
	.B(reg_write_data[4]), 
	.A(\reg_array[3][4] ));
   MX2X1 U217 (.Y(n400), 
	.S0(n335), 
	.B(reg_write_data[3]), 
	.A(\reg_array[3][3] ));
   MX2X1 U218 (.Y(n401), 
	.S0(n335), 
	.B(reg_write_data[2]), 
	.A(\reg_array[3][2] ));
   MX2X1 U219 (.Y(n402), 
	.S0(n335), 
	.B(reg_write_data[1]), 
	.A(\reg_array[3][1] ));
   MX2X1 U220 (.Y(n403), 
	.S0(n335), 
	.B(reg_write_data[0]), 
	.A(\reg_array[3][0] ));
   AND3X1 U221 (.Y(n335), 
	.C(n334), 
	.B(n332), 
	.A(reg_write_dest[0]));
   MX2X1 U222 (.Y(n404), 
	.S0(n336), 
	.B(reg_write_data[15]), 
	.A(\reg_array[4][15] ));
   MX2X1 U223 (.Y(n405), 
	.S0(n336), 
	.B(reg_write_data[14]), 
	.A(\reg_array[4][14] ));
   MX2X1 U224 (.Y(n406), 
	.S0(n336), 
	.B(reg_write_data[13]), 
	.A(\reg_array[4][13] ));
   MX2X1 U225 (.Y(n407), 
	.S0(n336), 
	.B(reg_write_data[12]), 
	.A(\reg_array[4][12] ));
   MX2X1 U226 (.Y(n408), 
	.S0(n336), 
	.B(reg_write_data[11]), 
	.A(\reg_array[4][11] ));
   MX2X1 U227 (.Y(n409), 
	.S0(n336), 
	.B(reg_write_data[10]), 
	.A(\reg_array[4][10] ));
   MX2X1 U228 (.Y(n410), 
	.S0(n336), 
	.B(reg_write_data[9]), 
	.A(\reg_array[4][9] ));
   MX2X1 U229 (.Y(n411), 
	.S0(n336), 
	.B(reg_write_data[8]), 
	.A(\reg_array[4][8] ));
   MX2X1 U230 (.Y(n412), 
	.S0(n336), 
	.B(reg_write_data[7]), 
	.A(\reg_array[4][7] ));
   MX2X1 U231 (.Y(n413), 
	.S0(n336), 
	.B(reg_write_data[6]), 
	.A(\reg_array[4][6] ));
   MX2X1 U232 (.Y(n414), 
	.S0(n336), 
	.B(reg_write_data[5]), 
	.A(\reg_array[4][5] ));
   MX2X1 U233 (.Y(n415), 
	.S0(n336), 
	.B(reg_write_data[4]), 
	.A(\reg_array[4][4] ));
   MX2X1 U234 (.Y(n416), 
	.S0(n336), 
	.B(reg_write_data[3]), 
	.A(\reg_array[4][3] ));
   MX2X1 U235 (.Y(n417), 
	.S0(n336), 
	.B(reg_write_data[2]), 
	.A(\reg_array[4][2] ));
   MX2X1 U236 (.Y(n418), 
	.S0(n336), 
	.B(reg_write_data[1]), 
	.A(\reg_array[4][1] ));
   MX2X1 U237 (.Y(n419), 
	.S0(n336), 
	.B(reg_write_data[0]), 
	.A(\reg_array[4][0] ));
   AND3X1 U238 (.Y(n336), 
	.C(reg_write_dest[2]), 
	.B(n337), 
	.A(n330));
   NOR2BX1 U239 (.Y(n330), 
	.B(reg_write_dest[1]), 
	.AN(reg_write_en));
   MX2X1 U240 (.Y(n420), 
	.S0(n338), 
	.B(reg_write_data[15]), 
	.A(\reg_array[6][15] ));
   MX2X1 U241 (.Y(n421), 
	.S0(n338), 
	.B(reg_write_data[14]), 
	.A(\reg_array[6][14] ));
   MX2X1 U242 (.Y(n422), 
	.S0(n338), 
	.B(reg_write_data[13]), 
	.A(\reg_array[6][13] ));
   MX2X1 U243 (.Y(n423), 
	.S0(n338), 
	.B(reg_write_data[12]), 
	.A(\reg_array[6][12] ));
   MX2X1 U244 (.Y(n424), 
	.S0(n338), 
	.B(reg_write_data[11]), 
	.A(\reg_array[6][11] ));
   MX2X1 U245 (.Y(n425), 
	.S0(n338), 
	.B(reg_write_data[10]), 
	.A(\reg_array[6][10] ));
   MX2X1 U246 (.Y(n426), 
	.S0(n338), 
	.B(reg_write_data[9]), 
	.A(\reg_array[6][9] ));
   MX2X1 U247 (.Y(n427), 
	.S0(n338), 
	.B(reg_write_data[8]), 
	.A(\reg_array[6][8] ));
   MX2X1 U248 (.Y(n428), 
	.S0(n338), 
	.B(reg_write_data[7]), 
	.A(\reg_array[6][7] ));
   MX2X1 U249 (.Y(n429), 
	.S0(n338), 
	.B(reg_write_data[6]), 
	.A(\reg_array[6][6] ));
   MX2X1 U250 (.Y(n430), 
	.S0(n338), 
	.B(reg_write_data[5]), 
	.A(\reg_array[6][5] ));
   MX2X1 U251 (.Y(n431), 
	.S0(n338), 
	.B(reg_write_data[4]), 
	.A(\reg_array[6][4] ));
   MX2X1 U252 (.Y(n432), 
	.S0(n338), 
	.B(reg_write_data[3]), 
	.A(\reg_array[6][3] ));
   MX2X1 U253 (.Y(n433), 
	.S0(n338), 
	.B(reg_write_data[2]), 
	.A(\reg_array[6][2] ));
   MX2X1 U254 (.Y(n434), 
	.S0(n338), 
	.B(reg_write_data[1]), 
	.A(\reg_array[6][1] ));
   MX2X1 U255 (.Y(n435), 
	.S0(n338), 
	.B(reg_write_data[0]), 
	.A(\reg_array[6][0] ));
   AND3X1 U256 (.Y(n338), 
	.C(n334), 
	.B(n337), 
	.A(reg_write_dest[2]));
   MX2X1 U257 (.Y(n436), 
	.S0(n339), 
	.B(reg_write_data[15]), 
	.A(\reg_array[2][15] ));
   MX2X1 U258 (.Y(n437), 
	.S0(n339), 
	.B(reg_write_data[14]), 
	.A(\reg_array[2][14] ));
   MX2X1 U259 (.Y(n438), 
	.S0(n339), 
	.B(reg_write_data[13]), 
	.A(\reg_array[2][13] ));
   MX2X1 U260 (.Y(n439), 
	.S0(n339), 
	.B(reg_write_data[12]), 
	.A(\reg_array[2][12] ));
   MX2X1 U261 (.Y(n440), 
	.S0(n339), 
	.B(reg_write_data[11]), 
	.A(\reg_array[2][11] ));
   MX2X1 U262 (.Y(n441), 
	.S0(n339), 
	.B(reg_write_data[10]), 
	.A(\reg_array[2][10] ));
   MX2X1 U263 (.Y(n442), 
	.S0(n339), 
	.B(reg_write_data[9]), 
	.A(\reg_array[2][9] ));
   MX2X1 U264 (.Y(n443), 
	.S0(n339), 
	.B(reg_write_data[8]), 
	.A(\reg_array[2][8] ));
   MX2X1 U265 (.Y(n444), 
	.S0(n339), 
	.B(reg_write_data[7]), 
	.A(\reg_array[2][7] ));
   MX2X1 U266 (.Y(n445), 
	.S0(n339), 
	.B(reg_write_data[6]), 
	.A(\reg_array[2][6] ));
   MX2X1 U267 (.Y(n446), 
	.S0(n339), 
	.B(reg_write_data[5]), 
	.A(\reg_array[2][5] ));
   MX2X1 U268 (.Y(n447), 
	.S0(n339), 
	.B(reg_write_data[4]), 
	.A(\reg_array[2][4] ));
   MX2X1 U269 (.Y(n448), 
	.S0(n339), 
	.B(reg_write_data[3]), 
	.A(\reg_array[2][3] ));
   MX2X1 U270 (.Y(n449), 
	.S0(n339), 
	.B(reg_write_data[2]), 
	.A(\reg_array[2][2] ));
   MX2X1 U271 (.Y(n450), 
	.S0(n339), 
	.B(reg_write_data[1]), 
	.A(\reg_array[2][1] ));
   MX2X1 U272 (.Y(n451), 
	.S0(n339), 
	.B(reg_write_data[0]), 
	.A(\reg_array[2][0] ));
   AND3X1 U273 (.Y(n339), 
	.C(n334), 
	.B(n332), 
	.A(n337));
   AND2X1 U274 (.Y(n334), 
	.B(reg_write_en), 
	.A(reg_write_dest[1]));
   INVX1 U275 (.Y(n332), 
	.A(reg_write_dest[2]));
   INVX1 U276 (.Y(n337), 
	.A(reg_write_dest[0]));
   INVX1 U277 (.Y(n452), 
	.A(rst));
endmodule

module hazard_detection_unit (
	decoding_op_src1, 
	decoding_op_src2, 
	ex_op_dest, 
	mem_op_dest, 
	wb_op_dest, 
	pipeline_stall_n);
   input [2:0] decoding_op_src1;
   input [2:0] decoding_op_src2;
   input [2:0] ex_op_dest;
   input [2:0] mem_op_dest;
   input [2:0] wb_op_dest;
   output pipeline_stall_n;

   // Internal wires
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;

   NOR2X1 U2 (.Y(pipeline_stall_n), 
	.B(n32), 
	.A(n31));
   AOI31X1 U3 (.Y(n32), 
	.B0(n36), 
	.A2(n35), 
	.A1(n34), 
	.A0(n33));
   AOI31X1 U4 (.Y(n36), 
	.B0(n40), 
	.A2(n39), 
	.A1(n38), 
	.A0(n37));
   OAI33X1 U5 (.Y(n40), 
	.B2(n46), 
	.B1(n45), 
	.B0(n44), 
	.A2(n43), 
	.A1(n42), 
	.A0(n41));
   XNOR2X1 U6 (.Y(n46), 
	.B(n34), 
	.A(wb_op_dest[2]));
   XNOR2X1 U7 (.Y(n45), 
	.B(n35), 
	.A(wb_op_dest[0]));
   XNOR2X1 U8 (.Y(n44), 
	.B(n33), 
	.A(wb_op_dest[1]));
   XNOR2X1 U9 (.Y(n43), 
	.B(n34), 
	.A(mem_op_dest[2]));
   XNOR2X1 U10 (.Y(n42), 
	.B(n35), 
	.A(mem_op_dest[0]));
   XNOR2X1 U11 (.Y(n41), 
	.B(n33), 
	.A(mem_op_dest[1]));
   XNOR2X1 U12 (.Y(n39), 
	.B(decoding_op_src2[1]), 
	.A(ex_op_dest[1]));
   XNOR2X1 U13 (.Y(n38), 
	.B(decoding_op_src2[2]), 
	.A(ex_op_dest[2]));
   XNOR2X1 U14 (.Y(n37), 
	.B(decoding_op_src2[0]), 
	.A(ex_op_dest[0]));
   INVX1 U15 (.Y(n35), 
	.A(decoding_op_src2[0]));
   INVX1 U16 (.Y(n34), 
	.A(decoding_op_src2[2]));
   INVX1 U17 (.Y(n33), 
	.A(decoding_op_src2[1]));
   AOI31X1 U18 (.Y(n31), 
	.B0(n50), 
	.A2(n49), 
	.A1(n48), 
	.A0(n47));
   AOI31X1 U19 (.Y(n50), 
	.B0(n54), 
	.A2(n53), 
	.A1(n52), 
	.A0(n51));
   OAI33X1 U20 (.Y(n54), 
	.B2(n60), 
	.B1(n59), 
	.B0(n58), 
	.A2(n57), 
	.A1(n56), 
	.A0(n55));
   XNOR2X1 U21 (.Y(n60), 
	.B(n48), 
	.A(wb_op_dest[2]));
   XNOR2X1 U22 (.Y(n59), 
	.B(n49), 
	.A(wb_op_dest[0]));
   XNOR2X1 U23 (.Y(n58), 
	.B(n47), 
	.A(wb_op_dest[1]));
   XNOR2X1 U24 (.Y(n57), 
	.B(n48), 
	.A(mem_op_dest[2]));
   XNOR2X1 U25 (.Y(n56), 
	.B(n49), 
	.A(mem_op_dest[0]));
   XNOR2X1 U26 (.Y(n55), 
	.B(n47), 
	.A(mem_op_dest[1]));
   XNOR2X1 U27 (.Y(n53), 
	.B(decoding_op_src1[1]), 
	.A(ex_op_dest[1]));
   XNOR2X1 U28 (.Y(n52), 
	.B(decoding_op_src1[2]), 
	.A(ex_op_dest[2]));
   XNOR2X1 U29 (.Y(n51), 
	.B(decoding_op_src1[0]), 
	.A(ex_op_dest[0]));
   INVX1 U30 (.Y(n49), 
	.A(decoding_op_src1[0]));
   INVX1 U31 (.Y(n48), 
	.A(decoding_op_src1[2]));
   INVX1 U32 (.Y(n47), 
	.A(decoding_op_src1[1]));
endmodule

module mips_16_core_top (
	clk, 
	rst, 
	pc);
   input clk;
   input rst;
   output [7:0] pc;

   // Internal wires
   wire pipeline_stall_n;
   wire branch_taken;
   wire reg_write_en;
   wire [5:0] branch_offset_imm;
   wire [56:0] ID_pipeline_reg_out;
   wire [2:0] reg_read_addr_1;
   wire [2:0] reg_read_addr_2;
   wire [15:0] reg_read_data_1;
   wire [15:0] reg_read_data_2;
   wire [2:0] decoding_op_src1;
   wire [2:0] decoding_op_src2;
   wire [37:0] EX_pipeline_reg_out;
   wire [2:0] ex_op_dest;
   wire [36:0] MEM_pipeline_reg_out;
   wire [2:0] mem_op_dest;
   wire [2:0] reg_write_dest;
   wire [15:0] reg_write_data;
   wire [2:0] wb_op_dest;

   IF_stage IF_stage_inst (.clk(clk), 
	.rst(rst), 
	.instruction_fetch_en(pipeline_stall_n), 
	.branch_offset_imm({ branch_offset_imm[5],
		branch_offset_imm[4],
		branch_offset_imm[3],
		branch_offset_imm[2],
		branch_offset_imm[1],
		branch_offset_imm[0] }), 
	.branch_taken(branch_taken), 
	.pc({ pc[7],
		pc[6],
		pc[5],
		pc[4],
		pc[3],
		pc[2],
		pc[1],
		pc[0] }), 
	.instruction ());
   ID_stage ID_stage_inst (.clk(clk), 
	.rst(rst), 
	.instruction_decode_en(pipeline_stall_n), 
	.pipeline_reg_out({ ID_pipeline_reg_out[56],
		ID_pipeline_reg_out[55],
		ID_pipeline_reg_out[54],
		ID_pipeline_reg_out[53],
		ID_pipeline_reg_out[52],
		ID_pipeline_reg_out[51],
		ID_pipeline_reg_out[50],
		ID_pipeline_reg_out[49],
		ID_pipeline_reg_out[48],
		ID_pipeline_reg_out[47],
		ID_pipeline_reg_out[46],
		ID_pipeline_reg_out[45],
		ID_pipeline_reg_out[44],
		ID_pipeline_reg_out[43],
		ID_pipeline_reg_out[42],
		ID_pipeline_reg_out[41],
		ID_pipeline_reg_out[40],
		ID_pipeline_reg_out[39],
		ID_pipeline_reg_out[38],
		ID_pipeline_reg_out[37],
		ID_pipeline_reg_out[36],
		ID_pipeline_reg_out[35],
		ID_pipeline_reg_out[34],
		ID_pipeline_reg_out[33],
		ID_pipeline_reg_out[32],
		ID_pipeline_reg_out[31],
		ID_pipeline_reg_out[30],
		ID_pipeline_reg_out[29],
		ID_pipeline_reg_out[28],
		ID_pipeline_reg_out[27],
		ID_pipeline_reg_out[26],
		ID_pipeline_reg_out[25],
		ID_pipeline_reg_out[24],
		ID_pipeline_reg_out[23],
		ID_pipeline_reg_out[22],
		ID_pipeline_reg_out[21],
		ID_pipeline_reg_out[20],
		ID_pipeline_reg_out[19],
		ID_pipeline_reg_out[18],
		ID_pipeline_reg_out[17],
		ID_pipeline_reg_out[16],
		ID_pipeline_reg_out[15],
		ID_pipeline_reg_out[14],
		ID_pipeline_reg_out[13],
		ID_pipeline_reg_out[12],
		ID_pipeline_reg_out[11],
		ID_pipeline_reg_out[10],
		ID_pipeline_reg_out[9],
		ID_pipeline_reg_out[8],
		ID_pipeline_reg_out[7],
		ID_pipeline_reg_out[6],
		ID_pipeline_reg_out[5],
		ID_pipeline_reg_out[4],
		ID_pipeline_reg_out[3],
		ID_pipeline_reg_out[2],
		ID_pipeline_reg_out[1],
		ID_pipeline_reg_out[0] }), 
	.instruction({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.branch_offset_imm({ branch_offset_imm[5],
		branch_offset_imm[4],
		branch_offset_imm[3],
		branch_offset_imm[2],
		branch_offset_imm[1],
		branch_offset_imm[0] }), 
	.branch_taken(branch_taken), 
	.reg_read_addr_1({ reg_read_addr_1[2],
		reg_read_addr_1[1],
		reg_read_addr_1[0] }), 
	.reg_read_addr_2({ reg_read_addr_2[2],
		reg_read_addr_2[1],
		reg_read_addr_2[0] }), 
	.reg_read_data_1({ reg_read_data_1[15],
		reg_read_data_1[14],
		reg_read_data_1[13],
		reg_read_data_1[12],
		reg_read_data_1[11],
		reg_read_data_1[10],
		reg_read_data_1[9],
		reg_read_data_1[8],
		reg_read_data_1[7],
		reg_read_data_1[6],
		reg_read_data_1[5],
		reg_read_data_1[4],
		reg_read_data_1[3],
		reg_read_data_1[2],
		reg_read_data_1[1],
		reg_read_data_1[0] }), 
	.reg_read_data_2({ reg_read_data_2[15],
		reg_read_data_2[14],
		reg_read_data_2[13],
		reg_read_data_2[12],
		reg_read_data_2[11],
		reg_read_data_2[10],
		reg_read_data_2[9],
		reg_read_data_2[8],
		reg_read_data_2[7],
		reg_read_data_2[6],
		reg_read_data_2[5],
		reg_read_data_2[4],
		reg_read_data_2[3],
		reg_read_data_2[2],
		reg_read_data_2[1],
		reg_read_data_2[0] }), 
	.decoding_op_src1({ decoding_op_src1[2],
		decoding_op_src1[1],
		decoding_op_src1[0] }), 
	.decoding_op_src2({ decoding_op_src2[2],
		decoding_op_src2[1],
		decoding_op_src2[0] }));
   EX_stage EX_stage_inst (.clk(clk), 
	.rst(rst), 
	.pipeline_reg_in({ ID_pipeline_reg_out[56],
		ID_pipeline_reg_out[55],
		ID_pipeline_reg_out[54],
		ID_pipeline_reg_out[53],
		ID_pipeline_reg_out[52],
		ID_pipeline_reg_out[51],
		ID_pipeline_reg_out[50],
		ID_pipeline_reg_out[49],
		ID_pipeline_reg_out[48],
		ID_pipeline_reg_out[47],
		ID_pipeline_reg_out[46],
		ID_pipeline_reg_out[45],
		ID_pipeline_reg_out[44],
		ID_pipeline_reg_out[43],
		ID_pipeline_reg_out[42],
		ID_pipeline_reg_out[41],
		ID_pipeline_reg_out[40],
		ID_pipeline_reg_out[39],
		ID_pipeline_reg_out[38],
		ID_pipeline_reg_out[37],
		ID_pipeline_reg_out[36],
		ID_pipeline_reg_out[35],
		ID_pipeline_reg_out[34],
		ID_pipeline_reg_out[33],
		ID_pipeline_reg_out[32],
		ID_pipeline_reg_out[31],
		ID_pipeline_reg_out[30],
		ID_pipeline_reg_out[29],
		ID_pipeline_reg_out[28],
		ID_pipeline_reg_out[27],
		ID_pipeline_reg_out[26],
		ID_pipeline_reg_out[25],
		ID_pipeline_reg_out[24],
		ID_pipeline_reg_out[23],
		ID_pipeline_reg_out[22],
		ID_pipeline_reg_out[21],
		ID_pipeline_reg_out[20],
		ID_pipeline_reg_out[19],
		ID_pipeline_reg_out[18],
		ID_pipeline_reg_out[17],
		ID_pipeline_reg_out[16],
		ID_pipeline_reg_out[15],
		ID_pipeline_reg_out[14],
		ID_pipeline_reg_out[13],
		ID_pipeline_reg_out[12],
		ID_pipeline_reg_out[11],
		ID_pipeline_reg_out[10],
		ID_pipeline_reg_out[9],
		ID_pipeline_reg_out[8],
		ID_pipeline_reg_out[7],
		ID_pipeline_reg_out[6],
		ID_pipeline_reg_out[5],
		ID_pipeline_reg_out[4],
		ID_pipeline_reg_out[3],
		ID_pipeline_reg_out[2],
		ID_pipeline_reg_out[1],
		ID_pipeline_reg_out[0] }), 
	.pipeline_reg_out({ EX_pipeline_reg_out[37],
		EX_pipeline_reg_out[36],
		EX_pipeline_reg_out[35],
		EX_pipeline_reg_out[34],
		EX_pipeline_reg_out[33],
		EX_pipeline_reg_out[32],
		EX_pipeline_reg_out[31],
		EX_pipeline_reg_out[30],
		EX_pipeline_reg_out[29],
		EX_pipeline_reg_out[28],
		EX_pipeline_reg_out[27],
		EX_pipeline_reg_out[26],
		EX_pipeline_reg_out[25],
		EX_pipeline_reg_out[24],
		EX_pipeline_reg_out[23],
		EX_pipeline_reg_out[22],
		EX_pipeline_reg_out[21],
		EX_pipeline_reg_out[20],
		EX_pipeline_reg_out[19],
		EX_pipeline_reg_out[18],
		EX_pipeline_reg_out[17],
		EX_pipeline_reg_out[16],
		EX_pipeline_reg_out[15],
		EX_pipeline_reg_out[14],
		EX_pipeline_reg_out[13],
		EX_pipeline_reg_out[12],
		EX_pipeline_reg_out[11],
		EX_pipeline_reg_out[10],
		EX_pipeline_reg_out[9],
		EX_pipeline_reg_out[8],
		EX_pipeline_reg_out[7],
		EX_pipeline_reg_out[6],
		EX_pipeline_reg_out[5],
		EX_pipeline_reg_out[4],
		EX_pipeline_reg_out[3],
		EX_pipeline_reg_out[2],
		EX_pipeline_reg_out[1],
		EX_pipeline_reg_out[0] }), 
	.ex_op_dest({ ex_op_dest[2],
		ex_op_dest[1],
		ex_op_dest[0] }));
   MEM_stage MEM_stage_inst (.clk(clk), 
	.rst(rst), 
	.pipeline_reg_in({ EX_pipeline_reg_out[37],
		EX_pipeline_reg_out[36],
		EX_pipeline_reg_out[35],
		EX_pipeline_reg_out[34],
		EX_pipeline_reg_out[33],
		EX_pipeline_reg_out[32],
		EX_pipeline_reg_out[31],
		EX_pipeline_reg_out[30],
		EX_pipeline_reg_out[29],
		EX_pipeline_reg_out[28],
		EX_pipeline_reg_out[27],
		EX_pipeline_reg_out[26],
		EX_pipeline_reg_out[25],
		EX_pipeline_reg_out[24],
		EX_pipeline_reg_out[23],
		EX_pipeline_reg_out[22],
		EX_pipeline_reg_out[21],
		EX_pipeline_reg_out[20],
		EX_pipeline_reg_out[19],
		EX_pipeline_reg_out[18],
		EX_pipeline_reg_out[17],
		EX_pipeline_reg_out[16],
		EX_pipeline_reg_out[15],
		EX_pipeline_reg_out[14],
		EX_pipeline_reg_out[13],
		EX_pipeline_reg_out[12],
		EX_pipeline_reg_out[11],
		EX_pipeline_reg_out[10],
		EX_pipeline_reg_out[9],
		EX_pipeline_reg_out[8],
		EX_pipeline_reg_out[7],
		EX_pipeline_reg_out[6],
		EX_pipeline_reg_out[5],
		EX_pipeline_reg_out[4],
		EX_pipeline_reg_out[3],
		EX_pipeline_reg_out[2],
		EX_pipeline_reg_out[1],
		EX_pipeline_reg_out[0] }), 
	.pipeline_reg_out({ MEM_pipeline_reg_out[36],
		MEM_pipeline_reg_out[35],
		MEM_pipeline_reg_out[34],
		MEM_pipeline_reg_out[33],
		MEM_pipeline_reg_out[32],
		MEM_pipeline_reg_out[31],
		MEM_pipeline_reg_out[30],
		MEM_pipeline_reg_out[29],
		MEM_pipeline_reg_out[28],
		MEM_pipeline_reg_out[27],
		MEM_pipeline_reg_out[26],
		MEM_pipeline_reg_out[25],
		MEM_pipeline_reg_out[24],
		MEM_pipeline_reg_out[23],
		MEM_pipeline_reg_out[22],
		MEM_pipeline_reg_out[21],
		MEM_pipeline_reg_out[20],
		MEM_pipeline_reg_out[19],
		MEM_pipeline_reg_out[18],
		MEM_pipeline_reg_out[17],
		MEM_pipeline_reg_out[16],
		MEM_pipeline_reg_out[15],
		MEM_pipeline_reg_out[14],
		MEM_pipeline_reg_out[13],
		MEM_pipeline_reg_out[12],
		MEM_pipeline_reg_out[11],
		MEM_pipeline_reg_out[10],
		MEM_pipeline_reg_out[9],
		MEM_pipeline_reg_out[8],
		MEM_pipeline_reg_out[7],
		MEM_pipeline_reg_out[6],
		MEM_pipeline_reg_out[5],
		MEM_pipeline_reg_out[4],
		MEM_pipeline_reg_out[3],
		MEM_pipeline_reg_out[2],
		MEM_pipeline_reg_out[1],
		MEM_pipeline_reg_out[0] }), 
	.mem_op_dest({ mem_op_dest[2],
		mem_op_dest[1],
		mem_op_dest[0] }));
   WB_stage WB_stage_inst (.pipeline_reg_in({ MEM_pipeline_reg_out[36],
		MEM_pipeline_reg_out[35],
		MEM_pipeline_reg_out[34],
		MEM_pipeline_reg_out[33],
		MEM_pipeline_reg_out[32],
		MEM_pipeline_reg_out[31],
		MEM_pipeline_reg_out[30],
		MEM_pipeline_reg_out[29],
		MEM_pipeline_reg_out[28],
		MEM_pipeline_reg_out[27],
		MEM_pipeline_reg_out[26],
		MEM_pipeline_reg_out[25],
		MEM_pipeline_reg_out[24],
		MEM_pipeline_reg_out[23],
		MEM_pipeline_reg_out[22],
		MEM_pipeline_reg_out[21],
		MEM_pipeline_reg_out[20],
		MEM_pipeline_reg_out[19],
		MEM_pipeline_reg_out[18],
		MEM_pipeline_reg_out[17],
		MEM_pipeline_reg_out[16],
		MEM_pipeline_reg_out[15],
		MEM_pipeline_reg_out[14],
		MEM_pipeline_reg_out[13],
		MEM_pipeline_reg_out[12],
		MEM_pipeline_reg_out[11],
		MEM_pipeline_reg_out[10],
		MEM_pipeline_reg_out[9],
		MEM_pipeline_reg_out[8],
		MEM_pipeline_reg_out[7],
		MEM_pipeline_reg_out[6],
		MEM_pipeline_reg_out[5],
		MEM_pipeline_reg_out[4],
		MEM_pipeline_reg_out[3],
		MEM_pipeline_reg_out[2],
		MEM_pipeline_reg_out[1],
		MEM_pipeline_reg_out[0] }), 
	.reg_write_en(reg_write_en), 
	.reg_write_dest({ reg_write_dest[2],
		reg_write_dest[1],
		reg_write_dest[0] }), 
	.reg_write_data({ reg_write_data[15],
		reg_write_data[14],
		reg_write_data[13],
		reg_write_data[12],
		reg_write_data[11],
		reg_write_data[10],
		reg_write_data[9],
		reg_write_data[8],
		reg_write_data[7],
		reg_write_data[6],
		reg_write_data[5],
		reg_write_data[4],
		reg_write_data[3],
		reg_write_data[2],
		reg_write_data[1],
		reg_write_data[0] }), 
	.wb_op_dest({ wb_op_dest[2],
		wb_op_dest[1],
		wb_op_dest[0] }));
   register_file register_file_inst (.clk(clk), 
	.rst(rst), 
	.reg_write_en(reg_write_en), 
	.reg_write_dest({ reg_write_dest[2],
		reg_write_dest[1],
		reg_write_dest[0] }), 
	.reg_write_data({ reg_write_data[15],
		reg_write_data[14],
		reg_write_data[13],
		reg_write_data[12],
		reg_write_data[11],
		reg_write_data[10],
		reg_write_data[9],
		reg_write_data[8],
		reg_write_data[7],
		reg_write_data[6],
		reg_write_data[5],
		reg_write_data[4],
		reg_write_data[3],
		reg_write_data[2],
		reg_write_data[1],
		reg_write_data[0] }), 
	.reg_read_addr_1({ reg_read_addr_1[2],
		reg_read_addr_1[1],
		reg_read_addr_1[0] }), 
	.reg_read_data_1({ reg_read_data_1[15],
		reg_read_data_1[14],
		reg_read_data_1[13],
		reg_read_data_1[12],
		reg_read_data_1[11],
		reg_read_data_1[10],
		reg_read_data_1[9],
		reg_read_data_1[8],
		reg_read_data_1[7],
		reg_read_data_1[6],
		reg_read_data_1[5],
		reg_read_data_1[4],
		reg_read_data_1[3],
		reg_read_data_1[2],
		reg_read_data_1[1],
		reg_read_data_1[0] }), 
	.reg_read_addr_2({ reg_read_addr_2[2],
		reg_read_addr_2[1],
		reg_read_addr_2[0] }), 
	.reg_read_data_2({ reg_read_data_2[15],
		reg_read_data_2[14],
		reg_read_data_2[13],
		reg_read_data_2[12],
		reg_read_data_2[11],
		reg_read_data_2[10],
		reg_read_data_2[9],
		reg_read_data_2[8],
		reg_read_data_2[7],
		reg_read_data_2[6],
		reg_read_data_2[5],
		reg_read_data_2[4],
		reg_read_data_2[3],
		reg_read_data_2[2],
		reg_read_data_2[1],
		reg_read_data_2[0] }));
   hazard_detection_unit hazard_detection_unit_inst (.decoding_op_src1({ decoding_op_src1[2],
		decoding_op_src1[1],
		decoding_op_src1[0] }), 
	.decoding_op_src2({ decoding_op_src2[2],
		decoding_op_src2[1],
		decoding_op_src2[0] }), 
	.ex_op_dest({ ex_op_dest[2],
		ex_op_dest[1],
		ex_op_dest[0] }), 
	.mem_op_dest({ mem_op_dest[2],
		mem_op_dest[1],
		mem_op_dest[0] }), 
	.wb_op_dest({ wb_op_dest[2],
		wb_op_dest[1],
		wb_op_dest[0] }), 
	.pipeline_stall_n(pipeline_stall_n));
endmodule

