
module instruction_mem ( clk, pc, instruction );
  input [7:0] pc;
  output [15:0] instruction;
  input clk;

  assign instruction[0] = 1'b0;
  assign instruction[1] = 1'b0;
  assign instruction[2] = 1'b0;
  assign instruction[3] = 1'b0;
  assign instruction[4] = 1'b0;
  assign instruction[5] = 1'b0;
  assign instruction[6] = 1'b0;
  assign instruction[7] = 1'b0;
  assign instruction[8] = 1'b0;
  assign instruction[9] = 1'b0;
  assign instruction[10] = 1'b0;
  assign instruction[11] = 1'b0;
  assign instruction[12] = 1'b0;
  assign instruction[13] = 1'b0;
  assign instruction[14] = 1'b0;
  assign instruction[15] = 1'b0;

endmodule


module IF_stage_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module IF_stage_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module IF_stage ( clk, rst, instruction_fetch_en, branch_offset_imm, 
        branch_taken, pc, instruction );
  input [5:0] branch_offset_imm;
  output [7:0] pc;
  output [15:0] instruction;
  input clk, rst, instruction_fetch_en, branch_taken;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n23, n2, n3;
  assign instruction[15] = 1'b0;
  assign instruction[14] = 1'b0;
  assign instruction[13] = 1'b0;
  assign instruction[12] = 1'b0;
  assign instruction[11] = 1'b0;
  assign instruction[10] = 1'b0;
  assign instruction[9] = 1'b0;
  assign instruction[8] = 1'b0;
  assign instruction[7] = 1'b0;
  assign instruction[6] = 1'b0;
  assign instruction[5] = 1'b0;
  assign instruction[4] = 1'b0;
  assign instruction[3] = 1'b0;
  assign instruction[2] = 1'b0;
  assign instruction[1] = 1'b0;
  assign instruction[0] = 1'b0;

  instruction_mem imem ( .clk(clk), .pc(pc) );
  IF_stage_DW01_inc_0 add_39 ( .A(pc), .SUM({N21, N20, N19, N18, N17, N16, N15, 
        N14}) );
  IF_stage_DW01_add_0 add_37 ( .A(pc), .B({branch_offset_imm[5], 
        branch_offset_imm[5], branch_offset_imm}), .CI(1'b0), .SUM({N13, N12, 
        N11, N10, N9, N8, N7, N6}) );
  DFFRHQX1 \pc_reg[7]  ( .D(n21), .CK(clk), .RN(n3), .Q(pc[7]) );
  DFFRHQX1 \pc_reg[4]  ( .D(n17), .CK(clk), .RN(n3), .Q(pc[4]) );
  DFFRHQX1 \pc_reg[5]  ( .D(n16), .CK(clk), .RN(n3), .Q(pc[5]) );
  DFFRHQX1 \pc_reg[6]  ( .D(n15), .CK(clk), .RN(n3), .Q(pc[6]) );
  DFFRHQX1 \pc_reg[1]  ( .D(n20), .CK(clk), .RN(n3), .Q(pc[1]) );
  DFFRHQX1 \pc_reg[2]  ( .D(n19), .CK(clk), .RN(n3), .Q(pc[2]) );
  DFFRHQX1 \pc_reg[3]  ( .D(n18), .CK(clk), .RN(n3), .Q(pc[3]) );
  DFFRHQX2 \pc_reg[0]  ( .D(n23), .CK(clk), .RN(n3), .Q(pc[0]) );
  CLKINVX3 U3 ( .A(instruction_fetch_en), .Y(n2) );
  NOR2X2 U4 ( .A(n2), .B(branch_taken), .Y(n6) );
  AND2X2 U6 ( .A(branch_taken), .B(instruction_fetch_en), .Y(n7) );
  OAI2BB1X1 U7 ( .A0N(pc[6]), .A1N(n2), .B0(n5), .Y(n15) );
  AOI22X1 U8 ( .A0(N20), .A1(n6), .B0(N12), .B1(n7), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(pc[5]), .A1N(n2), .B0(n8), .Y(n16) );
  AOI22X1 U10 ( .A0(N19), .A1(n6), .B0(N11), .B1(n7), .Y(n8) );
  OAI2BB1X1 U11 ( .A0N(pc[4]), .A1N(n2), .B0(n9), .Y(n17) );
  AOI22X1 U12 ( .A0(N18), .A1(n6), .B0(N10), .B1(n7), .Y(n9) );
  OAI2BB1X1 U13 ( .A0N(pc[3]), .A1N(n2), .B0(n10), .Y(n18) );
  AOI22X1 U14 ( .A0(N17), .A1(n6), .B0(N9), .B1(n7), .Y(n10) );
  OAI2BB1X1 U15 ( .A0N(pc[2]), .A1N(n2), .B0(n11), .Y(n19) );
  AOI22X1 U16 ( .A0(N16), .A1(n6), .B0(N8), .B1(n7), .Y(n11) );
  OAI2BB1X1 U17 ( .A0N(pc[1]), .A1N(n2), .B0(n12), .Y(n20) );
  AOI22X1 U18 ( .A0(N15), .A1(n6), .B0(N7), .B1(n7), .Y(n12) );
  OAI2BB1X1 U19 ( .A0N(pc[7]), .A1N(n2), .B0(n13), .Y(n21) );
  AOI22X1 U20 ( .A0(N21), .A1(n6), .B0(N13), .B1(n7), .Y(n13) );
  OAI2BB1X1 U21 ( .A0N(pc[0]), .A1N(n2), .B0(n14), .Y(n23) );
  AOI22X1 U22 ( .A0(N14), .A1(n6), .B0(N6), .B1(n7), .Y(n14) );
  CLKINVX3 U23 ( .A(rst), .Y(n3) );
endmodule


module ID_stage ( clk, rst, instruction_decode_en, pipeline_reg_out, 
        instruction, branch_offset_imm, branch_taken, reg_read_addr_1, 
        reg_read_addr_2, reg_read_data_1, reg_read_data_2, decoding_op_src1, 
        decoding_op_src2 );
  output [56:0] pipeline_reg_out;
  input [15:0] instruction;
  output [5:0] branch_offset_imm;
  output [2:0] reg_read_addr_1;
  output [2:0] reg_read_addr_2;
  input [15:0] reg_read_data_1;
  input [15:0] reg_read_data_2;
  output [2:0] decoding_op_src1;
  output [2:0] decoding_op_src2;
  input clk, rst, instruction_decode_en;
  output branch_taken;
  wire   write_back_en, n2, n3, n4, n5, n6, n9, n11, n12, n13, n14, n15, n16,
         n17, n18, n22, n23, n26, n27, n29, n30, n31, n32, n33, n34, n35, n37,
         n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n73, n74, n75, n78,
         n80, n1, n7, n8, n10, n19, n20, n21, n24, n25, n28, n36, n43, n49,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n76, n77, n79, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n93, n94, n95, n96, n97, n98;
  wire   [15:9] instruction_reg;
  wire   [2:0] ir_dest_with_bubble;
  wire   [2:0] ex_alu_cmd;
  wire   [15:0] ex_alu_src2;
  assign decoding_op_src1[2] = reg_read_addr_1[2];
  assign decoding_op_src1[1] = reg_read_addr_1[1];
  assign decoding_op_src1[0] = reg_read_addr_1[0];

  DFFRHQX4 \pipeline_reg_out_reg[38]  ( .D(reg_read_data_1[0]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[38]) );
  DFFRHQX1 \instruction_reg_reg[2]  ( .D(n64), .CK(clk), .RN(n8), .Q(
        branch_offset_imm[2]) );
  DFFRHQX1 \instruction_reg_reg[1]  ( .D(n49), .CK(clk), .RN(n8), .Q(
        branch_offset_imm[1]) );
  DFFRHQX1 \instruction_reg_reg[0]  ( .D(n43), .CK(clk), .RN(n8), .Q(
        branch_offset_imm[0]) );
  DFFRHQX1 \pipeline_reg_out_reg[56]  ( .D(ex_alu_cmd[2]), .CK(clk), .RN(n8), 
        .Q(pipeline_reg_out[56]) );
  DFFRHQX1 \pipeline_reg_out_reg[54]  ( .D(ex_alu_cmd[0]), .CK(clk), .RN(n8), 
        .Q(pipeline_reg_out[54]) );
  DFFRHQX2 \pipeline_reg_out_reg[55]  ( .D(ex_alu_cmd[1]), .CK(clk), .RN(n8), 
        .Q(pipeline_reg_out[55]) );
  DFFRHQX1 \pipeline_reg_out_reg[48]  ( .D(reg_read_data_1[10]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[48]) );
  DFFRHQX1 \pipeline_reg_out_reg[47]  ( .D(reg_read_data_1[9]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[47]) );
  DFFRHQX1 \pipeline_reg_out_reg[46]  ( .D(reg_read_data_1[8]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[46]) );
  DFFRHQX1 \pipeline_reg_out_reg[45]  ( .D(reg_read_data_1[7]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[45]) );
  DFFRHQX1 \pipeline_reg_out_reg[44]  ( .D(reg_read_data_1[6]), .CK(clk), .RN(
        n98), .Q(pipeline_reg_out[44]) );
  DFFRHQX1 \pipeline_reg_out_reg[43]  ( .D(reg_read_data_1[5]), .CK(clk), .RN(
        n98), .Q(pipeline_reg_out[43]) );
  DFFRHQX1 \pipeline_reg_out_reg[42]  ( .D(reg_read_data_1[4]), .CK(clk), .RN(
        n98), .Q(pipeline_reg_out[42]) );
  DFFRHQX1 \pipeline_reg_out_reg[41]  ( .D(reg_read_data_1[3]), .CK(clk), .RN(
        n7), .Q(pipeline_reg_out[41]) );
  DFFRHQX1 \pipeline_reg_out_reg[40]  ( .D(reg_read_data_1[2]), .CK(clk), .RN(
        n7), .Q(pipeline_reg_out[40]) );
  DFFRHQX1 \pipeline_reg_out_reg[52]  ( .D(reg_read_data_1[14]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[52]) );
  DFFRHQX1 \pipeline_reg_out_reg[51]  ( .D(reg_read_data_1[13]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[51]) );
  DFFRHQX1 \pipeline_reg_out_reg[50]  ( .D(reg_read_data_1[12]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[50]) );
  DFFRHQX1 \pipeline_reg_out_reg[49]  ( .D(reg_read_data_1[11]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[49]) );
  DFFRHQX1 \pipeline_reg_out_reg[39]  ( .D(reg_read_data_1[1]), .CK(clk), .RN(
        n19), .Q(pipeline_reg_out[39]) );
  DFFRHQX1 \pipeline_reg_out_reg[25]  ( .D(n77), .CK(clk), .RN(n10), .Q(
        pipeline_reg_out[25]) );
  DFFRHQX1 \pipeline_reg_out_reg[24]  ( .D(n79), .CK(clk), .RN(n10), .Q(
        pipeline_reg_out[24]) );
  DFFRHQX1 \pipeline_reg_out_reg[23]  ( .D(n81), .CK(clk), .RN(n10), .Q(
        pipeline_reg_out[23]) );
  DFFRHQX1 \pipeline_reg_out_reg[22]  ( .D(n82), .CK(clk), .RN(n10), .Q(
        pipeline_reg_out[22]) );
  DFFRHQX1 \pipeline_reg_out_reg[53]  ( .D(reg_read_data_1[15]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[53]) );
  DFFRHQX1 \pipeline_reg_out_reg[3]  ( .D(ir_dest_with_bubble[2]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[3]) );
  DFFRHQX1 \pipeline_reg_out_reg[2]  ( .D(ir_dest_with_bubble[1]), .CK(clk), 
        .RN(n19), .Q(pipeline_reg_out[2]) );
  DFFRHQX1 \pipeline_reg_out_reg[1]  ( .D(ir_dest_with_bubble[0]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[1]) );
  DFFRHQX1 \pipeline_reg_out_reg[26]  ( .D(n76), .CK(clk), .RN(n10), .Q(
        pipeline_reg_out[26]) );
  DFFRHQX1 \instruction_reg_reg[14]  ( .D(n78), .CK(clk), .RN(n7), .Q(
        instruction_reg[14]) );
  DFFRHQX1 \instruction_reg_reg[11]  ( .D(n75), .CK(clk), .RN(n7), .Q(
        instruction_reg[11]) );
  DFFRHQX1 \instruction_reg_reg[10]  ( .D(n74), .CK(clk), .RN(n7), .Q(
        instruction_reg[10]) );
  DFFRHQX1 \instruction_reg_reg[9]  ( .D(n73), .CK(clk), .RN(n7), .Q(
        instruction_reg[9]) );
  DFFRHQX1 \instruction_reg_reg[7]  ( .D(n69), .CK(clk), .RN(n7), .Q(
        reg_read_addr_1[1]) );
  DFFRHQX1 \instruction_reg_reg[6]  ( .D(n68), .CK(clk), .RN(n7), .Q(
        reg_read_addr_1[0]) );
  DFFRHQX1 \instruction_reg_reg[15]  ( .D(n80), .CK(clk), .RN(n19), .Q(
        instruction_reg[15]) );
  DFFRHQX2 \instruction_reg_reg[13]  ( .D(n72), .CK(clk), .RN(n7), .Q(
        instruction_reg[13]) );
  DFFRHQX2 \instruction_reg_reg[5]  ( .D(n67), .CK(clk), .RN(n7), .Q(
        branch_offset_imm[5]) );
  DFFRHQX2 \instruction_reg_reg[12]  ( .D(n71), .CK(clk), .RN(n7), .Q(
        instruction_reg[12]) );
  DFFRHQX2 \pipeline_reg_out_reg[27]  ( .D(ex_alu_src2[5]), .CK(clk), .RN(n10), 
        .Q(pipeline_reg_out[27]) );
  DFFRHQX2 \pipeline_reg_out_reg[28]  ( .D(ex_alu_src2[6]), .CK(clk), .RN(n10), 
        .Q(pipeline_reg_out[28]) );
  DFFRHQX2 \pipeline_reg_out_reg[29]  ( .D(ex_alu_src2[7]), .CK(clk), .RN(n10), 
        .Q(pipeline_reg_out[29]) );
  DFFRHQX2 \pipeline_reg_out_reg[32]  ( .D(ex_alu_src2[10]), .CK(clk), .RN(n10), .Q(pipeline_reg_out[32]) );
  DFFRHQX2 \pipeline_reg_out_reg[35]  ( .D(ex_alu_src2[13]), .CK(clk), .RN(n7), 
        .Q(pipeline_reg_out[35]) );
  DFFRHQX2 \pipeline_reg_out_reg[30]  ( .D(ex_alu_src2[8]), .CK(clk), .RN(n10), 
        .Q(pipeline_reg_out[30]) );
  DFFRHQX2 \pipeline_reg_out_reg[36]  ( .D(ex_alu_src2[14]), .CK(clk), .RN(n7), 
        .Q(pipeline_reg_out[36]) );
  DFFRHQX2 \pipeline_reg_out_reg[33]  ( .D(ex_alu_src2[11]), .CK(clk), .RN(n7), 
        .Q(pipeline_reg_out[33]) );
  DFFRHQX2 \pipeline_reg_out_reg[31]  ( .D(ex_alu_src2[9]), .CK(clk), .RN(n98), 
        .Q(pipeline_reg_out[31]) );
  DFFRHQX2 \pipeline_reg_out_reg[34]  ( .D(ex_alu_src2[12]), .CK(clk), .RN(n98), .Q(pipeline_reg_out[34]) );
  DFFRHQX1 \pipeline_reg_out_reg[20]  ( .D(reg_read_data_2[15]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[20]) );
  DFFRHQX1 \pipeline_reg_out_reg[19]  ( .D(reg_read_data_2[14]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[19]) );
  DFFRHQX1 \pipeline_reg_out_reg[18]  ( .D(reg_read_data_2[13]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[18]) );
  DFFRHQX1 \pipeline_reg_out_reg[17]  ( .D(reg_read_data_2[12]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[17]) );
  DFFRHQX1 \pipeline_reg_out_reg[16]  ( .D(reg_read_data_2[11]), .CK(clk), 
        .RN(n10), .Q(pipeline_reg_out[16]) );
  DFFRHQX1 \pipeline_reg_out_reg[15]  ( .D(reg_read_data_2[10]), .CK(clk), 
        .RN(n8), .Q(pipeline_reg_out[15]) );
  DFFRHQX1 \pipeline_reg_out_reg[14]  ( .D(reg_read_data_2[9]), .CK(clk), .RN(
        n10), .Q(pipeline_reg_out[14]) );
  DFFRHQX1 \pipeline_reg_out_reg[13]  ( .D(reg_read_data_2[8]), .CK(clk), .RN(
        n10), .Q(pipeline_reg_out[13]) );
  DFFRHQX1 \pipeline_reg_out_reg[12]  ( .D(reg_read_data_2[7]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[12]) );
  DFFRHQX1 \pipeline_reg_out_reg[11]  ( .D(reg_read_data_2[6]), .CK(clk), .RN(
        n19), .Q(pipeline_reg_out[11]) );
  DFFRHQX1 \pipeline_reg_out_reg[10]  ( .D(reg_read_data_2[5]), .CK(clk), .RN(
        n10), .Q(pipeline_reg_out[10]) );
  DFFRHQX1 \pipeline_reg_out_reg[9]  ( .D(reg_read_data_2[4]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[9]) );
  DFFRHQX1 \pipeline_reg_out_reg[8]  ( .D(reg_read_data_2[3]), .CK(clk), .RN(
        n19), .Q(pipeline_reg_out[8]) );
  DFFRHQX1 \pipeline_reg_out_reg[7]  ( .D(reg_read_data_2[2]), .CK(clk), .RN(
        n10), .Q(pipeline_reg_out[7]) );
  DFFRHQX1 \pipeline_reg_out_reg[6]  ( .D(reg_read_data_2[1]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[6]) );
  DFFRHQX1 \pipeline_reg_out_reg[5]  ( .D(reg_read_data_2[0]), .CK(clk), .RN(
        n8), .Q(pipeline_reg_out[5]) );
  DFFRHQX1 \instruction_reg_reg[8]  ( .D(n70), .CK(clk), .RN(n7), .Q(
        reg_read_addr_1[2]) );
  DFFRHQX1 \instruction_reg_reg[4]  ( .D(n66), .CK(clk), .RN(n7), .Q(
        branch_offset_imm[4]) );
  DFFRHQX1 \instruction_reg_reg[3]  ( .D(n65), .CK(clk), .RN(n7), .Q(
        branch_offset_imm[3]) );
  DFFRHQX1 \pipeline_reg_out_reg[21]  ( .D(n93), .CK(clk), .RN(n10), .Q(
        pipeline_reg_out[21]) );
  DFFRHQX1 \pipeline_reg_out_reg[4]  ( .D(write_back_en), .CK(clk), .RN(n8), 
        .Q(pipeline_reg_out[4]) );
  DFFRHQX1 \pipeline_reg_out_reg[0]  ( .D(n85), .CK(clk), .RN(n19), .Q(
        pipeline_reg_out[0]) );
  DFFRHQX2 \pipeline_reg_out_reg[37]  ( .D(ex_alu_src2[15]), .CK(clk), .RN(n8), 
        .Q(pipeline_reg_out[37]) );
  INVX4 U3 ( .A(rst), .Y(n10) );
  INVX4 U4 ( .A(rst), .Y(n8) );
  NAND2X2 U5 ( .A(branch_offset_imm[5]), .B(n27), .Y(n1) );
  OAI21XL U6 ( .A0(n52), .A1(n89), .B0(n53), .Y(n50) );
  CLKINVX3 U7 ( .A(n28), .Y(n24) );
  INVX1 U8 ( .A(n20), .Y(n28) );
  INVX1 U9 ( .A(n24), .Y(n25) );
  INVX1 U10 ( .A(n20), .Y(n36) );
  NOR2X1 U11 ( .A(n84), .B(n86), .Y(n3) );
  OAI31X1 U12 ( .A0(n46), .A1(n6), .A2(n84), .B0(n47), .Y(ex_alu_cmd[2]) );
  NAND2X1 U13 ( .A(n86), .B(n7), .Y(n46) );
  NOR4BX1 U14 ( .AN(n19), .B(n3), .C(n4), .D(n5), .Y(write_back_en) );
  AND3X2 U15 ( .A(n6), .B(n86), .C(n84), .Y(n5) );
  NOR2X1 U16 ( .A(n87), .B(n88), .Y(n6) );
  INVX1 U17 ( .A(n21), .Y(n20) );
  INVX1 U18 ( .A(instruction_decode_en), .Y(n21) );
  NAND4X1 U19 ( .A(n6), .B(n42), .C(n84), .D(n7), .Y(n47) );
  NOR2X1 U20 ( .A(n87), .B(n44), .Y(n41) );
  INVX1 U21 ( .A(n44), .Y(n84) );
  INVX1 U22 ( .A(n42), .Y(n86) );
  AND2X2 U23 ( .A(n39), .B(n88), .Y(n4) );
  OAI31X1 U24 ( .A0(n46), .A1(n88), .A2(n41), .B0(n47), .Y(ex_alu_cmd[0]) );
  OAI21XL U25 ( .A0(n48), .A1(n46), .B0(n47), .Y(ex_alu_cmd[1]) );
  AOI22X1 U26 ( .A0(n6), .A1(n44), .B0(n88), .B1(n87), .Y(n48) );
  INVX1 U27 ( .A(n2), .Y(n85) );
  CLKINVX3 U28 ( .A(rst), .Y(n7) );
  INVX1 U29 ( .A(rst), .Y(n19) );
  NOR2X1 U30 ( .A(n33), .B(n50), .Y(decoding_op_src2[2]) );
  NOR2X1 U31 ( .A(n35), .B(n50), .Y(decoding_op_src2[0]) );
  NOR2X1 U32 ( .A(n34), .B(n50), .Y(decoding_op_src2[1]) );
  CLKINVX3 U33 ( .A(n27), .Y(n83) );
  INVX1 U34 ( .A(n51), .Y(n93) );
  INVX1 U35 ( .A(n38), .Y(n88) );
  INVX1 U36 ( .A(n45), .Y(n87) );
  NOR2X1 U37 ( .A(n94), .B(n25), .Y(n44) );
  NOR3X1 U38 ( .A(n86), .B(n44), .C(n45), .Y(n39) );
  NOR2X1 U39 ( .A(n89), .B(n25), .Y(n42) );
  NAND3X1 U40 ( .A(n38), .B(n7), .C(n39), .Y(n2) );
  NOR4BX1 U41 ( .AN(n60), .B(n61), .C(reg_read_data_1[11]), .D(
        reg_read_data_1[10]), .Y(n59) );
  OR3XL U42 ( .A(reg_read_data_1[12]), .B(reg_read_data_1[14]), .C(
        reg_read_data_1[13]), .Y(n61) );
  NOR4BX1 U43 ( .AN(n55), .B(n89), .C(reg_read_data_1[0]), .D(n62), .Y(n60) );
  AOI31X1 U44 ( .A0(n95), .A1(n97), .A2(n96), .B0(n28), .Y(n62) );
  AND4X2 U45 ( .A(n56), .B(n57), .C(n58), .D(n59), .Y(branch_taken) );
  NOR2X1 U46 ( .A(reg_read_data_1[1]), .B(reg_read_data_1[15]), .Y(n56) );
  NOR3X1 U47 ( .A(reg_read_data_1[2]), .B(reg_read_data_1[4]), .C(
        reg_read_data_1[3]), .Y(n57) );
  NOR4BX1 U48 ( .AN(n63), .B(reg_read_data_1[6]), .C(reg_read_data_1[5]), .D(
        reg_read_data_1[7]), .Y(n58) );
  OAI2BB1XL U49 ( .A0N(reg_read_data_2[5]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[5]) );
  OAI2BB1XL U50 ( .A0N(reg_read_data_2[6]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[6]) );
  OAI2BB1XL U51 ( .A0N(reg_read_data_2[7]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[7]) );
  OAI2BB1XL U52 ( .A0N(reg_read_data_2[8]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[8]) );
  OAI2BB1XL U53 ( .A0N(reg_read_data_2[9]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[9]) );
  OAI2BB1XL U54 ( .A0N(reg_read_data_2[10]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[10]) );
  OAI2BB1XL U55 ( .A0N(reg_read_data_2[11]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[11]) );
  OAI2BB1XL U56 ( .A0N(reg_read_data_2[12]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[12]) );
  OAI2BB1XL U57 ( .A0N(reg_read_data_2[13]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[13]) );
  OAI2BB1XL U58 ( .A0N(reg_read_data_2[14]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[14]) );
  OAI2BB1XL U59 ( .A0N(reg_read_data_2[15]), .A1N(n83), .B0(n1), .Y(
        ex_alu_src2[15]) );
  NOR2X1 U60 ( .A(reg_read_data_1[9]), .B(reg_read_data_1[8]), .Y(n63) );
  NOR2X1 U61 ( .A(n21), .B(n95), .Y(ir_dest_with_bubble[2]) );
  NOR2X1 U62 ( .A(n25), .B(n97), .Y(ir_dest_with_bubble[0]) );
  NOR2X1 U63 ( .A(n21), .B(n96), .Y(ir_dest_with_bubble[1]) );
  INVX1 U64 ( .A(n35), .Y(reg_read_addr_2[0]) );
  INVX1 U65 ( .A(n34), .Y(reg_read_addr_2[1]) );
  INVX1 U66 ( .A(n33), .Y(reg_read_addr_2[2]) );
  OAI21X2 U67 ( .A0(n37), .A1(rst), .B0(n2), .Y(n27) );
  AOI211X1 U68 ( .A0(n3), .A1(n6), .B0(n4), .C0(n40), .Y(n37) );
  AND3X2 U69 ( .A(n41), .B(n42), .C(n88), .Y(n40) );
  NAND4X1 U70 ( .A(instruction_reg[12]), .B(instruction_reg[15]), .C(
        instruction_reg[13]), .D(n94), .Y(n51) );
  AOI22X1 U71 ( .A0(n51), .A1(branch_offset_imm[5]), .B0(instruction_reg[11]), 
        .B1(n93), .Y(n33) );
  AOI22X1 U72 ( .A0(n51), .A1(branch_offset_imm[3]), .B0(instruction_reg[9]), 
        .B1(n93), .Y(n35) );
  AOI22X1 U73 ( .A0(n51), .A1(branch_offset_imm[4]), .B0(instruction_reg[10]), 
        .B1(n93), .Y(n34) );
  NAND2X1 U74 ( .A(instruction_reg[12]), .B(n24), .Y(n38) );
  NAND2X1 U75 ( .A(instruction_reg[13]), .B(n24), .Y(n45) );
  INVX1 U76 ( .A(n26), .Y(n82) );
  AOI22X1 U77 ( .A0(n27), .A1(branch_offset_imm[0]), .B0(reg_read_data_2[0]), 
        .B1(n83), .Y(n26) );
  INVX1 U78 ( .A(n29), .Y(n81) );
  AOI22X1 U79 ( .A0(n27), .A1(branch_offset_imm[1]), .B0(reg_read_data_2[1]), 
        .B1(n83), .Y(n29) );
  INVX1 U80 ( .A(n30), .Y(n79) );
  AOI22X1 U81 ( .A0(n27), .A1(branch_offset_imm[2]), .B0(reg_read_data_2[2]), 
        .B1(n83), .Y(n30) );
  INVX1 U82 ( .A(n31), .Y(n77) );
  AOI22X1 U83 ( .A0(n27), .A1(branch_offset_imm[3]), .B0(reg_read_data_2[3]), 
        .B1(n83), .Y(n31) );
  INVX1 U84 ( .A(n32), .Y(n76) );
  AOI22X1 U85 ( .A0(n27), .A1(branch_offset_imm[4]), .B0(reg_read_data_2[4]), 
        .B1(n83), .Y(n32) );
  NOR3X1 U86 ( .A(instruction_reg[12]), .B(instruction_reg[13]), .C(n94), .Y(
        n55) );
  INVX1 U87 ( .A(instruction_reg[14]), .Y(n94) );
  INVX1 U88 ( .A(instruction_reg[15]), .Y(n89) );
  OR4X2 U89 ( .A(instruction_reg[12]), .B(instruction_reg[13]), .C(
        instruction_reg[14]), .D(instruction_reg[15]), .Y(n53) );
  AOI21X1 U90 ( .A0(n54), .A1(n94), .B0(n55), .Y(n52) );
  XOR2X1 U91 ( .A(instruction_reg[13]), .B(instruction_reg[12]), .Y(n54) );
  INVX1 U92 ( .A(n9), .Y(n43) );
  AOI22X1 U93 ( .A0(n36), .A1(branch_offset_imm[0]), .B0(instruction[0]), .B1(
        n20), .Y(n9) );
  OAI2BB2X1 U94 ( .B0(instruction_decode_en), .B1(n89), .A0N(instruction[15]), 
        .A1N(n24), .Y(n80) );
  OAI2BB2X1 U95 ( .B0(instruction_decode_en), .B1(n94), .A0N(instruction[14]), 
        .A1N(n24), .Y(n78) );
  OAI2BB2X1 U96 ( .B0(n20), .B1(n95), .A0N(instruction[11]), .A1N(n24), .Y(n75) );
  OAI2BB2X1 U97 ( .B0(n20), .B1(n97), .A0N(instruction[9]), .A1N(n24), .Y(n73)
         );
  OAI2BB2X1 U98 ( .B0(n20), .B1(n96), .A0N(instruction[10]), .A1N(n24), .Y(n74) );
  INVX1 U99 ( .A(n18), .Y(n70) );
  AOI22X1 U100 ( .A0(instruction[8]), .A1(n24), .B0(reg_read_addr_1[2]), .B1(
        n25), .Y(n18) );
  INVX1 U101 ( .A(n15), .Y(n67) );
  AOI22X1 U102 ( .A0(n36), .A1(branch_offset_imm[5]), .B0(instruction[5]), 
        .B1(n24), .Y(n15) );
  INVX1 U103 ( .A(n22), .Y(n71) );
  AOI22X1 U104 ( .A0(n25), .A1(instruction_reg[12]), .B0(instruction[12]), 
        .B1(n20), .Y(n22) );
  INVX1 U105 ( .A(n23), .Y(n72) );
  AOI22X1 U106 ( .A0(n25), .A1(instruction_reg[13]), .B0(instruction[13]), 
        .B1(n24), .Y(n23) );
  INVX1 U107 ( .A(n13), .Y(n65) );
  AOI22X1 U108 ( .A0(n28), .A1(branch_offset_imm[3]), .B0(instruction[3]), 
        .B1(instruction_decode_en), .Y(n13) );
  INVX1 U109 ( .A(n14), .Y(n66) );
  AOI22X1 U110 ( .A0(n36), .A1(branch_offset_imm[4]), .B0(instruction[4]), 
        .B1(n24), .Y(n14) );
  INVX1 U111 ( .A(n11), .Y(n49) );
  AOI22X1 U112 ( .A0(n21), .A1(branch_offset_imm[1]), .B0(instruction[1]), 
        .B1(n24), .Y(n11) );
  INVX1 U113 ( .A(n12), .Y(n64) );
  AOI22X1 U114 ( .A0(n25), .A1(branch_offset_imm[2]), .B0(instruction[2]), 
        .B1(n24), .Y(n12) );
  INVX1 U115 ( .A(n16), .Y(n68) );
  AOI22X1 U116 ( .A0(instruction[6]), .A1(n24), .B0(reg_read_addr_1[0]), .B1(
        n21), .Y(n16) );
  INVX1 U117 ( .A(n17), .Y(n69) );
  AOI22X1 U118 ( .A0(instruction[7]), .A1(n24), .B0(reg_read_addr_1[1]), .B1(
        n21), .Y(n17) );
  INVX1 U119 ( .A(rst), .Y(n98) );
  INVX1 U120 ( .A(instruction_reg[11]), .Y(n95) );
  INVX1 U121 ( .A(instruction_reg[9]), .Y(n97) );
  INVX1 U122 ( .A(instruction_reg[10]), .Y(n96) );
endmodule


module alu_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [15:0] A;
  input [15:0] SH;
  output [15:0] B;
  input DATA_TC, SH_TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  NOR2X4 U3 ( .A(SH[0]), .B(SH[1]), .Y(n3) );
  NOR2X4 U4 ( .A(n25), .B(SH[1]), .Y(n4) );
  OR2X2 U5 ( .A(n57), .B(n22), .Y(n5) );
  OAI22XL U6 ( .A0(n26), .A1(n20), .B0(n27), .B1(n5), .Y(B[9]) );
  AOI221XL U7 ( .A0(A[4]), .A1(n4), .B0(A[3]), .B1(n3), .C0(n43), .Y(n41) );
  AOI22XL U8 ( .A0(A[13]), .A1(n4), .B0(A[12]), .B1(n3), .Y(n70) );
  AOI22XL U9 ( .A0(A[12]), .A1(n4), .B0(A[11]), .B1(n3), .Y(n58) );
  AOI22XL U10 ( .A0(A[2]), .A1(n4), .B0(A[1]), .B1(n3), .Y(n55) );
  AOI22XL U11 ( .A0(A[3]), .A1(n4), .B0(A[2]), .B1(n3), .Y(n51) );
  NAND2XL U12 ( .A(n3), .B(A[15]), .Y(n31) );
  AOI22XL U13 ( .A0(A[8]), .A1(n4), .B0(A[7]), .B1(n3), .Y(n42) );
  AOI22XL U14 ( .A0(A[6]), .A1(n4), .B0(A[5]), .B1(n3), .Y(n54) );
  AOI22XL U15 ( .A0(A[7]), .A1(n4), .B0(A[6]), .B1(n3), .Y(n49) );
  AOI22XL U16 ( .A0(A[10]), .A1(n4), .B0(A[9]), .B1(n3), .Y(n56) );
  AOI22XL U17 ( .A0(A[11]), .A1(n4), .B0(A[10]), .B1(n3), .Y(n59) );
  AOI22XL U18 ( .A0(A[5]), .A1(n4), .B0(A[4]), .B1(n3), .Y(n62) );
  AOI22XL U19 ( .A0(A[9]), .A1(n4), .B0(A[8]), .B1(n3), .Y(n65) );
  AOI22XL U20 ( .A0(A[1]), .A1(n4), .B0(A[0]), .B1(n3), .Y(n63) );
  CLKINVX3 U21 ( .A(n47), .Y(n20) );
  CLKINVX3 U22 ( .A(n44), .Y(n23) );
  CLKINVX3 U23 ( .A(n50), .Y(n24) );
  INVX1 U24 ( .A(n40), .Y(n19) );
  INVX1 U25 ( .A(n70), .Y(n6) );
  INVX1 U26 ( .A(n65), .Y(n10) );
  INVX1 U27 ( .A(n56), .Y(n9) );
  INVX1 U28 ( .A(n59), .Y(n8) );
  INVX1 U29 ( .A(n58), .Y(n7) );
  INVX1 U30 ( .A(n62), .Y(n15) );
  INVX1 U31 ( .A(n54), .Y(n13) );
  INVX1 U32 ( .A(n49), .Y(n12) );
  INVX1 U33 ( .A(A[2]), .Y(n18) );
  INVX1 U34 ( .A(SH[0]), .Y(n25) );
  INVX1 U35 ( .A(n42), .Y(n11) );
  INVX1 U36 ( .A(SH[2]), .Y(n22) );
  INVX1 U37 ( .A(A[5]), .Y(n14) );
  INVX1 U38 ( .A(A[3]), .Y(n17) );
  INVX1 U39 ( .A(A[4]), .Y(n16) );
  INVX1 U40 ( .A(SH[15]), .Y(n21) );
  OAI22X1 U41 ( .A0(n28), .A1(n20), .B0(n29), .B1(n5), .Y(B[8]) );
  OAI222XL U42 ( .A0(n30), .A1(n5), .B0(n31), .B1(n32), .C0(n33), .C1(n20), 
        .Y(B[7]) );
  OAI222XL U43 ( .A0(n34), .A1(n5), .B0(n35), .B1(n32), .C0(n36), .C1(n20), 
        .Y(B[6]) );
  OAI222XL U44 ( .A0(n26), .A1(n5), .B0(n27), .B1(n32), .C0(n37), .C1(n20), 
        .Y(B[5]) );
  OAI222XL U45 ( .A0(n28), .A1(n5), .B0(n29), .B1(n32), .C0(n38), .C1(n20), 
        .Y(B[4]) );
  OAI222XL U46 ( .A0(n39), .A1(n40), .B0(n41), .B1(n20), .C0(n33), .C1(n5), 
        .Y(B[3]) );
  AOI221X1 U47 ( .A0(n24), .A1(A[10]), .B0(n23), .B1(A[9]), .C0(n11), .Y(n33)
         );
  OAI2BB2X1 U48 ( .B0(n44), .B1(n14), .A0N(n24), .A1N(A[6]), .Y(n43) );
  OAI221XL U49 ( .A0(n35), .A1(n45), .B0(n34), .B1(n32), .C0(n46), .Y(B[2]) );
  AOI2BB2X1 U50 ( .B0(n47), .B1(n48), .A0N(n5), .A1N(n36), .Y(n46) );
  AOI221X1 U51 ( .A0(n24), .A1(A[9]), .B0(n23), .B1(A[8]), .C0(n12), .Y(n36)
         );
  OAI221XL U52 ( .A0(n50), .A1(n14), .B0(n44), .B1(n16), .C0(n51), .Y(n48) );
  OAI221XL U53 ( .A0(n27), .A1(n45), .B0(n26), .B1(n32), .C0(n52), .Y(B[1]) );
  AOI2BB2X1 U54 ( .B0(n47), .B1(n53), .A0N(n5), .A1N(n37), .Y(n52) );
  AOI221X1 U55 ( .A0(n24), .A1(A[8]), .B0(n23), .B1(A[7]), .C0(n13), .Y(n37)
         );
  OAI221XL U56 ( .A0(n50), .A1(n16), .B0(n44), .B1(n17), .C0(n55), .Y(n53) );
  AOI221X1 U57 ( .A0(n24), .A1(A[12]), .B0(n23), .B1(A[11]), .C0(n9), .Y(n26)
         );
  NOR2X1 U58 ( .A(n20), .B(n31), .Y(B[15]) );
  NOR2X1 U59 ( .A(n35), .B(n20), .Y(B[14]) );
  NOR2X1 U60 ( .A(n27), .B(n20), .Y(B[13]) );
  AOI222X1 U61 ( .A0(n4), .A1(A[14]), .B0(n23), .B1(A[15]), .C0(n3), .C1(A[13]), .Y(n27) );
  NOR2X1 U62 ( .A(n29), .B(n20), .Y(B[12]) );
  NOR2X1 U63 ( .A(n39), .B(n57), .Y(B[11]) );
  MX2X1 U64 ( .A(n31), .B(n30), .S0(n22), .Y(n39) );
  AOI221X1 U65 ( .A0(A[14]), .A1(n24), .B0(n23), .B1(A[13]), .C0(n7), .Y(n30)
         );
  OAI22X1 U66 ( .A0(n34), .A1(n20), .B0(n35), .B1(n5), .Y(B[10]) );
  AOI22X1 U67 ( .A0(A[14]), .A1(n3), .B0(A[15]), .B1(n4), .Y(n35) );
  AOI221X1 U68 ( .A0(A[13]), .A1(n24), .B0(n23), .B1(A[12]), .C0(n8), .Y(n34)
         );
  OAI221XL U69 ( .A0(n29), .A1(n45), .B0(n28), .B1(n32), .C0(n60), .Y(B[0]) );
  AOI2BB2X1 U70 ( .B0(n47), .B1(n61), .A0N(n5), .A1N(n38), .Y(n60) );
  AOI221X1 U71 ( .A0(n24), .A1(A[7]), .B0(n23), .B1(A[6]), .C0(n15), .Y(n38)
         );
  OAI221XL U72 ( .A0(n50), .A1(n17), .B0(n44), .B1(n18), .C0(n63), .Y(n61) );
  NOR2X1 U73 ( .A(n57), .B(SH[2]), .Y(n47) );
  NAND3BX1 U74 ( .AN(SH[3]), .B(n21), .C(n64), .Y(n57) );
  NAND2X1 U75 ( .A(n19), .B(n22), .Y(n32) );
  AOI221X1 U76 ( .A0(n24), .A1(A[11]), .B0(n23), .B1(A[10]), .C0(n10), .Y(n28)
         );
  NAND2X1 U77 ( .A(n19), .B(SH[2]), .Y(n45) );
  NAND3X1 U78 ( .A(SH[3]), .B(n21), .C(n64), .Y(n40) );
  AND4X1 U79 ( .A(n66), .B(n67), .C(n68), .D(n69), .Y(n64) );
  NOR3X1 U80 ( .A(SH[7]), .B(SH[9]), .C(SH[8]), .Y(n69) );
  NOR3X1 U81 ( .A(SH[4]), .B(SH[6]), .C(SH[5]), .Y(n68) );
  NOR3X1 U82 ( .A(SH[12]), .B(SH[14]), .C(SH[13]), .Y(n67) );
  NOR2X1 U83 ( .A(SH[11]), .B(SH[10]), .Y(n66) );
  AOI221X1 U84 ( .A0(A[15]), .A1(n24), .B0(n23), .B1(A[14]), .C0(n6), .Y(n29)
         );
  NAND2X1 U85 ( .A(n25), .B(SH[1]), .Y(n44) );
  NAND2X1 U86 ( .A(SH[0]), .B(SH[1]), .Y(n50) );
endmodule


module alu_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [15:0] A;
  input [15:0] SH;
  output [15:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[6][15] , \ML_int[6][14] , \ML_int[6][13] , \ML_int[6][12] ,
         \ML_int[6][11] , \ML_int[6][10] , \ML_int[6][9] , \ML_int[6][8] ,
         \ML_int[6][7] , \ML_int[6][6] , \ML_int[6][5] , \ML_int[6][4] ,
         \ML_int[6][3] , \ML_int[6][2] , \ML_int[6][1] , \ML_int[6][0] , n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [4:0] SHMAG;
  assign B[15] = \ML_int[6][15] ;
  assign B[14] = \ML_int[6][14] ;
  assign B[13] = \ML_int[6][13] ;
  assign B[12] = \ML_int[6][12] ;
  assign B[11] = \ML_int[6][11] ;
  assign B[10] = \ML_int[6][10] ;
  assign B[9] = \ML_int[6][9] ;
  assign B[8] = \ML_int[6][8] ;
  assign B[7] = \ML_int[6][7] ;
  assign B[6] = \ML_int[6][6] ;
  assign B[5] = \ML_int[6][5] ;
  assign B[4] = \ML_int[6][4] ;
  assign B[3] = \ML_int[6][3] ;
  assign B[2] = \ML_int[6][2] ;
  assign B[1] = \ML_int[6][1] ;
  assign B[0] = \ML_int[6][0] ;

  MX2X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S0(n8), .Y(\ML_int[1][1] ) );
  MX2X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S0(n8), .Y(\ML_int[1][15] ) );
  MX2X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S0(n8), .Y(\ML_int[1][14] ) );
  MX2X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S0(n8), .Y(\ML_int[1][13] ) );
  MX2X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S0(n8), .Y(\ML_int[1][12] ) );
  MX2X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S0(n9), .Y(
        \ML_int[2][3] ) );
  MX2X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S0(n9), .Y(
        \ML_int[2][2] ) );
  MX2X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S0(n8), .Y(\ML_int[1][5] ) );
  MX2X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S0(n8), .Y(\ML_int[1][4] ) );
  MX2X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S0(n8), .Y(\ML_int[1][11] ) );
  MX2X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S0(n8), .Y(\ML_int[1][9] ) );
  MX2X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S0(n8), .Y(\ML_int[1][10] ) );
  MX2X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S0(n8), .Y(\ML_int[1][8] ) );
  MX2X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S0(n8), .Y(\ML_int[1][7] ) );
  MX2X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S0(n8), .Y(\ML_int[1][6] ) );
  MX2X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S0(n8), .Y(\ML_int[1][3] ) );
  MX2X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S0(n8), .Y(\ML_int[1][2] ) );
  MX2X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S0(n9), .Y(
        \ML_int[2][15] ) );
  MX2X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S0(n10), .Y(
        \ML_int[3][15] ) );
  MX2X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S0(n11), .Y(
        \ML_int[4][15] ) );
  MX2X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S0(n9), .Y(
        \ML_int[2][14] ) );
  MX2X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S0(n10), .Y(
        \ML_int[3][14] ) );
  MX2X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S0(n11), .Y(
        \ML_int[4][14] ) );
  MX2X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S0(n9), .Y(
        \ML_int[2][13] ) );
  MX2X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S0(n10), .Y(
        \ML_int[3][13] ) );
  MX2X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S0(n11), .Y(
        \ML_int[4][13] ) );
  MX2X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S0(n9), .Y(
        \ML_int[2][12] ) );
  MX2X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S0(n10), .Y(
        \ML_int[3][12] ) );
  MX2X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S0(n11), .Y(
        \ML_int[4][12] ) );
  MX2X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S0(n10), .Y(
        \ML_int[3][7] ) );
  MX2X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S0(n10), .Y(
        \ML_int[3][6] ) );
  MX2X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S0(n10), .Y(
        \ML_int[3][5] ) );
  MX2X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S0(n10), .Y(
        \ML_int[3][4] ) );
  MX2X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S0(n9), .Y(
        \ML_int[2][7] ) );
  MX2X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S0(n9), .Y(
        \ML_int[2][6] ) );
  MX2X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S0(n9), .Y(
        \ML_int[2][5] ) );
  MX2X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S0(n9), .Y(
        \ML_int[2][4] ) );
  MX2X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S0(n9), .Y(
        \ML_int[2][11] ) );
  MX2X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S0(n9), .Y(
        \ML_int[2][10] ) );
  MX2X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S0(n9), .Y(
        \ML_int[2][9] ) );
  MX2X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S0(n9), .Y(
        \ML_int[2][8] ) );
  NAND2X2 U3 ( .A(n7), .B(SHMAG[3]), .Y(n16) );
  NOR2XL U4 ( .A(n16), .B(n20), .Y(\ML_int[6][0] ) );
  NOR2XL U5 ( .A(n16), .B(n19), .Y(\ML_int[6][1] ) );
  NOR2XL U6 ( .A(n16), .B(n18), .Y(\ML_int[6][2] ) );
  NOR2XL U7 ( .A(n16), .B(n17), .Y(\ML_int[6][3] ) );
  NOR2BXL U8 ( .AN(\ML_int[3][4] ), .B(n16), .Y(\ML_int[6][4] ) );
  NOR2BXL U9 ( .AN(\ML_int[3][5] ), .B(n16), .Y(\ML_int[6][5] ) );
  NOR2BXL U10 ( .AN(\ML_int[3][6] ), .B(n16), .Y(\ML_int[6][6] ) );
  NOR2BXL U11 ( .AN(\ML_int[3][7] ), .B(n16), .Y(\ML_int[6][7] ) );
  CLKINVX3 U12 ( .A(SHMAG[1]), .Y(n9) );
  CLKINVX3 U13 ( .A(SHMAG[2]), .Y(n10) );
  CLKINVX3 U14 ( .A(SHMAG[0]), .Y(n8) );
  CLKINVX3 U15 ( .A(SHMAG[3]), .Y(n11) );
  MXI2X1 U16 ( .A(n3), .B(n20), .S0(n11), .Y(\ML_int[4][8] ) );
  MXI2X1 U17 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S0(n10), .Y(n3) );
  MXI2X1 U18 ( .A(n4), .B(n19), .S0(n11), .Y(\ML_int[4][9] ) );
  MXI2X1 U19 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S0(n10), .Y(n4) );
  MXI2X1 U20 ( .A(n5), .B(n18), .S0(n11), .Y(\ML_int[4][10] ) );
  MXI2X1 U21 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S0(n10), .Y(n5) );
  MXI2X1 U22 ( .A(n6), .B(n17), .S0(n11), .Y(\ML_int[4][11] ) );
  MXI2X1 U23 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S0(n10), .Y(n6) );
  INVX1 U24 ( .A(SH[7]), .Y(n12) );
  INVX1 U25 ( .A(SH[5]), .Y(n14) );
  INVX1 U26 ( .A(SH[6]), .Y(n13) );
  BUFX3 U27 ( .A(n15), .Y(n7) );
  NOR2BX1 U28 ( .AN(SHMAG[4]), .B(SH[15]), .Y(n15) );
  AND2X1 U29 ( .A(\ML_int[4][9] ), .B(n7), .Y(\ML_int[6][9] ) );
  AND2X1 U30 ( .A(\ML_int[4][8] ), .B(n7), .Y(\ML_int[6][8] ) );
  AND2X1 U31 ( .A(\ML_int[4][15] ), .B(n7), .Y(\ML_int[6][15] ) );
  AND2X1 U32 ( .A(\ML_int[4][14] ), .B(n7), .Y(\ML_int[6][14] ) );
  AND2X1 U33 ( .A(\ML_int[4][13] ), .B(n7), .Y(\ML_int[6][13] ) );
  AND2X1 U34 ( .A(\ML_int[4][12] ), .B(n7), .Y(\ML_int[6][12] ) );
  AND2X1 U35 ( .A(\ML_int[4][11] ), .B(n7), .Y(\ML_int[6][11] ) );
  AND2X1 U36 ( .A(\ML_int[4][10] ), .B(n7), .Y(\ML_int[6][10] ) );
  AOI21X1 U37 ( .A0(SH[3]), .A1(n21), .B0(n22), .Y(SHMAG[3]) );
  AOI21X1 U38 ( .A0(SH[4]), .A1(n21), .B0(n22), .Y(SHMAG[4]) );
  NAND2X1 U39 ( .A(\ML_int[2][3] ), .B(SHMAG[2]), .Y(n17) );
  NAND2X1 U40 ( .A(\ML_int[2][2] ), .B(SHMAG[2]), .Y(n18) );
  NAND2X1 U41 ( .A(\ML_int[2][1] ), .B(SHMAG[2]), .Y(n19) );
  NAND2X1 U42 ( .A(\ML_int[2][0] ), .B(SHMAG[2]), .Y(n20) );
  AOI21X1 U43 ( .A0(SH[2]), .A1(n21), .B0(n22), .Y(SHMAG[2]) );
  AND2X1 U44 ( .A(\ML_int[1][1] ), .B(SHMAG[1]), .Y(\ML_int[2][1] ) );
  AND2X1 U45 ( .A(\ML_int[1][0] ), .B(SHMAG[1]), .Y(\ML_int[2][0] ) );
  AOI21X1 U46 ( .A0(SH[1]), .A1(n21), .B0(n22), .Y(SHMAG[1]) );
  AND2X1 U47 ( .A(A[0]), .B(SHMAG[0]), .Y(\ML_int[1][0] ) );
  AOI21X1 U48 ( .A0(SH[0]), .A1(n21), .B0(n22), .Y(SHMAG[0]) );
  AOI2BB1X1 U49 ( .A0N(n23), .A1N(n24), .B0(SH[15]), .Y(n22) );
  OR4X1 U50 ( .A(n25), .B(SH[10]), .C(SH[11]), .D(SH[12]), .Y(n24) );
  OR2X1 U51 ( .A(SH[14]), .B(SH[13]), .Y(n25) );
  NAND4X1 U52 ( .A(n14), .B(n13), .C(n26), .D(n12), .Y(n23) );
  NOR2X1 U53 ( .A(SH[9]), .B(SH[8]), .Y(n26) );
  NAND2X1 U54 ( .A(SH[15]), .B(n27), .Y(n21) );
  NAND4BXL U55 ( .AN(n28), .B(SH[9]), .C(SH[8]), .D(n29), .Y(n27) );
  NOR3X1 U56 ( .A(n12), .B(n14), .C(n13), .Y(n29) );
  NAND3BX1 U57 ( .AN(n30), .B(SH[13]), .C(SH[14]), .Y(n28) );
  NAND3X1 U58 ( .A(SH[11]), .B(SH[10]), .C(SH[12]), .Y(n30) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [16:0] carry;

  ADDFX2 U2_14 ( .A(A[14]), .B(n2), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFX2 U2_13 ( .A(A[13]), .B(n3), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFX2 U2_12 ( .A(A[12]), .B(n4), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFX2 U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFX2 U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFX2 U2_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFX2 U2_8 ( .A(A[8]), .B(n8), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFX2 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  XOR3X2 U2_15 ( .A(A[15]), .B(n1), .C(carry[15]), .Y(DIFF[15]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFX2 U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFX2 U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFX2 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  INVX1 U1 ( .A(B[0]), .Y(n16) );
  INVX1 U2 ( .A(B[2]), .Y(n14) );
  INVX1 U3 ( .A(B[3]), .Y(n13) );
  INVX1 U4 ( .A(B[4]), .Y(n12) );
  INVX1 U5 ( .A(B[1]), .Y(n15) );
  OR2X2 U6 ( .A(A[0]), .B(n16), .Y(carry[1]) );
  INVX1 U7 ( .A(B[15]), .Y(n1) );
  INVX1 U8 ( .A(B[5]), .Y(n11) );
  INVX1 U9 ( .A(B[6]), .Y(n10) );
  INVX1 U10 ( .A(B[7]), .Y(n9) );
  INVX1 U11 ( .A(B[8]), .Y(n8) );
  INVX1 U12 ( .A(B[9]), .Y(n7) );
  INVX1 U13 ( .A(B[10]), .Y(n6) );
  INVX1 U14 ( .A(B[11]), .Y(n5) );
  INVX1 U15 ( .A(B[12]), .Y(n4) );
  INVX1 U16 ( .A(B[13]), .Y(n3) );
  INVX1 U17 ( .A(B[14]), .Y(n2) );
  XNOR2X1 U18 ( .A(n16), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;

  wire   [15:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  XOR3X2 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu ( a, b, cmd, r );
  input [15:0] a;
  input [15:0] b;
  input [2:0] cmd;
  output [15:0] r;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n29, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n61, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249;

  alu_DW_rash_0 srl_40 ( .A({n35, n34, n33, n29, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, a[0]}), .DATA_TC(1'b0), .SH({b[15:5], n16, 
        n15, n14, n13, n12}), .SH_TC(1'b0), .B({N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147}) );
  alu_DW01_ash_0 sll_36 ( .A({n35, n34, n33, n29, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, a[0]}), .DATA_TC(1'b0), .SH({b[15:5], n16, 
        n15, n14, n13, n12}), .SH_TC(1'b0), .B({N130, N129, N128, N127, N126, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115}) );
  alu_DW01_sub_0 sub_28 ( .A({n35, n34, n33, n29, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, a[0]}), .B({b[15:5], n16, n15, n14, n13, n12}), .CI(1'b0), .DIFF({N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51}) );
  alu_DW01_add_0 add_26 ( .A({n35, n34, n33, n29, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, a[0]}), .B({b[15:5], n16, n15, n14, n13, n12}), .CI(1'b0), .SUM({N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35}) );
  OAI221XL U3 ( .A0(n5), .A1(n191), .B0(n193), .B1(n2), .C0(n140), .Y(n165) );
  OAI221XL U4 ( .A0(n5), .A1(n187), .B0(n189), .B1(n2), .C0(n45), .Y(n160) );
  AOI222X1 U5 ( .A0(n1), .A1(n33), .B0(n4), .B1(n34), .C0(n13), .C1(n35), .Y(
        n244) );
  OAI221XL U6 ( .A0(n5), .A1(n180), .B0(n2), .B1(n181), .C0(n43), .Y(n44) );
  AOI222X1 U7 ( .A0(N41), .A1(n55), .B0(N121), .B1(n56), .C0(N57), .C1(n57), 
        .Y(n77) );
  AOI222X1 U8 ( .A0(N42), .A1(n55), .B0(N122), .B1(n56), .C0(N58), .C1(n57), 
        .Y(n72) );
  AOI222X1 U12 ( .A0(N46), .A1(n55), .B0(N126), .B1(n56), .C0(N62), .C1(n57), 
        .Y(n127) );
  AOI222X1 U13 ( .A0(N49), .A1(n55), .B0(N129), .B1(n56), .C0(N65), .C1(n57), 
        .Y(n112) );
  AOI222X1 U14 ( .A0(N47), .A1(n55), .B0(N127), .B1(n56), .C0(N63), .C1(n57), 
        .Y(n122) );
  AOI222X1 U15 ( .A0(N48), .A1(n55), .B0(N128), .B1(n56), .C0(N64), .C1(n57), 
        .Y(n117) );
  AOI222X1 U16 ( .A0(N39), .A1(n55), .B0(N119), .B1(n56), .C0(N55), .C1(n57), 
        .Y(n87) );
  AOI222X1 U17 ( .A0(N40), .A1(n55), .B0(N120), .B1(n56), .C0(N56), .C1(n57), 
        .Y(n82) );
  AOI222X1 U18 ( .A0(N43), .A1(n55), .B0(N123), .B1(n56), .C0(N59), .C1(n57), 
        .Y(n67) );
  AOI222X1 U19 ( .A0(N37), .A1(n55), .B0(N117), .B1(n56), .C0(N53), .C1(n57), 
        .Y(n97) );
  AOI222X1 U20 ( .A0(N38), .A1(n55), .B0(N118), .B1(n56), .C0(N54), .C1(n57), 
        .Y(n92) );
  AOI222X1 U21 ( .A0(N36), .A1(n55), .B0(N116), .B1(n56), .C0(N52), .C1(n57), 
        .Y(n102) );
  NOR2X4 U22 ( .A(n12), .B(n13), .Y(n1) );
  NAND2X2 U23 ( .A(n12), .B(n13), .Y(n2) );
  NAND2X4 U24 ( .A(cmd[1]), .B(n245), .Y(n3) );
  NOR2X4 U25 ( .A(n168), .B(n13), .Y(n4) );
  NAND2X2 U26 ( .A(n168), .B(n13), .Y(n5) );
  NAND4X2 U27 ( .A(n51), .B(n50), .C(n49), .D(n48), .Y(n162) );
  CLKINVX3 U28 ( .A(n7), .Y(n64) );
  CLKINVX3 U29 ( .A(n10), .Y(n57) );
  CLKINVX3 U30 ( .A(n9), .Y(n56) );
  CLKINVX3 U31 ( .A(n8), .Y(n55) );
  OAI221XL U32 ( .A0(n5), .A1(n189), .B0(n2), .B1(n191), .C0(n145), .Y(n161)
         );
  OAI221XL U33 ( .A0(n5), .A1(n181), .B0(n2), .B1(n183), .C0(n146), .Y(n147)
         );
  OAI221XL U34 ( .A0(n195), .A1(n5), .B0(n206), .B1(n2), .C0(n42), .Y(n207) );
  CLKINVX3 U35 ( .A(n6), .Y(n63) );
  AOI2BB1XL U36 ( .A0N(n175), .A1N(n234), .B0(n242), .Y(n209) );
  OAI32XL U37 ( .A0(n164), .A1(n203), .A2(n163), .B0(n162), .B1(n233), .Y(n228) );
  OAI32XL U38 ( .A0(n230), .A1(n172), .A2(n162), .B0(n244), .B1(n163), .Y(n231) );
  OAI33XL U39 ( .A0(n164), .A1(n234), .A2(n163), .B0(n233), .B1(n13), .B2(n162), .Y(n235) );
  AOI22XL U40 ( .A0(n25), .A1(n4), .B0(n24), .B1(n1), .Y(n45) );
  AOI22XL U41 ( .A0(n33), .A1(n4), .B0(n29), .B1(n1), .Y(n42) );
  AOI22XL U42 ( .A0(n26), .A1(n4), .B0(n25), .B1(n1), .Y(n145) );
  NOR2XL U43 ( .A(n61), .B(n162), .Y(N131) );
  AOI21XL U44 ( .A0(n223), .A1(n222), .B0(n162), .Y(N133) );
  AOI31XL U45 ( .A0(n233), .A1(n219), .A2(n218), .B0(n162), .Y(N132) );
  AOI22XL U46 ( .A0(n27), .A1(n4), .B0(n26), .B1(n1), .Y(n140) );
  AOI22XL U47 ( .A0(n22), .A1(n4), .B0(n21), .B1(n1), .Y(n146) );
  AOI22XL U48 ( .A0(n29), .A1(n4), .B0(n27), .B1(n1), .Y(n141) );
  AOI22XL U49 ( .A0(n23), .A1(n4), .B0(n22), .B1(n1), .Y(n151) );
  AOI22XL U50 ( .A0(n24), .A1(n4), .B0(n23), .B1(n1), .Y(n156) );
  AOI22XL U51 ( .A0(n21), .A1(n4), .B0(n20), .B1(n1), .Y(n43) );
  AOI21XL U52 ( .A0(n227), .A1(n226), .B0(n162), .Y(N134) );
  AOI21XL U53 ( .A0(n35), .A1(n1), .B0(n202), .Y(n224) );
  AOI22XL U54 ( .A0(n18), .A1(n4), .B0(n17), .B1(n1), .Y(n144) );
  AOI22XL U55 ( .A0(n19), .A1(n4), .B0(n18), .B1(n1), .Y(n149) );
  AOI22XL U56 ( .A0(n20), .A1(n4), .B0(n19), .B1(n1), .Y(n153) );
  NAND2XL U57 ( .A(n35), .B(n2), .Y(n230) );
  AOI22XL U58 ( .A0(n17), .A1(n4), .B0(a[0]), .B1(n1), .Y(n46) );
  INVX1 U59 ( .A(n211), .Y(n205) );
  INVX1 U60 ( .A(n166), .Y(n175) );
  INVX1 U61 ( .A(n219), .Y(n204) );
  INVX1 U62 ( .A(n220), .Y(n200) );
  INVX1 U63 ( .A(n241), .Y(n201) );
  INVX1 U64 ( .A(n143), .Y(n174) );
  BUFX3 U65 ( .A(n167), .Y(n11) );
  NAND3BX1 U66 ( .AN(n163), .B(n169), .C(n170), .Y(n167) );
  INVX1 U67 ( .A(n161), .Y(n192) );
  INVX1 U68 ( .A(n164), .Y(n171) );
  INVX1 U69 ( .A(n165), .Y(n194) );
  INVX1 U70 ( .A(n160), .Y(n190) );
  INVX1 U71 ( .A(n230), .Y(n198) );
  INVX1 U72 ( .A(n210), .Y(n202) );
  INVX1 U73 ( .A(n224), .Y(n199) );
  CLKINVX3 U74 ( .A(n41), .Y(n39) );
  CLKINVX3 U75 ( .A(n38), .Y(n36) );
  INVX1 U76 ( .A(n38), .Y(n37) );
  INVX1 U77 ( .A(n41), .Y(n40) );
  INVX1 U78 ( .A(n238), .Y(n197) );
  INVX1 U79 ( .A(n162), .Y(n173) );
  NAND3X1 U80 ( .A(n85), .B(n86), .C(n87), .Y(r[4]) );
  AOI22X1 U81 ( .A0(n20), .A1(n88), .B0(n16), .B1(n89), .Y(n86) );
  AOI22XL U82 ( .A0(N151), .A1(n63), .B0(N135), .B1(n64), .Y(n85) );
  INVX1 U83 ( .A(n16), .Y(n172) );
  NAND3X1 U84 ( .A(n100), .B(n101), .C(n102), .Y(r[1]) );
  AOI22X1 U85 ( .A0(n17), .A1(n103), .B0(n13), .B1(n104), .Y(n101) );
  AOI22XL U86 ( .A0(N148), .A1(n63), .B0(N132), .B1(n64), .Y(n100) );
  NAND3X1 U87 ( .A(n95), .B(n96), .C(n97), .Y(r[2]) );
  AOI22X1 U88 ( .A0(n18), .A1(n98), .B0(n14), .B1(n99), .Y(n96) );
  AOI22XL U89 ( .A0(N149), .A1(n63), .B0(N133), .B1(n64), .Y(n95) );
  NAND3X1 U90 ( .A(n90), .B(n91), .C(n92), .Y(r[3]) );
  AOI22X1 U91 ( .A0(n19), .A1(n93), .B0(n15), .B1(n94), .Y(n91) );
  AOI22XL U92 ( .A0(N150), .A1(n63), .B0(N134), .B1(n64), .Y(n90) );
  INVX1 U93 ( .A(n35), .Y(n206) );
  INVX1 U94 ( .A(n15), .Y(n170) );
  INVX1 U95 ( .A(n14), .Y(n169) );
  INVX1 U96 ( .A(n12), .Y(n168) );
  INVX1 U97 ( .A(n27), .Y(n189) );
  INVX1 U98 ( .A(n29), .Y(n191) );
  INVX1 U99 ( .A(n147), .Y(n184) );
  INVX1 U100 ( .A(n157), .Y(n188) );
  INVX1 U101 ( .A(n142), .Y(n196) );
  INVX1 U102 ( .A(n207), .Y(n203) );
  INVX1 U103 ( .A(n44), .Y(n182) );
  INVX1 U104 ( .A(n152), .Y(n186) );
  INVX1 U105 ( .A(n33), .Y(n193) );
  INVX1 U106 ( .A(n34), .Y(n195) );
  INVX1 U107 ( .A(n24), .Y(n183) );
  INVX1 U108 ( .A(n23), .Y(n181) );
  INVX1 U109 ( .A(n26), .Y(n187) );
  INVX1 U110 ( .A(n25), .Y(n185) );
  INVX1 U111 ( .A(n22), .Y(n180) );
  OAI221XL U112 ( .A0(n25), .A1(n39), .B0(n185), .B1(n3), .C0(n36), .Y(n59) );
  OAI221XL U113 ( .A0(n17), .A1(n39), .B0(n3), .B1(n248), .C0(n36), .Y(n104)
         );
  INVX1 U114 ( .A(n17), .Y(n248) );
  OAI221XL U115 ( .A0(n18), .A1(n39), .B0(n3), .B1(n176), .C0(n36), .Y(n99) );
  OAI221XL U116 ( .A0(n19), .A1(n39), .B0(n3), .B1(n177), .C0(n36), .Y(n94) );
  OAI221XL U117 ( .A0(n20), .A1(n39), .B0(n3), .B1(n178), .C0(n36), .Y(n89) );
  OAI221XL U118 ( .A0(n21), .A1(n39), .B0(n3), .B1(n179), .C0(n36), .Y(n84) );
  OAI221XL U119 ( .A0(n22), .A1(n39), .B0(n3), .B1(n180), .C0(n36), .Y(n79) );
  OAI221XL U120 ( .A0(n23), .A1(n39), .B0(n3), .B1(n181), .C0(n36), .Y(n74) );
  OAI221XL U121 ( .A0(n24), .A1(n39), .B0(n3), .B1(n183), .C0(n36), .Y(n69) );
  OAI221XL U122 ( .A0(n26), .A1(n40), .B0(n3), .B1(n187), .C0(n37), .Y(n134)
         );
  OAI221XL U123 ( .A0(n27), .A1(n40), .B0(n3), .B1(n189), .C0(n37), .Y(n129)
         );
  OAI221XL U124 ( .A0(n29), .A1(n40), .B0(n3), .B1(n191), .C0(n37), .Y(n124)
         );
  OAI221XL U125 ( .A0(n33), .A1(n40), .B0(n3), .B1(n193), .C0(n37), .Y(n119)
         );
  OAI221XL U126 ( .A0(n34), .A1(n40), .B0(n3), .B1(n195), .C0(n37), .Y(n114)
         );
  OAI221XL U127 ( .A0(n35), .A1(n39), .B0(n3), .B1(n206), .C0(n37), .Y(n109)
         );
  OAI21XL U128 ( .A0(n13), .A1(n39), .B0(n36), .Y(n103) );
  OAI21XL U129 ( .A0(n12), .A1(n39), .B0(n36), .Y(n138) );
  OAI21XL U130 ( .A0(n14), .A1(n39), .B0(n36), .Y(n98) );
  OAI21XL U131 ( .A0(n15), .A1(n39), .B0(n36), .Y(n93) );
  OAI21XL U132 ( .A0(n16), .A1(n39), .B0(n36), .Y(n88) );
  INVX1 U133 ( .A(n19), .Y(n177) );
  INVX1 U134 ( .A(n20), .Y(n178) );
  INVX1 U135 ( .A(n21), .Y(n179) );
  INVX1 U136 ( .A(n18), .Y(n176) );
  INVX1 U137 ( .A(n60), .Y(n41) );
  INVX1 U138 ( .A(n62), .Y(n38) );
  OR3XL U139 ( .A(n247), .B(n245), .C(n246), .Y(n6) );
  NAND3X1 U140 ( .A(n110), .B(n111), .C(n112), .Y(r[14]) );
  AOI22X1 U141 ( .A0(n34), .A1(n113), .B0(b[14]), .B1(n114), .Y(n111) );
  AOI22XL U142 ( .A0(N161), .A1(n63), .B0(N145), .B1(n64), .Y(n110) );
  NAND3X1 U143 ( .A(n125), .B(n126), .C(n127), .Y(r[11]) );
  AOI22X1 U144 ( .A0(n27), .A1(n128), .B0(b[11]), .B1(n129), .Y(n126) );
  AOI22XL U145 ( .A0(N158), .A1(n63), .B0(N142), .B1(n64), .Y(n125) );
  NAND3X1 U146 ( .A(n75), .B(n76), .C(n77), .Y(r[6]) );
  AOI22X1 U147 ( .A0(n22), .A1(n78), .B0(b[6]), .B1(n79), .Y(n76) );
  AOI22XL U148 ( .A0(N153), .A1(n63), .B0(N137), .B1(n64), .Y(n75) );
  NAND3X1 U149 ( .A(n80), .B(n81), .C(n82), .Y(r[5]) );
  AOI22X1 U150 ( .A0(n21), .A1(n83), .B0(b[5]), .B1(n84), .Y(n81) );
  AOI22XL U151 ( .A0(N152), .A1(n63), .B0(N136), .B1(n64), .Y(n80) );
  NAND3X1 U152 ( .A(n70), .B(n71), .C(n72), .Y(r[7]) );
  AOI22X1 U153 ( .A0(n23), .A1(n73), .B0(b[7]), .B1(n74), .Y(n71) );
  AOI22XL U154 ( .A0(N154), .A1(n63), .B0(N138), .B1(n64), .Y(n70) );
  NAND3X1 U155 ( .A(n65), .B(n66), .C(n67), .Y(r[8]) );
  AOI22X1 U156 ( .A0(n24), .A1(n68), .B0(b[8]), .B1(n69), .Y(n66) );
  AOI22XL U157 ( .A0(N155), .A1(n63), .B0(N139), .B1(n64), .Y(n65) );
  NAND3X1 U158 ( .A(n120), .B(n121), .C(n122), .Y(r[12]) );
  AOI22X1 U159 ( .A0(n29), .A1(n123), .B0(b[12]), .B1(n124), .Y(n121) );
  AOI22XL U160 ( .A0(N159), .A1(n63), .B0(N143), .B1(n64), .Y(n120) );
  NAND3X1 U161 ( .A(n115), .B(n116), .C(n117), .Y(r[13]) );
  AOI22X1 U162 ( .A0(n33), .A1(n118), .B0(b[13]), .B1(n119), .Y(n116) );
  AOI22XL U163 ( .A0(N160), .A1(n63), .B0(N144), .B1(n64), .Y(n115) );
  NAND3X1 U164 ( .A(n52), .B(n53), .C(n54), .Y(r[9]) );
  AOI22X1 U165 ( .A0(n25), .A1(n58), .B0(b[9]), .B1(n59), .Y(n53) );
  AOI222XL U166 ( .A0(N44), .A1(n55), .B0(N124), .B1(n56), .C0(N60), .C1(n57), 
        .Y(n54) );
  AOI22XL U167 ( .A0(N156), .A1(n63), .B0(N140), .B1(n64), .Y(n52) );
  NAND3X1 U168 ( .A(n130), .B(n131), .C(n132), .Y(r[10]) );
  AOI22X1 U169 ( .A0(n26), .A1(n133), .B0(b[10]), .B1(n134), .Y(n131) );
  AOI222XL U170 ( .A0(N45), .A1(n55), .B0(N125), .B1(n56), .C0(N61), .C1(n57), 
        .Y(n132) );
  AOI22XL U171 ( .A0(N157), .A1(n63), .B0(N141), .B1(n64), .Y(n130) );
  NAND3X1 U172 ( .A(n135), .B(n136), .C(n137), .Y(r[0]) );
  AOI22X1 U173 ( .A0(a[0]), .A1(n138), .B0(n12), .B1(n139), .Y(n136) );
  AOI22XL U174 ( .A0(N147), .A1(n63), .B0(N131), .B1(n64), .Y(n135) );
  AOI222XL U175 ( .A0(N35), .A1(n55), .B0(N115), .B1(n56), .C0(N51), .C1(n57), 
        .Y(n137) );
  NAND3X1 U176 ( .A(n105), .B(n106), .C(n107), .Y(r[15]) );
  AOI22X1 U177 ( .A0(n35), .A1(n108), .B0(b[15]), .B1(n109), .Y(n106) );
  AOI222XL U178 ( .A0(N50), .A1(n55), .B0(N130), .B1(n56), .C0(N66), .C1(n57), 
        .Y(n107) );
  AOI22XL U179 ( .A0(N162), .A1(n63), .B0(N146), .B1(n64), .Y(n105) );
  BUFX3 U180 ( .A(b[4]), .Y(n16) );
  BUFX3 U181 ( .A(a[15]), .Y(n35) );
  BUFX3 U182 ( .A(b[1]), .Y(n13) );
  BUFX3 U183 ( .A(b[2]), .Y(n14) );
  BUFX3 U184 ( .A(a[13]), .Y(n33) );
  BUFX3 U185 ( .A(a[14]), .Y(n34) );
  BUFX3 U186 ( .A(a[11]), .Y(n27) );
  BUFX3 U187 ( .A(a[12]), .Y(n29) );
  BUFX3 U188 ( .A(b[0]), .Y(n12) );
  BUFX3 U189 ( .A(b[3]), .Y(n15) );
  BUFX3 U190 ( .A(a[1]), .Y(n17) );
  BUFX3 U191 ( .A(a[7]), .Y(n23) );
  BUFX3 U192 ( .A(a[8]), .Y(n24) );
  BUFX3 U193 ( .A(a[9]), .Y(n25) );
  BUFX3 U194 ( .A(a[10]), .Y(n26) );
  BUFX3 U195 ( .A(a[6]), .Y(n22) );
  BUFX3 U196 ( .A(a[3]), .Y(n19) );
  BUFX3 U197 ( .A(a[4]), .Y(n20) );
  BUFX3 U198 ( .A(a[2]), .Y(n18) );
  BUFX3 U199 ( .A(a[5]), .Y(n21) );
  OAI221XL U200 ( .A0(a[0]), .A1(n39), .B0(n3), .B1(n249), .C0(n36), .Y(n139)
         );
  INVX1 U201 ( .A(a[0]), .Y(n249) );
  INVX1 U202 ( .A(cmd[2]), .Y(n245) );
  INVX1 U203 ( .A(cmd[1]), .Y(n246) );
  NAND3X1 U204 ( .A(cmd[0]), .B(n245), .C(cmd[1]), .Y(n62) );
  NAND3X1 U205 ( .A(n247), .B(n246), .C(cmd[2]), .Y(n60) );
  INVX1 U206 ( .A(cmd[0]), .Y(n247) );
  OAI21XL U207 ( .A0(b[15]), .A1(n39), .B0(n36), .Y(n108) );
  OAI21XL U208 ( .A0(b[12]), .A1(n60), .B0(n36), .Y(n123) );
  OAI21XL U209 ( .A0(b[9]), .A1(n60), .B0(n62), .Y(n58) );
  OAI21XL U210 ( .A0(b[11]), .A1(n60), .B0(n62), .Y(n128) );
  OAI21XL U211 ( .A0(b[8]), .A1(n60), .B0(n62), .Y(n68) );
  OAI21XL U212 ( .A0(b[14]), .A1(n60), .B0(n62), .Y(n113) );
  OAI21XL U213 ( .A0(b[13]), .A1(n40), .B0(n62), .Y(n118) );
  OAI21XL U214 ( .A0(b[10]), .A1(n60), .B0(n62), .Y(n133) );
  OAI21XL U215 ( .A0(b[7]), .A1(n39), .B0(n36), .Y(n73) );
  OAI21XL U216 ( .A0(b[6]), .A1(n39), .B0(n36), .Y(n78) );
  OAI21XL U217 ( .A0(b[5]), .A1(n39), .B0(n36), .Y(n83) );
  OR3XL U218 ( .A(n245), .B(cmd[0]), .C(n246), .Y(n7) );
  OR3XL U219 ( .A(cmd[1]), .B(cmd[2]), .C(cmd[0]), .Y(n8) );
  OR3XL U220 ( .A(n245), .B(cmd[1]), .C(n247), .Y(n9) );
  OR3XL U221 ( .A(cmd[1]), .B(cmd[2]), .C(n247), .Y(n10) );
  NAND2X1 U222 ( .A(n15), .B(n14), .Y(n159) );
  NAND2X1 U223 ( .A(n170), .B(n14), .Y(n158) );
  NAND2X1 U224 ( .A(n15), .B(n169), .Y(n164) );
  NOR3X1 U225 ( .A(n14), .B(n16), .C(n15), .Y(n155) );
  OAI221XL U226 ( .A0(n5), .A1(n176), .B0(n2), .B1(n177), .C0(n46), .Y(n47) );
  NOR2X1 U227 ( .A(b[11]), .B(b[10]), .Y(n51) );
  NOR3X1 U228 ( .A(b[12]), .B(b[14]), .C(b[13]), .Y(n50) );
  NOR3X1 U229 ( .A(b[15]), .B(b[6]), .C(b[5]), .Y(n49) );
  NOR3X1 U230 ( .A(b[7]), .B(b[9]), .C(b[8]), .Y(n48) );
  NAND2X1 U231 ( .A(n173), .B(n172), .Y(n163) );
  NAND3X1 U232 ( .A(n16), .B(n170), .C(n173), .Y(n143) );
  NOR2X1 U233 ( .A(n158), .B(n163), .Y(n166) );
  OAI221XL U234 ( .A0(n193), .A1(n5), .B0(n195), .B1(n2), .C0(n141), .Y(n142)
         );
  OAI221XL U235 ( .A0(n5), .A1(n177), .B0(n2), .B1(n178), .C0(n144), .Y(n148)
         );
  OAI221XL U236 ( .A0(n5), .A1(n178), .B0(n2), .B1(n179), .C0(n149), .Y(n150)
         );
  OAI221XL U237 ( .A0(n5), .A1(n183), .B0(n2), .B1(n185), .C0(n151), .Y(n152)
         );
  OAI221XL U238 ( .A0(n5), .A1(n179), .B0(n2), .B1(n180), .C0(n153), .Y(n154)
         );
  OAI221XL U239 ( .A0(n5), .A1(n185), .B0(n2), .B1(n187), .C0(n156), .Y(n157)
         );
  NAND2X1 U240 ( .A(n205), .B(n214), .Y(N146) );
  NAND4X1 U241 ( .A(n1), .B(n202), .C(n173), .D(n170), .Y(n214) );
  OAI221XL U242 ( .A0(n13), .A1(n241), .B0(n234), .B1(n11), .C0(n213), .Y(N145) );
  OAI221XL U243 ( .A0(n196), .A1(n11), .B0(n224), .B1(n143), .C0(n213), .Y(
        N142) );
  OAI221XL U244 ( .A0(n244), .A1(n175), .B0(n192), .B1(n11), .C0(n243), .Y(
        N140) );
  OAI211X1 U245 ( .A0(n184), .A1(n11), .B0(n237), .C0(n232), .Y(N136) );
  AOI22X1 U246 ( .A0(n171), .A1(n231), .B0(n166), .B1(n161), .Y(n232) );
  OAI211X1 U247 ( .A0(n244), .A1(n11), .B0(n212), .C0(n213), .Y(N144) );
  NAND3X1 U248 ( .A(n174), .B(n169), .C(n198), .Y(n212) );
  AOI211X1 U249 ( .A0(n198), .A1(n174), .B0(n242), .C0(n201), .Y(n243) );
  OAI211X1 U250 ( .A0(n196), .A1(n175), .B0(n239), .C0(n197), .Y(N138) );
  OAI21XL U251 ( .A0(n11), .A1(n188), .B0(n240), .Y(n238) );
  NAND4X1 U252 ( .A(n171), .B(n1), .C(n35), .D(n173), .Y(n239) );
  AOI221X1 U253 ( .A0(n208), .A1(n172), .B0(n155), .B1(n47), .C0(n215), .Y(n61) );
  OAI222XL U254 ( .A0(n203), .A1(n159), .B0(n182), .B1(n158), .C0(n190), .C1(
        n164), .Y(n208) );
  OAI211X1 U255 ( .A0(n203), .A1(n11), .B0(n241), .C0(n213), .Y(N143) );
  NAND2X1 U256 ( .A(n174), .B(n202), .Y(n241) );
  OAI221XL U257 ( .A0(n203), .A1(n175), .B0(n190), .B1(n11), .C0(n240), .Y(
        N139) );
  AOI21X1 U258 ( .A0(n35), .A1(n174), .B0(n242), .Y(n240) );
  AOI21X1 U259 ( .A0(n155), .A1(n148), .B0(n217), .Y(n218) );
  MX2X1 U260 ( .A(n198), .B(n216), .S0(n172), .Y(n217) );
  OAI222XL U261 ( .A0(n164), .A1(n192), .B0(n158), .B1(n184), .C0(n159), .C1(
        n244), .Y(n216) );
  MXI2X1 U262 ( .A(n221), .B(n220), .S0(n16), .Y(n222) );
  OAI222XL U263 ( .A0(n234), .A1(n159), .B0(n186), .B1(n158), .C0(n194), .C1(
        n164), .Y(n221) );
  AOI21X1 U264 ( .A0(n155), .A1(n150), .B0(n204), .Y(n223) );
  MXI2X1 U265 ( .A(n225), .B(n199), .S0(n16), .Y(n226) );
  OAI222XL U266 ( .A0(n206), .A1(n159), .B0(n188), .B1(n158), .C0(n196), .C1(
        n164), .Y(n225) );
  AOI21X1 U267 ( .A0(n155), .A1(n154), .B0(n204), .Y(n227) );
  NAND2X1 U268 ( .A(n215), .B(n170), .Y(n219) );
  OAI211X1 U269 ( .A0(n186), .A1(n11), .B0(n237), .C0(n236), .Y(N137) );
  AOI21X1 U270 ( .A0(n166), .A1(n165), .B0(n235), .Y(n236) );
  OAI211X1 U271 ( .A0(n182), .A1(n11), .B0(n237), .C0(n229), .Y(N135) );
  AOI21X1 U272 ( .A0(n166), .A1(n160), .B0(n228), .Y(n229) );
  NAND2X1 U273 ( .A(n215), .B(n169), .Y(n233) );
  NOR2X1 U274 ( .A(n206), .B(n172), .Y(n215) );
  AOI22X1 U275 ( .A0(n35), .A1(n174), .B0(n14), .B1(n242), .Y(n237) );
  OAI221XL U276 ( .A0(n194), .A1(n11), .B0(n200), .B1(n143), .C0(n209), .Y(
        N141) );
  MXI2X1 U277 ( .A(n35), .B(n34), .S0(n1), .Y(n234) );
  OAI21XL U278 ( .A0(n13), .A1(n206), .B0(n210), .Y(n220) );
  NAND2X1 U279 ( .A(n35), .B(n169), .Y(n210) );
  AOI21X1 U280 ( .A0(n14), .A1(n211), .B0(n242), .Y(n213) );
  NOR2X1 U281 ( .A(n205), .B(n170), .Y(n242) );
  NOR2X1 U282 ( .A(n206), .B(n163), .Y(n211) );
endmodule


module EX_stage ( clk, rst, pipeline_reg_in, pipeline_reg_out, ex_op_dest );
  input [56:0] pipeline_reg_in;
  output [37:0] pipeline_reg_out;
  output [2:0] ex_op_dest;
  input clk, rst;
  wire   pipeline_reg_in_0, \pipeline_reg_in[3] , \pipeline_reg_in[2] ,
         \pipeline_reg_in[1] , n39;
  wire   [15:0] ex_alu_result;
  assign pipeline_reg_in_0 = pipeline_reg_in[0];
  assign ex_op_dest[2] = \pipeline_reg_in[3] ;
  assign \pipeline_reg_in[3]  = pipeline_reg_in[3];
  assign ex_op_dest[1] = \pipeline_reg_in[2] ;
  assign \pipeline_reg_in[2]  = pipeline_reg_in[2];
  assign ex_op_dest[0] = \pipeline_reg_in[1] ;
  assign \pipeline_reg_in[1]  = pipeline_reg_in[1];

  alu alu_inst ( .a(pipeline_reg_in[53:38]), .b(pipeline_reg_in[37:22]), .cmd(
        pipeline_reg_in[56:54]), .r(ex_alu_result) );
  DFFTRXL \pipeline_reg_out_reg[1]  ( .D(\pipeline_reg_in[1] ), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[1]) );
  DFFTRXL \pipeline_reg_out_reg[0]  ( .D(pipeline_reg_in_0), .RN(n39), .CK(clk), .Q(pipeline_reg_out[0]) );
  DFFTRXL \pipeline_reg_out_reg[13]  ( .D(pipeline_reg_in[13]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[13]) );
  DFFTRXL \pipeline_reg_out_reg[12]  ( .D(pipeline_reg_in[12]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[12]) );
  DFFTRXL \pipeline_reg_out_reg[11]  ( .D(pipeline_reg_in[11]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[11]) );
  DFFTRXL \pipeline_reg_out_reg[10]  ( .D(pipeline_reg_in[10]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[10]) );
  DFFTRXL \pipeline_reg_out_reg[9]  ( .D(pipeline_reg_in[9]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[9]) );
  DFFTRXL \pipeline_reg_out_reg[8]  ( .D(pipeline_reg_in[8]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[8]) );
  DFFTRXL \pipeline_reg_out_reg[7]  ( .D(pipeline_reg_in[7]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[7]) );
  DFFTRXL \pipeline_reg_out_reg[6]  ( .D(pipeline_reg_in[6]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[6]) );
  DFFTRXL \pipeline_reg_out_reg[5]  ( .D(pipeline_reg_in[5]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[5]) );
  DFFTRXL \pipeline_reg_out_reg[4]  ( .D(pipeline_reg_in[4]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[4]) );
  DFFTRXL \pipeline_reg_out_reg[3]  ( .D(\pipeline_reg_in[3] ), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[3]) );
  DFFTRXL \pipeline_reg_out_reg[2]  ( .D(\pipeline_reg_in[2] ), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[2]) );
  DFFTRXL \pipeline_reg_out_reg[21]  ( .D(pipeline_reg_in[21]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[21]) );
  DFFTRXL \pipeline_reg_out_reg[20]  ( .D(pipeline_reg_in[20]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[20]) );
  DFFTRXL \pipeline_reg_out_reg[19]  ( .D(pipeline_reg_in[19]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[19]) );
  DFFTRXL \pipeline_reg_out_reg[18]  ( .D(pipeline_reg_in[18]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[18]) );
  DFFTRXL \pipeline_reg_out_reg[17]  ( .D(pipeline_reg_in[17]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[17]) );
  DFFTRXL \pipeline_reg_out_reg[16]  ( .D(pipeline_reg_in[16]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[16]) );
  DFFTRXL \pipeline_reg_out_reg[15]  ( .D(pipeline_reg_in[15]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[15]) );
  DFFTRXL \pipeline_reg_out_reg[14]  ( .D(pipeline_reg_in[14]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[14]) );
  DFFTRXL \pipeline_reg_out_reg[22]  ( .D(ex_alu_result[0]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[22]) );
  DFFTRXL \pipeline_reg_out_reg[23]  ( .D(ex_alu_result[1]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[23]) );
  DFFTRXL \pipeline_reg_out_reg[25]  ( .D(ex_alu_result[3]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[25]) );
  DFFTRXL \pipeline_reg_out_reg[24]  ( .D(ex_alu_result[2]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[24]) );
  DFFTRXL \pipeline_reg_out_reg[37]  ( .D(ex_alu_result[15]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[37]) );
  DFFTRXL \pipeline_reg_out_reg[31]  ( .D(ex_alu_result[9]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[31]) );
  DFFTRXL \pipeline_reg_out_reg[32]  ( .D(ex_alu_result[10]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[32]) );
  DFFTRXL \pipeline_reg_out_reg[30]  ( .D(ex_alu_result[8]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[30]) );
  DFFTRXL \pipeline_reg_out_reg[27]  ( .D(ex_alu_result[5]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[27]) );
  DFFTRXL \pipeline_reg_out_reg[26]  ( .D(ex_alu_result[4]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[26]) );
  DFFTRXL \pipeline_reg_out_reg[35]  ( .D(ex_alu_result[13]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[35]) );
  DFFTRXL \pipeline_reg_out_reg[34]  ( .D(ex_alu_result[12]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[34]) );
  DFFTRXL \pipeline_reg_out_reg[36]  ( .D(ex_alu_result[14]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[36]) );
  DFFTRXL \pipeline_reg_out_reg[33]  ( .D(ex_alu_result[11]), .RN(n39), .CK(
        clk), .Q(pipeline_reg_out[33]) );
  DFFTRX4 \pipeline_reg_out_reg[29]  ( .D(ex_alu_result[7]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[29]) );
  DFFTRX4 \pipeline_reg_out_reg[28]  ( .D(ex_alu_result[6]), .RN(n39), .CK(clk), .Q(pipeline_reg_out[28]) );
  INVX8 U3 ( .A(rst), .Y(n39) );
endmodule


module data_mem ( clk, mem_access_addr, mem_write_data, mem_write_en, 
        mem_read_data );
  input [15:0] mem_access_addr;
  input [15:0] mem_write_data;
  output [15:0] mem_read_data;
  input clk, mem_write_en;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \ram[255][15] ,
         \ram[255][14] , \ram[255][13] , \ram[255][12] , \ram[255][11] ,
         \ram[255][10] , \ram[255][9] , \ram[255][8] , \ram[255][7] ,
         \ram[255][6] , \ram[255][5] , \ram[255][4] , \ram[255][3] ,
         \ram[255][2] , \ram[255][1] , \ram[255][0] , \ram[254][15] ,
         \ram[254][14] , \ram[254][13] , \ram[254][12] , \ram[254][11] ,
         \ram[254][10] , \ram[254][9] , \ram[254][8] , \ram[254][7] ,
         \ram[254][6] , \ram[254][5] , \ram[254][4] , \ram[254][3] ,
         \ram[254][2] , \ram[254][1] , \ram[254][0] , \ram[253][15] ,
         \ram[253][14] , \ram[253][13] , \ram[253][12] , \ram[253][11] ,
         \ram[253][10] , \ram[253][9] , \ram[253][8] , \ram[253][7] ,
         \ram[253][6] , \ram[253][5] , \ram[253][4] , \ram[253][3] ,
         \ram[253][2] , \ram[253][1] , \ram[253][0] , \ram[252][15] ,
         \ram[252][14] , \ram[252][13] , \ram[252][12] , \ram[252][11] ,
         \ram[252][10] , \ram[252][9] , \ram[252][8] , \ram[252][7] ,
         \ram[252][6] , \ram[252][5] , \ram[252][4] , \ram[252][3] ,
         \ram[252][2] , \ram[252][1] , \ram[252][0] , \ram[251][15] ,
         \ram[251][14] , \ram[251][13] , \ram[251][12] , \ram[251][11] ,
         \ram[251][10] , \ram[251][9] , \ram[251][8] , \ram[251][7] ,
         \ram[251][6] , \ram[251][5] , \ram[251][4] , \ram[251][3] ,
         \ram[251][2] , \ram[251][1] , \ram[251][0] , \ram[250][15] ,
         \ram[250][14] , \ram[250][13] , \ram[250][12] , \ram[250][11] ,
         \ram[250][10] , \ram[250][9] , \ram[250][8] , \ram[250][7] ,
         \ram[250][6] , \ram[250][5] , \ram[250][4] , \ram[250][3] ,
         \ram[250][2] , \ram[250][1] , \ram[250][0] , \ram[249][15] ,
         \ram[249][14] , \ram[249][13] , \ram[249][12] , \ram[249][11] ,
         \ram[249][10] , \ram[249][9] , \ram[249][8] , \ram[249][7] ,
         \ram[249][6] , \ram[249][5] , \ram[249][4] , \ram[249][3] ,
         \ram[249][2] , \ram[249][1] , \ram[249][0] , \ram[248][15] ,
         \ram[248][14] , \ram[248][13] , \ram[248][12] , \ram[248][11] ,
         \ram[248][10] , \ram[248][9] , \ram[248][8] , \ram[248][7] ,
         \ram[248][6] , \ram[248][5] , \ram[248][4] , \ram[248][3] ,
         \ram[248][2] , \ram[248][1] , \ram[248][0] , \ram[247][15] ,
         \ram[247][14] , \ram[247][13] , \ram[247][12] , \ram[247][11] ,
         \ram[247][10] , \ram[247][9] , \ram[247][8] , \ram[247][7] ,
         \ram[247][6] , \ram[247][5] , \ram[247][4] , \ram[247][3] ,
         \ram[247][2] , \ram[247][1] , \ram[247][0] , \ram[246][15] ,
         \ram[246][14] , \ram[246][13] , \ram[246][12] , \ram[246][11] ,
         \ram[246][10] , \ram[246][9] , \ram[246][8] , \ram[246][7] ,
         \ram[246][6] , \ram[246][5] , \ram[246][4] , \ram[246][3] ,
         \ram[246][2] , \ram[246][1] , \ram[246][0] , \ram[245][15] ,
         \ram[245][14] , \ram[245][13] , \ram[245][12] , \ram[245][11] ,
         \ram[245][10] , \ram[245][9] , \ram[245][8] , \ram[245][7] ,
         \ram[245][6] , \ram[245][5] , \ram[245][4] , \ram[245][3] ,
         \ram[245][2] , \ram[245][1] , \ram[245][0] , \ram[244][15] ,
         \ram[244][14] , \ram[244][13] , \ram[244][12] , \ram[244][11] ,
         \ram[244][10] , \ram[244][9] , \ram[244][8] , \ram[244][7] ,
         \ram[244][6] , \ram[244][5] , \ram[244][4] , \ram[244][3] ,
         \ram[244][2] , \ram[244][1] , \ram[244][0] , \ram[243][15] ,
         \ram[243][14] , \ram[243][13] , \ram[243][12] , \ram[243][11] ,
         \ram[243][10] , \ram[243][9] , \ram[243][8] , \ram[243][7] ,
         \ram[243][6] , \ram[243][5] , \ram[243][4] , \ram[243][3] ,
         \ram[243][2] , \ram[243][1] , \ram[243][0] , \ram[242][15] ,
         \ram[242][14] , \ram[242][13] , \ram[242][12] , \ram[242][11] ,
         \ram[242][10] , \ram[242][9] , \ram[242][8] , \ram[242][7] ,
         \ram[242][6] , \ram[242][5] , \ram[242][4] , \ram[242][3] ,
         \ram[242][2] , \ram[242][1] , \ram[242][0] , \ram[241][15] ,
         \ram[241][14] , \ram[241][13] , \ram[241][12] , \ram[241][11] ,
         \ram[241][10] , \ram[241][9] , \ram[241][8] , \ram[241][7] ,
         \ram[241][6] , \ram[241][5] , \ram[241][4] , \ram[241][3] ,
         \ram[241][2] , \ram[241][1] , \ram[241][0] , \ram[240][15] ,
         \ram[240][14] , \ram[240][13] , \ram[240][12] , \ram[240][11] ,
         \ram[240][10] , \ram[240][9] , \ram[240][8] , \ram[240][7] ,
         \ram[240][6] , \ram[240][5] , \ram[240][4] , \ram[240][3] ,
         \ram[240][2] , \ram[240][1] , \ram[240][0] , \ram[239][15] ,
         \ram[239][14] , \ram[239][13] , \ram[239][12] , \ram[239][11] ,
         \ram[239][10] , \ram[239][9] , \ram[239][8] , \ram[239][7] ,
         \ram[239][6] , \ram[239][5] , \ram[239][4] , \ram[239][3] ,
         \ram[239][2] , \ram[239][1] , \ram[239][0] , \ram[238][15] ,
         \ram[238][14] , \ram[238][13] , \ram[238][12] , \ram[238][11] ,
         \ram[238][10] , \ram[238][9] , \ram[238][8] , \ram[238][7] ,
         \ram[238][6] , \ram[238][5] , \ram[238][4] , \ram[238][3] ,
         \ram[238][2] , \ram[238][1] , \ram[238][0] , \ram[237][15] ,
         \ram[237][14] , \ram[237][13] , \ram[237][12] , \ram[237][11] ,
         \ram[237][10] , \ram[237][9] , \ram[237][8] , \ram[237][7] ,
         \ram[237][6] , \ram[237][5] , \ram[237][4] , \ram[237][3] ,
         \ram[237][2] , \ram[237][1] , \ram[237][0] , \ram[236][15] ,
         \ram[236][14] , \ram[236][13] , \ram[236][12] , \ram[236][11] ,
         \ram[236][10] , \ram[236][9] , \ram[236][8] , \ram[236][7] ,
         \ram[236][6] , \ram[236][5] , \ram[236][4] , \ram[236][3] ,
         \ram[236][2] , \ram[236][1] , \ram[236][0] , \ram[235][15] ,
         \ram[235][14] , \ram[235][13] , \ram[235][12] , \ram[235][11] ,
         \ram[235][10] , \ram[235][9] , \ram[235][8] , \ram[235][7] ,
         \ram[235][6] , \ram[235][5] , \ram[235][4] , \ram[235][3] ,
         \ram[235][2] , \ram[235][1] , \ram[235][0] , \ram[234][15] ,
         \ram[234][14] , \ram[234][13] , \ram[234][12] , \ram[234][11] ,
         \ram[234][10] , \ram[234][9] , \ram[234][8] , \ram[234][7] ,
         \ram[234][6] , \ram[234][5] , \ram[234][4] , \ram[234][3] ,
         \ram[234][2] , \ram[234][1] , \ram[234][0] , \ram[233][15] ,
         \ram[233][14] , \ram[233][13] , \ram[233][12] , \ram[233][11] ,
         \ram[233][10] , \ram[233][9] , \ram[233][8] , \ram[233][7] ,
         \ram[233][6] , \ram[233][5] , \ram[233][4] , \ram[233][3] ,
         \ram[233][2] , \ram[233][1] , \ram[233][0] , \ram[232][15] ,
         \ram[232][14] , \ram[232][13] , \ram[232][12] , \ram[232][11] ,
         \ram[232][10] , \ram[232][9] , \ram[232][8] , \ram[232][7] ,
         \ram[232][6] , \ram[232][5] , \ram[232][4] , \ram[232][3] ,
         \ram[232][2] , \ram[232][1] , \ram[232][0] , \ram[231][15] ,
         \ram[231][14] , \ram[231][13] , \ram[231][12] , \ram[231][11] ,
         \ram[231][10] , \ram[231][9] , \ram[231][8] , \ram[231][7] ,
         \ram[231][6] , \ram[231][5] , \ram[231][4] , \ram[231][3] ,
         \ram[231][2] , \ram[231][1] , \ram[231][0] , \ram[230][15] ,
         \ram[230][14] , \ram[230][13] , \ram[230][12] , \ram[230][11] ,
         \ram[230][10] , \ram[230][9] , \ram[230][8] , \ram[230][7] ,
         \ram[230][6] , \ram[230][5] , \ram[230][4] , \ram[230][3] ,
         \ram[230][2] , \ram[230][1] , \ram[230][0] , \ram[229][15] ,
         \ram[229][14] , \ram[229][13] , \ram[229][12] , \ram[229][11] ,
         \ram[229][10] , \ram[229][9] , \ram[229][8] , \ram[229][7] ,
         \ram[229][6] , \ram[229][5] , \ram[229][4] , \ram[229][3] ,
         \ram[229][2] , \ram[229][1] , \ram[229][0] , \ram[228][15] ,
         \ram[228][14] , \ram[228][13] , \ram[228][12] , \ram[228][11] ,
         \ram[228][10] , \ram[228][9] , \ram[228][8] , \ram[228][7] ,
         \ram[228][6] , \ram[228][5] , \ram[228][4] , \ram[228][3] ,
         \ram[228][2] , \ram[228][1] , \ram[228][0] , \ram[227][15] ,
         \ram[227][14] , \ram[227][13] , \ram[227][12] , \ram[227][11] ,
         \ram[227][10] , \ram[227][9] , \ram[227][8] , \ram[227][7] ,
         \ram[227][6] , \ram[227][5] , \ram[227][4] , \ram[227][3] ,
         \ram[227][2] , \ram[227][1] , \ram[227][0] , \ram[226][15] ,
         \ram[226][14] , \ram[226][13] , \ram[226][12] , \ram[226][11] ,
         \ram[226][10] , \ram[226][9] , \ram[226][8] , \ram[226][7] ,
         \ram[226][6] , \ram[226][5] , \ram[226][4] , \ram[226][3] ,
         \ram[226][2] , \ram[226][1] , \ram[226][0] , \ram[225][15] ,
         \ram[225][14] , \ram[225][13] , \ram[225][12] , \ram[225][11] ,
         \ram[225][10] , \ram[225][9] , \ram[225][8] , \ram[225][7] ,
         \ram[225][6] , \ram[225][5] , \ram[225][4] , \ram[225][3] ,
         \ram[225][2] , \ram[225][1] , \ram[225][0] , \ram[224][15] ,
         \ram[224][14] , \ram[224][13] , \ram[224][12] , \ram[224][11] ,
         \ram[224][10] , \ram[224][9] , \ram[224][8] , \ram[224][7] ,
         \ram[224][6] , \ram[224][5] , \ram[224][4] , \ram[224][3] ,
         \ram[224][2] , \ram[224][1] , \ram[224][0] , \ram[223][15] ,
         \ram[223][14] , \ram[223][13] , \ram[223][12] , \ram[223][11] ,
         \ram[223][10] , \ram[223][9] , \ram[223][8] , \ram[223][7] ,
         \ram[223][6] , \ram[223][5] , \ram[223][4] , \ram[223][3] ,
         \ram[223][2] , \ram[223][1] , \ram[223][0] , \ram[222][15] ,
         \ram[222][14] , \ram[222][13] , \ram[222][12] , \ram[222][11] ,
         \ram[222][10] , \ram[222][9] , \ram[222][8] , \ram[222][7] ,
         \ram[222][6] , \ram[222][5] , \ram[222][4] , \ram[222][3] ,
         \ram[222][2] , \ram[222][1] , \ram[222][0] , \ram[221][15] ,
         \ram[221][14] , \ram[221][13] , \ram[221][12] , \ram[221][11] ,
         \ram[221][10] , \ram[221][9] , \ram[221][8] , \ram[221][7] ,
         \ram[221][6] , \ram[221][5] , \ram[221][4] , \ram[221][3] ,
         \ram[221][2] , \ram[221][1] , \ram[221][0] , \ram[220][15] ,
         \ram[220][14] , \ram[220][13] , \ram[220][12] , \ram[220][11] ,
         \ram[220][10] , \ram[220][9] , \ram[220][8] , \ram[220][7] ,
         \ram[220][6] , \ram[220][5] , \ram[220][4] , \ram[220][3] ,
         \ram[220][2] , \ram[220][1] , \ram[220][0] , \ram[219][15] ,
         \ram[219][14] , \ram[219][13] , \ram[219][12] , \ram[219][11] ,
         \ram[219][10] , \ram[219][9] , \ram[219][8] , \ram[219][7] ,
         \ram[219][6] , \ram[219][5] , \ram[219][4] , \ram[219][3] ,
         \ram[219][2] , \ram[219][1] , \ram[219][0] , \ram[218][15] ,
         \ram[218][14] , \ram[218][13] , \ram[218][12] , \ram[218][11] ,
         \ram[218][10] , \ram[218][9] , \ram[218][8] , \ram[218][7] ,
         \ram[218][6] , \ram[218][5] , \ram[218][4] , \ram[218][3] ,
         \ram[218][2] , \ram[218][1] , \ram[218][0] , \ram[217][15] ,
         \ram[217][14] , \ram[217][13] , \ram[217][12] , \ram[217][11] ,
         \ram[217][10] , \ram[217][9] , \ram[217][8] , \ram[217][7] ,
         \ram[217][6] , \ram[217][5] , \ram[217][4] , \ram[217][3] ,
         \ram[217][2] , \ram[217][1] , \ram[217][0] , \ram[216][15] ,
         \ram[216][14] , \ram[216][13] , \ram[216][12] , \ram[216][11] ,
         \ram[216][10] , \ram[216][9] , \ram[216][8] , \ram[216][7] ,
         \ram[216][6] , \ram[216][5] , \ram[216][4] , \ram[216][3] ,
         \ram[216][2] , \ram[216][1] , \ram[216][0] , \ram[215][15] ,
         \ram[215][14] , \ram[215][13] , \ram[215][12] , \ram[215][11] ,
         \ram[215][10] , \ram[215][9] , \ram[215][8] , \ram[215][7] ,
         \ram[215][6] , \ram[215][5] , \ram[215][4] , \ram[215][3] ,
         \ram[215][2] , \ram[215][1] , \ram[215][0] , \ram[214][15] ,
         \ram[214][14] , \ram[214][13] , \ram[214][12] , \ram[214][11] ,
         \ram[214][10] , \ram[214][9] , \ram[214][8] , \ram[214][7] ,
         \ram[214][6] , \ram[214][5] , \ram[214][4] , \ram[214][3] ,
         \ram[214][2] , \ram[214][1] , \ram[214][0] , \ram[213][15] ,
         \ram[213][14] , \ram[213][13] , \ram[213][12] , \ram[213][11] ,
         \ram[213][10] , \ram[213][9] , \ram[213][8] , \ram[213][7] ,
         \ram[213][6] , \ram[213][5] , \ram[213][4] , \ram[213][3] ,
         \ram[213][2] , \ram[213][1] , \ram[213][0] , \ram[212][15] ,
         \ram[212][14] , \ram[212][13] , \ram[212][12] , \ram[212][11] ,
         \ram[212][10] , \ram[212][9] , \ram[212][8] , \ram[212][7] ,
         \ram[212][6] , \ram[212][5] , \ram[212][4] , \ram[212][3] ,
         \ram[212][2] , \ram[212][1] , \ram[212][0] , \ram[211][15] ,
         \ram[211][14] , \ram[211][13] , \ram[211][12] , \ram[211][11] ,
         \ram[211][10] , \ram[211][9] , \ram[211][8] , \ram[211][7] ,
         \ram[211][6] , \ram[211][5] , \ram[211][4] , \ram[211][3] ,
         \ram[211][2] , \ram[211][1] , \ram[211][0] , \ram[210][15] ,
         \ram[210][14] , \ram[210][13] , \ram[210][12] , \ram[210][11] ,
         \ram[210][10] , \ram[210][9] , \ram[210][8] , \ram[210][7] ,
         \ram[210][6] , \ram[210][5] , \ram[210][4] , \ram[210][3] ,
         \ram[210][2] , \ram[210][1] , \ram[210][0] , \ram[209][15] ,
         \ram[209][14] , \ram[209][13] , \ram[209][12] , \ram[209][11] ,
         \ram[209][10] , \ram[209][9] , \ram[209][8] , \ram[209][7] ,
         \ram[209][6] , \ram[209][5] , \ram[209][4] , \ram[209][3] ,
         \ram[209][2] , \ram[209][1] , \ram[209][0] , \ram[208][15] ,
         \ram[208][14] , \ram[208][13] , \ram[208][12] , \ram[208][11] ,
         \ram[208][10] , \ram[208][9] , \ram[208][8] , \ram[208][7] ,
         \ram[208][6] , \ram[208][5] , \ram[208][4] , \ram[208][3] ,
         \ram[208][2] , \ram[208][1] , \ram[208][0] , \ram[207][15] ,
         \ram[207][14] , \ram[207][13] , \ram[207][12] , \ram[207][11] ,
         \ram[207][10] , \ram[207][9] , \ram[207][8] , \ram[207][7] ,
         \ram[207][6] , \ram[207][5] , \ram[207][4] , \ram[207][3] ,
         \ram[207][2] , \ram[207][1] , \ram[207][0] , \ram[206][15] ,
         \ram[206][14] , \ram[206][13] , \ram[206][12] , \ram[206][11] ,
         \ram[206][10] , \ram[206][9] , \ram[206][8] , \ram[206][7] ,
         \ram[206][6] , \ram[206][5] , \ram[206][4] , \ram[206][3] ,
         \ram[206][2] , \ram[206][1] , \ram[206][0] , \ram[205][15] ,
         \ram[205][14] , \ram[205][13] , \ram[205][12] , \ram[205][11] ,
         \ram[205][10] , \ram[205][9] , \ram[205][8] , \ram[205][7] ,
         \ram[205][6] , \ram[205][5] , \ram[205][4] , \ram[205][3] ,
         \ram[205][2] , \ram[205][1] , \ram[205][0] , \ram[204][15] ,
         \ram[204][14] , \ram[204][13] , \ram[204][12] , \ram[204][11] ,
         \ram[204][10] , \ram[204][9] , \ram[204][8] , \ram[204][7] ,
         \ram[204][6] , \ram[204][5] , \ram[204][4] , \ram[204][3] ,
         \ram[204][2] , \ram[204][1] , \ram[204][0] , \ram[203][15] ,
         \ram[203][14] , \ram[203][13] , \ram[203][12] , \ram[203][11] ,
         \ram[203][10] , \ram[203][9] , \ram[203][8] , \ram[203][7] ,
         \ram[203][6] , \ram[203][5] , \ram[203][4] , \ram[203][3] ,
         \ram[203][2] , \ram[203][1] , \ram[203][0] , \ram[202][15] ,
         \ram[202][14] , \ram[202][13] , \ram[202][12] , \ram[202][11] ,
         \ram[202][10] , \ram[202][9] , \ram[202][8] , \ram[202][7] ,
         \ram[202][6] , \ram[202][5] , \ram[202][4] , \ram[202][3] ,
         \ram[202][2] , \ram[202][1] , \ram[202][0] , \ram[201][15] ,
         \ram[201][14] , \ram[201][13] , \ram[201][12] , \ram[201][11] ,
         \ram[201][10] , \ram[201][9] , \ram[201][8] , \ram[201][7] ,
         \ram[201][6] , \ram[201][5] , \ram[201][4] , \ram[201][3] ,
         \ram[201][2] , \ram[201][1] , \ram[201][0] , \ram[200][15] ,
         \ram[200][14] , \ram[200][13] , \ram[200][12] , \ram[200][11] ,
         \ram[200][10] , \ram[200][9] , \ram[200][8] , \ram[200][7] ,
         \ram[200][6] , \ram[200][5] , \ram[200][4] , \ram[200][3] ,
         \ram[200][2] , \ram[200][1] , \ram[200][0] , \ram[199][15] ,
         \ram[199][14] , \ram[199][13] , \ram[199][12] , \ram[199][11] ,
         \ram[199][10] , \ram[199][9] , \ram[199][8] , \ram[199][7] ,
         \ram[199][6] , \ram[199][5] , \ram[199][4] , \ram[199][3] ,
         \ram[199][2] , \ram[199][1] , \ram[199][0] , \ram[198][15] ,
         \ram[198][14] , \ram[198][13] , \ram[198][12] , \ram[198][11] ,
         \ram[198][10] , \ram[198][9] , \ram[198][8] , \ram[198][7] ,
         \ram[198][6] , \ram[198][5] , \ram[198][4] , \ram[198][3] ,
         \ram[198][2] , \ram[198][1] , \ram[198][0] , \ram[197][15] ,
         \ram[197][14] , \ram[197][13] , \ram[197][12] , \ram[197][11] ,
         \ram[197][10] , \ram[197][9] , \ram[197][8] , \ram[197][7] ,
         \ram[197][6] , \ram[197][5] , \ram[197][4] , \ram[197][3] ,
         \ram[197][2] , \ram[197][1] , \ram[197][0] , \ram[196][15] ,
         \ram[196][14] , \ram[196][13] , \ram[196][12] , \ram[196][11] ,
         \ram[196][10] , \ram[196][9] , \ram[196][8] , \ram[196][7] ,
         \ram[196][6] , \ram[196][5] , \ram[196][4] , \ram[196][3] ,
         \ram[196][2] , \ram[196][1] , \ram[196][0] , \ram[195][15] ,
         \ram[195][14] , \ram[195][13] , \ram[195][12] , \ram[195][11] ,
         \ram[195][10] , \ram[195][9] , \ram[195][8] , \ram[195][7] ,
         \ram[195][6] , \ram[195][5] , \ram[195][4] , \ram[195][3] ,
         \ram[195][2] , \ram[195][1] , \ram[195][0] , \ram[194][15] ,
         \ram[194][14] , \ram[194][13] , \ram[194][12] , \ram[194][11] ,
         \ram[194][10] , \ram[194][9] , \ram[194][8] , \ram[194][7] ,
         \ram[194][6] , \ram[194][5] , \ram[194][4] , \ram[194][3] ,
         \ram[194][2] , \ram[194][1] , \ram[194][0] , \ram[193][15] ,
         \ram[193][14] , \ram[193][13] , \ram[193][12] , \ram[193][11] ,
         \ram[193][10] , \ram[193][9] , \ram[193][8] , \ram[193][7] ,
         \ram[193][6] , \ram[193][5] , \ram[193][4] , \ram[193][3] ,
         \ram[193][2] , \ram[193][1] , \ram[193][0] , \ram[192][15] ,
         \ram[192][14] , \ram[192][13] , \ram[192][12] , \ram[192][11] ,
         \ram[192][10] , \ram[192][9] , \ram[192][8] , \ram[192][7] ,
         \ram[192][6] , \ram[192][5] , \ram[192][4] , \ram[192][3] ,
         \ram[192][2] , \ram[192][1] , \ram[192][0] , \ram[191][15] ,
         \ram[191][14] , \ram[191][13] , \ram[191][12] , \ram[191][11] ,
         \ram[191][10] , \ram[191][9] , \ram[191][8] , \ram[191][7] ,
         \ram[191][6] , \ram[191][5] , \ram[191][4] , \ram[191][3] ,
         \ram[191][2] , \ram[191][1] , \ram[191][0] , \ram[190][15] ,
         \ram[190][14] , \ram[190][13] , \ram[190][12] , \ram[190][11] ,
         \ram[190][10] , \ram[190][9] , \ram[190][8] , \ram[190][7] ,
         \ram[190][6] , \ram[190][5] , \ram[190][4] , \ram[190][3] ,
         \ram[190][2] , \ram[190][1] , \ram[190][0] , \ram[189][15] ,
         \ram[189][14] , \ram[189][13] , \ram[189][12] , \ram[189][11] ,
         \ram[189][10] , \ram[189][9] , \ram[189][8] , \ram[189][7] ,
         \ram[189][6] , \ram[189][5] , \ram[189][4] , \ram[189][3] ,
         \ram[189][2] , \ram[189][1] , \ram[189][0] , \ram[188][15] ,
         \ram[188][14] , \ram[188][13] , \ram[188][12] , \ram[188][11] ,
         \ram[188][10] , \ram[188][9] , \ram[188][8] , \ram[188][7] ,
         \ram[188][6] , \ram[188][5] , \ram[188][4] , \ram[188][3] ,
         \ram[188][2] , \ram[188][1] , \ram[188][0] , \ram[187][15] ,
         \ram[187][14] , \ram[187][13] , \ram[187][12] , \ram[187][11] ,
         \ram[187][10] , \ram[187][9] , \ram[187][8] , \ram[187][7] ,
         \ram[187][6] , \ram[187][5] , \ram[187][4] , \ram[187][3] ,
         \ram[187][2] , \ram[187][1] , \ram[187][0] , \ram[186][15] ,
         \ram[186][14] , \ram[186][13] , \ram[186][12] , \ram[186][11] ,
         \ram[186][10] , \ram[186][9] , \ram[186][8] , \ram[186][7] ,
         \ram[186][6] , \ram[186][5] , \ram[186][4] , \ram[186][3] ,
         \ram[186][2] , \ram[186][1] , \ram[186][0] , \ram[185][15] ,
         \ram[185][14] , \ram[185][13] , \ram[185][12] , \ram[185][11] ,
         \ram[185][10] , \ram[185][9] , \ram[185][8] , \ram[185][7] ,
         \ram[185][6] , \ram[185][5] , \ram[185][4] , \ram[185][3] ,
         \ram[185][2] , \ram[185][1] , \ram[185][0] , \ram[184][15] ,
         \ram[184][14] , \ram[184][13] , \ram[184][12] , \ram[184][11] ,
         \ram[184][10] , \ram[184][9] , \ram[184][8] , \ram[184][7] ,
         \ram[184][6] , \ram[184][5] , \ram[184][4] , \ram[184][3] ,
         \ram[184][2] , \ram[184][1] , \ram[184][0] , \ram[183][15] ,
         \ram[183][14] , \ram[183][13] , \ram[183][12] , \ram[183][11] ,
         \ram[183][10] , \ram[183][9] , \ram[183][8] , \ram[183][7] ,
         \ram[183][6] , \ram[183][5] , \ram[183][4] , \ram[183][3] ,
         \ram[183][2] , \ram[183][1] , \ram[183][0] , \ram[182][15] ,
         \ram[182][14] , \ram[182][13] , \ram[182][12] , \ram[182][11] ,
         \ram[182][10] , \ram[182][9] , \ram[182][8] , \ram[182][7] ,
         \ram[182][6] , \ram[182][5] , \ram[182][4] , \ram[182][3] ,
         \ram[182][2] , \ram[182][1] , \ram[182][0] , \ram[181][15] ,
         \ram[181][14] , \ram[181][13] , \ram[181][12] , \ram[181][11] ,
         \ram[181][10] , \ram[181][9] , \ram[181][8] , \ram[181][7] ,
         \ram[181][6] , \ram[181][5] , \ram[181][4] , \ram[181][3] ,
         \ram[181][2] , \ram[181][1] , \ram[181][0] , \ram[180][15] ,
         \ram[180][14] , \ram[180][13] , \ram[180][12] , \ram[180][11] ,
         \ram[180][10] , \ram[180][9] , \ram[180][8] , \ram[180][7] ,
         \ram[180][6] , \ram[180][5] , \ram[180][4] , \ram[180][3] ,
         \ram[180][2] , \ram[180][1] , \ram[180][0] , \ram[179][15] ,
         \ram[179][14] , \ram[179][13] , \ram[179][12] , \ram[179][11] ,
         \ram[179][10] , \ram[179][9] , \ram[179][8] , \ram[179][7] ,
         \ram[179][6] , \ram[179][5] , \ram[179][4] , \ram[179][3] ,
         \ram[179][2] , \ram[179][1] , \ram[179][0] , \ram[178][15] ,
         \ram[178][14] , \ram[178][13] , \ram[178][12] , \ram[178][11] ,
         \ram[178][10] , \ram[178][9] , \ram[178][8] , \ram[178][7] ,
         \ram[178][6] , \ram[178][5] , \ram[178][4] , \ram[178][3] ,
         \ram[178][2] , \ram[178][1] , \ram[178][0] , \ram[177][15] ,
         \ram[177][14] , \ram[177][13] , \ram[177][12] , \ram[177][11] ,
         \ram[177][10] , \ram[177][9] , \ram[177][8] , \ram[177][7] ,
         \ram[177][6] , \ram[177][5] , \ram[177][4] , \ram[177][3] ,
         \ram[177][2] , \ram[177][1] , \ram[177][0] , \ram[176][15] ,
         \ram[176][14] , \ram[176][13] , \ram[176][12] , \ram[176][11] ,
         \ram[176][10] , \ram[176][9] , \ram[176][8] , \ram[176][7] ,
         \ram[176][6] , \ram[176][5] , \ram[176][4] , \ram[176][3] ,
         \ram[176][2] , \ram[176][1] , \ram[176][0] , \ram[175][15] ,
         \ram[175][14] , \ram[175][13] , \ram[175][12] , \ram[175][11] ,
         \ram[175][10] , \ram[175][9] , \ram[175][8] , \ram[175][7] ,
         \ram[175][6] , \ram[175][5] , \ram[175][4] , \ram[175][3] ,
         \ram[175][2] , \ram[175][1] , \ram[175][0] , \ram[174][15] ,
         \ram[174][14] , \ram[174][13] , \ram[174][12] , \ram[174][11] ,
         \ram[174][10] , \ram[174][9] , \ram[174][8] , \ram[174][7] ,
         \ram[174][6] , \ram[174][5] , \ram[174][4] , \ram[174][3] ,
         \ram[174][2] , \ram[174][1] , \ram[174][0] , \ram[173][15] ,
         \ram[173][14] , \ram[173][13] , \ram[173][12] , \ram[173][11] ,
         \ram[173][10] , \ram[173][9] , \ram[173][8] , \ram[173][7] ,
         \ram[173][6] , \ram[173][5] , \ram[173][4] , \ram[173][3] ,
         \ram[173][2] , \ram[173][1] , \ram[173][0] , \ram[172][15] ,
         \ram[172][14] , \ram[172][13] , \ram[172][12] , \ram[172][11] ,
         \ram[172][10] , \ram[172][9] , \ram[172][8] , \ram[172][7] ,
         \ram[172][6] , \ram[172][5] , \ram[172][4] , \ram[172][3] ,
         \ram[172][2] , \ram[172][1] , \ram[172][0] , \ram[171][15] ,
         \ram[171][14] , \ram[171][13] , \ram[171][12] , \ram[171][11] ,
         \ram[171][10] , \ram[171][9] , \ram[171][8] , \ram[171][7] ,
         \ram[171][6] , \ram[171][5] , \ram[171][4] , \ram[171][3] ,
         \ram[171][2] , \ram[171][1] , \ram[171][0] , \ram[170][15] ,
         \ram[170][14] , \ram[170][13] , \ram[170][12] , \ram[170][11] ,
         \ram[170][10] , \ram[170][9] , \ram[170][8] , \ram[170][7] ,
         \ram[170][6] , \ram[170][5] , \ram[170][4] , \ram[170][3] ,
         \ram[170][2] , \ram[170][1] , \ram[170][0] , \ram[169][15] ,
         \ram[169][14] , \ram[169][13] , \ram[169][12] , \ram[169][11] ,
         \ram[169][10] , \ram[169][9] , \ram[169][8] , \ram[169][7] ,
         \ram[169][6] , \ram[169][5] , \ram[169][4] , \ram[169][3] ,
         \ram[169][2] , \ram[169][1] , \ram[169][0] , \ram[168][15] ,
         \ram[168][14] , \ram[168][13] , \ram[168][12] , \ram[168][11] ,
         \ram[168][10] , \ram[168][9] , \ram[168][8] , \ram[168][7] ,
         \ram[168][6] , \ram[168][5] , \ram[168][4] , \ram[168][3] ,
         \ram[168][2] , \ram[168][1] , \ram[168][0] , \ram[167][15] ,
         \ram[167][14] , \ram[167][13] , \ram[167][12] , \ram[167][11] ,
         \ram[167][10] , \ram[167][9] , \ram[167][8] , \ram[167][7] ,
         \ram[167][6] , \ram[167][5] , \ram[167][4] , \ram[167][3] ,
         \ram[167][2] , \ram[167][1] , \ram[167][0] , \ram[166][15] ,
         \ram[166][14] , \ram[166][13] , \ram[166][12] , \ram[166][11] ,
         \ram[166][10] , \ram[166][9] , \ram[166][8] , \ram[166][7] ,
         \ram[166][6] , \ram[166][5] , \ram[166][4] , \ram[166][3] ,
         \ram[166][2] , \ram[166][1] , \ram[166][0] , \ram[165][15] ,
         \ram[165][14] , \ram[165][13] , \ram[165][12] , \ram[165][11] ,
         \ram[165][10] , \ram[165][9] , \ram[165][8] , \ram[165][7] ,
         \ram[165][6] , \ram[165][5] , \ram[165][4] , \ram[165][3] ,
         \ram[165][2] , \ram[165][1] , \ram[165][0] , \ram[164][15] ,
         \ram[164][14] , \ram[164][13] , \ram[164][12] , \ram[164][11] ,
         \ram[164][10] , \ram[164][9] , \ram[164][8] , \ram[164][7] ,
         \ram[164][6] , \ram[164][5] , \ram[164][4] , \ram[164][3] ,
         \ram[164][2] , \ram[164][1] , \ram[164][0] , \ram[163][15] ,
         \ram[163][14] , \ram[163][13] , \ram[163][12] , \ram[163][11] ,
         \ram[163][10] , \ram[163][9] , \ram[163][8] , \ram[163][7] ,
         \ram[163][6] , \ram[163][5] , \ram[163][4] , \ram[163][3] ,
         \ram[163][2] , \ram[163][1] , \ram[163][0] , \ram[162][15] ,
         \ram[162][14] , \ram[162][13] , \ram[162][12] , \ram[162][11] ,
         \ram[162][10] , \ram[162][9] , \ram[162][8] , \ram[162][7] ,
         \ram[162][6] , \ram[162][5] , \ram[162][4] , \ram[162][3] ,
         \ram[162][2] , \ram[162][1] , \ram[162][0] , \ram[161][15] ,
         \ram[161][14] , \ram[161][13] , \ram[161][12] , \ram[161][11] ,
         \ram[161][10] , \ram[161][9] , \ram[161][8] , \ram[161][7] ,
         \ram[161][6] , \ram[161][5] , \ram[161][4] , \ram[161][3] ,
         \ram[161][2] , \ram[161][1] , \ram[161][0] , \ram[160][15] ,
         \ram[160][14] , \ram[160][13] , \ram[160][12] , \ram[160][11] ,
         \ram[160][10] , \ram[160][9] , \ram[160][8] , \ram[160][7] ,
         \ram[160][6] , \ram[160][5] , \ram[160][4] , \ram[160][3] ,
         \ram[160][2] , \ram[160][1] , \ram[160][0] , \ram[159][15] ,
         \ram[159][14] , \ram[159][13] , \ram[159][12] , \ram[159][11] ,
         \ram[159][10] , \ram[159][9] , \ram[159][8] , \ram[159][7] ,
         \ram[159][6] , \ram[159][5] , \ram[159][4] , \ram[159][3] ,
         \ram[159][2] , \ram[159][1] , \ram[159][0] , \ram[158][15] ,
         \ram[158][14] , \ram[158][13] , \ram[158][12] , \ram[158][11] ,
         \ram[158][10] , \ram[158][9] , \ram[158][8] , \ram[158][7] ,
         \ram[158][6] , \ram[158][5] , \ram[158][4] , \ram[158][3] ,
         \ram[158][2] , \ram[158][1] , \ram[158][0] , \ram[157][15] ,
         \ram[157][14] , \ram[157][13] , \ram[157][12] , \ram[157][11] ,
         \ram[157][10] , \ram[157][9] , \ram[157][8] , \ram[157][7] ,
         \ram[157][6] , \ram[157][5] , \ram[157][4] , \ram[157][3] ,
         \ram[157][2] , \ram[157][1] , \ram[157][0] , \ram[156][15] ,
         \ram[156][14] , \ram[156][13] , \ram[156][12] , \ram[156][11] ,
         \ram[156][10] , \ram[156][9] , \ram[156][8] , \ram[156][7] ,
         \ram[156][6] , \ram[156][5] , \ram[156][4] , \ram[156][3] ,
         \ram[156][2] , \ram[156][1] , \ram[156][0] , \ram[155][15] ,
         \ram[155][14] , \ram[155][13] , \ram[155][12] , \ram[155][11] ,
         \ram[155][10] , \ram[155][9] , \ram[155][8] , \ram[155][7] ,
         \ram[155][6] , \ram[155][5] , \ram[155][4] , \ram[155][3] ,
         \ram[155][2] , \ram[155][1] , \ram[155][0] , \ram[154][15] ,
         \ram[154][14] , \ram[154][13] , \ram[154][12] , \ram[154][11] ,
         \ram[154][10] , \ram[154][9] , \ram[154][8] , \ram[154][7] ,
         \ram[154][6] , \ram[154][5] , \ram[154][4] , \ram[154][3] ,
         \ram[154][2] , \ram[154][1] , \ram[154][0] , \ram[153][15] ,
         \ram[153][14] , \ram[153][13] , \ram[153][12] , \ram[153][11] ,
         \ram[153][10] , \ram[153][9] , \ram[153][8] , \ram[153][7] ,
         \ram[153][6] , \ram[153][5] , \ram[153][4] , \ram[153][3] ,
         \ram[153][2] , \ram[153][1] , \ram[153][0] , \ram[152][15] ,
         \ram[152][14] , \ram[152][13] , \ram[152][12] , \ram[152][11] ,
         \ram[152][10] , \ram[152][9] , \ram[152][8] , \ram[152][7] ,
         \ram[152][6] , \ram[152][5] , \ram[152][4] , \ram[152][3] ,
         \ram[152][2] , \ram[152][1] , \ram[152][0] , \ram[151][15] ,
         \ram[151][14] , \ram[151][13] , \ram[151][12] , \ram[151][11] ,
         \ram[151][10] , \ram[151][9] , \ram[151][8] , \ram[151][7] ,
         \ram[151][6] , \ram[151][5] , \ram[151][4] , \ram[151][3] ,
         \ram[151][2] , \ram[151][1] , \ram[151][0] , \ram[150][15] ,
         \ram[150][14] , \ram[150][13] , \ram[150][12] , \ram[150][11] ,
         \ram[150][10] , \ram[150][9] , \ram[150][8] , \ram[150][7] ,
         \ram[150][6] , \ram[150][5] , \ram[150][4] , \ram[150][3] ,
         \ram[150][2] , \ram[150][1] , \ram[150][0] , \ram[149][15] ,
         \ram[149][14] , \ram[149][13] , \ram[149][12] , \ram[149][11] ,
         \ram[149][10] , \ram[149][9] , \ram[149][8] , \ram[149][7] ,
         \ram[149][6] , \ram[149][5] , \ram[149][4] , \ram[149][3] ,
         \ram[149][2] , \ram[149][1] , \ram[149][0] , \ram[148][15] ,
         \ram[148][14] , \ram[148][13] , \ram[148][12] , \ram[148][11] ,
         \ram[148][10] , \ram[148][9] , \ram[148][8] , \ram[148][7] ,
         \ram[148][6] , \ram[148][5] , \ram[148][4] , \ram[148][3] ,
         \ram[148][2] , \ram[148][1] , \ram[148][0] , \ram[147][15] ,
         \ram[147][14] , \ram[147][13] , \ram[147][12] , \ram[147][11] ,
         \ram[147][10] , \ram[147][9] , \ram[147][8] , \ram[147][7] ,
         \ram[147][6] , \ram[147][5] , \ram[147][4] , \ram[147][3] ,
         \ram[147][2] , \ram[147][1] , \ram[147][0] , \ram[146][15] ,
         \ram[146][14] , \ram[146][13] , \ram[146][12] , \ram[146][11] ,
         \ram[146][10] , \ram[146][9] , \ram[146][8] , \ram[146][7] ,
         \ram[146][6] , \ram[146][5] , \ram[146][4] , \ram[146][3] ,
         \ram[146][2] , \ram[146][1] , \ram[146][0] , \ram[145][15] ,
         \ram[145][14] , \ram[145][13] , \ram[145][12] , \ram[145][11] ,
         \ram[145][10] , \ram[145][9] , \ram[145][8] , \ram[145][7] ,
         \ram[145][6] , \ram[145][5] , \ram[145][4] , \ram[145][3] ,
         \ram[145][2] , \ram[145][1] , \ram[145][0] , \ram[144][15] ,
         \ram[144][14] , \ram[144][13] , \ram[144][12] , \ram[144][11] ,
         \ram[144][10] , \ram[144][9] , \ram[144][8] , \ram[144][7] ,
         \ram[144][6] , \ram[144][5] , \ram[144][4] , \ram[144][3] ,
         \ram[144][2] , \ram[144][1] , \ram[144][0] , \ram[143][15] ,
         \ram[143][14] , \ram[143][13] , \ram[143][12] , \ram[143][11] ,
         \ram[143][10] , \ram[143][9] , \ram[143][8] , \ram[143][7] ,
         \ram[143][6] , \ram[143][5] , \ram[143][4] , \ram[143][3] ,
         \ram[143][2] , \ram[143][1] , \ram[143][0] , \ram[142][15] ,
         \ram[142][14] , \ram[142][13] , \ram[142][12] , \ram[142][11] ,
         \ram[142][10] , \ram[142][9] , \ram[142][8] , \ram[142][7] ,
         \ram[142][6] , \ram[142][5] , \ram[142][4] , \ram[142][3] ,
         \ram[142][2] , \ram[142][1] , \ram[142][0] , \ram[141][15] ,
         \ram[141][14] , \ram[141][13] , \ram[141][12] , \ram[141][11] ,
         \ram[141][10] , \ram[141][9] , \ram[141][8] , \ram[141][7] ,
         \ram[141][6] , \ram[141][5] , \ram[141][4] , \ram[141][3] ,
         \ram[141][2] , \ram[141][1] , \ram[141][0] , \ram[140][15] ,
         \ram[140][14] , \ram[140][13] , \ram[140][12] , \ram[140][11] ,
         \ram[140][10] , \ram[140][9] , \ram[140][8] , \ram[140][7] ,
         \ram[140][6] , \ram[140][5] , \ram[140][4] , \ram[140][3] ,
         \ram[140][2] , \ram[140][1] , \ram[140][0] , \ram[139][15] ,
         \ram[139][14] , \ram[139][13] , \ram[139][12] , \ram[139][11] ,
         \ram[139][10] , \ram[139][9] , \ram[139][8] , \ram[139][7] ,
         \ram[139][6] , \ram[139][5] , \ram[139][4] , \ram[139][3] ,
         \ram[139][2] , \ram[139][1] , \ram[139][0] , \ram[138][15] ,
         \ram[138][14] , \ram[138][13] , \ram[138][12] , \ram[138][11] ,
         \ram[138][10] , \ram[138][9] , \ram[138][8] , \ram[138][7] ,
         \ram[138][6] , \ram[138][5] , \ram[138][4] , \ram[138][3] ,
         \ram[138][2] , \ram[138][1] , \ram[138][0] , \ram[137][15] ,
         \ram[137][14] , \ram[137][13] , \ram[137][12] , \ram[137][11] ,
         \ram[137][10] , \ram[137][9] , \ram[137][8] , \ram[137][7] ,
         \ram[137][6] , \ram[137][5] , \ram[137][4] , \ram[137][3] ,
         \ram[137][2] , \ram[137][1] , \ram[137][0] , \ram[136][15] ,
         \ram[136][14] , \ram[136][13] , \ram[136][12] , \ram[136][11] ,
         \ram[136][10] , \ram[136][9] , \ram[136][8] , \ram[136][7] ,
         \ram[136][6] , \ram[136][5] , \ram[136][4] , \ram[136][3] ,
         \ram[136][2] , \ram[136][1] , \ram[136][0] , \ram[135][15] ,
         \ram[135][14] , \ram[135][13] , \ram[135][12] , \ram[135][11] ,
         \ram[135][10] , \ram[135][9] , \ram[135][8] , \ram[135][7] ,
         \ram[135][6] , \ram[135][5] , \ram[135][4] , \ram[135][3] ,
         \ram[135][2] , \ram[135][1] , \ram[135][0] , \ram[134][15] ,
         \ram[134][14] , \ram[134][13] , \ram[134][12] , \ram[134][11] ,
         \ram[134][10] , \ram[134][9] , \ram[134][8] , \ram[134][7] ,
         \ram[134][6] , \ram[134][5] , \ram[134][4] , \ram[134][3] ,
         \ram[134][2] , \ram[134][1] , \ram[134][0] , \ram[133][15] ,
         \ram[133][14] , \ram[133][13] , \ram[133][12] , \ram[133][11] ,
         \ram[133][10] , \ram[133][9] , \ram[133][8] , \ram[133][7] ,
         \ram[133][6] , \ram[133][5] , \ram[133][4] , \ram[133][3] ,
         \ram[133][2] , \ram[133][1] , \ram[133][0] , \ram[132][15] ,
         \ram[132][14] , \ram[132][13] , \ram[132][12] , \ram[132][11] ,
         \ram[132][10] , \ram[132][9] , \ram[132][8] , \ram[132][7] ,
         \ram[132][6] , \ram[132][5] , \ram[132][4] , \ram[132][3] ,
         \ram[132][2] , \ram[132][1] , \ram[132][0] , \ram[131][15] ,
         \ram[131][14] , \ram[131][13] , \ram[131][12] , \ram[131][11] ,
         \ram[131][10] , \ram[131][9] , \ram[131][8] , \ram[131][7] ,
         \ram[131][6] , \ram[131][5] , \ram[131][4] , \ram[131][3] ,
         \ram[131][2] , \ram[131][1] , \ram[131][0] , \ram[130][15] ,
         \ram[130][14] , \ram[130][13] , \ram[130][12] , \ram[130][11] ,
         \ram[130][10] , \ram[130][9] , \ram[130][8] , \ram[130][7] ,
         \ram[130][6] , \ram[130][5] , \ram[130][4] , \ram[130][3] ,
         \ram[130][2] , \ram[130][1] , \ram[130][0] , \ram[129][15] ,
         \ram[129][14] , \ram[129][13] , \ram[129][12] , \ram[129][11] ,
         \ram[129][10] , \ram[129][9] , \ram[129][8] , \ram[129][7] ,
         \ram[129][6] , \ram[129][5] , \ram[129][4] , \ram[129][3] ,
         \ram[129][2] , \ram[129][1] , \ram[129][0] , \ram[128][15] ,
         \ram[128][14] , \ram[128][13] , \ram[128][12] , \ram[128][11] ,
         \ram[128][10] , \ram[128][9] , \ram[128][8] , \ram[128][7] ,
         \ram[128][6] , \ram[128][5] , \ram[128][4] , \ram[128][3] ,
         \ram[128][2] , \ram[128][1] , \ram[128][0] , \ram[127][15] ,
         \ram[127][14] , \ram[127][13] , \ram[127][12] , \ram[127][11] ,
         \ram[127][10] , \ram[127][9] , \ram[127][8] , \ram[127][7] ,
         \ram[127][6] , \ram[127][5] , \ram[127][4] , \ram[127][3] ,
         \ram[127][2] , \ram[127][1] , \ram[127][0] , \ram[126][15] ,
         \ram[126][14] , \ram[126][13] , \ram[126][12] , \ram[126][11] ,
         \ram[126][10] , \ram[126][9] , \ram[126][8] , \ram[126][7] ,
         \ram[126][6] , \ram[126][5] , \ram[126][4] , \ram[126][3] ,
         \ram[126][2] , \ram[126][1] , \ram[126][0] , \ram[125][15] ,
         \ram[125][14] , \ram[125][13] , \ram[125][12] , \ram[125][11] ,
         \ram[125][10] , \ram[125][9] , \ram[125][8] , \ram[125][7] ,
         \ram[125][6] , \ram[125][5] , \ram[125][4] , \ram[125][3] ,
         \ram[125][2] , \ram[125][1] , \ram[125][0] , \ram[124][15] ,
         \ram[124][14] , \ram[124][13] , \ram[124][12] , \ram[124][11] ,
         \ram[124][10] , \ram[124][9] , \ram[124][8] , \ram[124][7] ,
         \ram[124][6] , \ram[124][5] , \ram[124][4] , \ram[124][3] ,
         \ram[124][2] , \ram[124][1] , \ram[124][0] , \ram[123][15] ,
         \ram[123][14] , \ram[123][13] , \ram[123][12] , \ram[123][11] ,
         \ram[123][10] , \ram[123][9] , \ram[123][8] , \ram[123][7] ,
         \ram[123][6] , \ram[123][5] , \ram[123][4] , \ram[123][3] ,
         \ram[123][2] , \ram[123][1] , \ram[123][0] , \ram[122][15] ,
         \ram[122][14] , \ram[122][13] , \ram[122][12] , \ram[122][11] ,
         \ram[122][10] , \ram[122][9] , \ram[122][8] , \ram[122][7] ,
         \ram[122][6] , \ram[122][5] , \ram[122][4] , \ram[122][3] ,
         \ram[122][2] , \ram[122][1] , \ram[122][0] , \ram[121][15] ,
         \ram[121][14] , \ram[121][13] , \ram[121][12] , \ram[121][11] ,
         \ram[121][10] , \ram[121][9] , \ram[121][8] , \ram[121][7] ,
         \ram[121][6] , \ram[121][5] , \ram[121][4] , \ram[121][3] ,
         \ram[121][2] , \ram[121][1] , \ram[121][0] , \ram[120][15] ,
         \ram[120][14] , \ram[120][13] , \ram[120][12] , \ram[120][11] ,
         \ram[120][10] , \ram[120][9] , \ram[120][8] , \ram[120][7] ,
         \ram[120][6] , \ram[120][5] , \ram[120][4] , \ram[120][3] ,
         \ram[120][2] , \ram[120][1] , \ram[120][0] , \ram[119][15] ,
         \ram[119][14] , \ram[119][13] , \ram[119][12] , \ram[119][11] ,
         \ram[119][10] , \ram[119][9] , \ram[119][8] , \ram[119][7] ,
         \ram[119][6] , \ram[119][5] , \ram[119][4] , \ram[119][3] ,
         \ram[119][2] , \ram[119][1] , \ram[119][0] , \ram[118][15] ,
         \ram[118][14] , \ram[118][13] , \ram[118][12] , \ram[118][11] ,
         \ram[118][10] , \ram[118][9] , \ram[118][8] , \ram[118][7] ,
         \ram[118][6] , \ram[118][5] , \ram[118][4] , \ram[118][3] ,
         \ram[118][2] , \ram[118][1] , \ram[118][0] , \ram[117][15] ,
         \ram[117][14] , \ram[117][13] , \ram[117][12] , \ram[117][11] ,
         \ram[117][10] , \ram[117][9] , \ram[117][8] , \ram[117][7] ,
         \ram[117][6] , \ram[117][5] , \ram[117][4] , \ram[117][3] ,
         \ram[117][2] , \ram[117][1] , \ram[117][0] , \ram[116][15] ,
         \ram[116][14] , \ram[116][13] , \ram[116][12] , \ram[116][11] ,
         \ram[116][10] , \ram[116][9] , \ram[116][8] , \ram[116][7] ,
         \ram[116][6] , \ram[116][5] , \ram[116][4] , \ram[116][3] ,
         \ram[116][2] , \ram[116][1] , \ram[116][0] , \ram[115][15] ,
         \ram[115][14] , \ram[115][13] , \ram[115][12] , \ram[115][11] ,
         \ram[115][10] , \ram[115][9] , \ram[115][8] , \ram[115][7] ,
         \ram[115][6] , \ram[115][5] , \ram[115][4] , \ram[115][3] ,
         \ram[115][2] , \ram[115][1] , \ram[115][0] , \ram[114][15] ,
         \ram[114][14] , \ram[114][13] , \ram[114][12] , \ram[114][11] ,
         \ram[114][10] , \ram[114][9] , \ram[114][8] , \ram[114][7] ,
         \ram[114][6] , \ram[114][5] , \ram[114][4] , \ram[114][3] ,
         \ram[114][2] , \ram[114][1] , \ram[114][0] , \ram[113][15] ,
         \ram[113][14] , \ram[113][13] , \ram[113][12] , \ram[113][11] ,
         \ram[113][10] , \ram[113][9] , \ram[113][8] , \ram[113][7] ,
         \ram[113][6] , \ram[113][5] , \ram[113][4] , \ram[113][3] ,
         \ram[113][2] , \ram[113][1] , \ram[113][0] , \ram[112][15] ,
         \ram[112][14] , \ram[112][13] , \ram[112][12] , \ram[112][11] ,
         \ram[112][10] , \ram[112][9] , \ram[112][8] , \ram[112][7] ,
         \ram[112][6] , \ram[112][5] , \ram[112][4] , \ram[112][3] ,
         \ram[112][2] , \ram[112][1] , \ram[112][0] , \ram[111][15] ,
         \ram[111][14] , \ram[111][13] , \ram[111][12] , \ram[111][11] ,
         \ram[111][10] , \ram[111][9] , \ram[111][8] , \ram[111][7] ,
         \ram[111][6] , \ram[111][5] , \ram[111][4] , \ram[111][3] ,
         \ram[111][2] , \ram[111][1] , \ram[111][0] , \ram[110][15] ,
         \ram[110][14] , \ram[110][13] , \ram[110][12] , \ram[110][11] ,
         \ram[110][10] , \ram[110][9] , \ram[110][8] , \ram[110][7] ,
         \ram[110][6] , \ram[110][5] , \ram[110][4] , \ram[110][3] ,
         \ram[110][2] , \ram[110][1] , \ram[110][0] , \ram[109][15] ,
         \ram[109][14] , \ram[109][13] , \ram[109][12] , \ram[109][11] ,
         \ram[109][10] , \ram[109][9] , \ram[109][8] , \ram[109][7] ,
         \ram[109][6] , \ram[109][5] , \ram[109][4] , \ram[109][3] ,
         \ram[109][2] , \ram[109][1] , \ram[109][0] , \ram[108][15] ,
         \ram[108][14] , \ram[108][13] , \ram[108][12] , \ram[108][11] ,
         \ram[108][10] , \ram[108][9] , \ram[108][8] , \ram[108][7] ,
         \ram[108][6] , \ram[108][5] , \ram[108][4] , \ram[108][3] ,
         \ram[108][2] , \ram[108][1] , \ram[108][0] , \ram[107][15] ,
         \ram[107][14] , \ram[107][13] , \ram[107][12] , \ram[107][11] ,
         \ram[107][10] , \ram[107][9] , \ram[107][8] , \ram[107][7] ,
         \ram[107][6] , \ram[107][5] , \ram[107][4] , \ram[107][3] ,
         \ram[107][2] , \ram[107][1] , \ram[107][0] , \ram[106][15] ,
         \ram[106][14] , \ram[106][13] , \ram[106][12] , \ram[106][11] ,
         \ram[106][10] , \ram[106][9] , \ram[106][8] , \ram[106][7] ,
         \ram[106][6] , \ram[106][5] , \ram[106][4] , \ram[106][3] ,
         \ram[106][2] , \ram[106][1] , \ram[106][0] , \ram[105][15] ,
         \ram[105][14] , \ram[105][13] , \ram[105][12] , \ram[105][11] ,
         \ram[105][10] , \ram[105][9] , \ram[105][8] , \ram[105][7] ,
         \ram[105][6] , \ram[105][5] , \ram[105][4] , \ram[105][3] ,
         \ram[105][2] , \ram[105][1] , \ram[105][0] , \ram[104][15] ,
         \ram[104][14] , \ram[104][13] , \ram[104][12] , \ram[104][11] ,
         \ram[104][10] , \ram[104][9] , \ram[104][8] , \ram[104][7] ,
         \ram[104][6] , \ram[104][5] , \ram[104][4] , \ram[104][3] ,
         \ram[104][2] , \ram[104][1] , \ram[104][0] , \ram[103][15] ,
         \ram[103][14] , \ram[103][13] , \ram[103][12] , \ram[103][11] ,
         \ram[103][10] , \ram[103][9] , \ram[103][8] , \ram[103][7] ,
         \ram[103][6] , \ram[103][5] , \ram[103][4] , \ram[103][3] ,
         \ram[103][2] , \ram[103][1] , \ram[103][0] , \ram[102][15] ,
         \ram[102][14] , \ram[102][13] , \ram[102][12] , \ram[102][11] ,
         \ram[102][10] , \ram[102][9] , \ram[102][8] , \ram[102][7] ,
         \ram[102][6] , \ram[102][5] , \ram[102][4] , \ram[102][3] ,
         \ram[102][2] , \ram[102][1] , \ram[102][0] , \ram[101][15] ,
         \ram[101][14] , \ram[101][13] , \ram[101][12] , \ram[101][11] ,
         \ram[101][10] , \ram[101][9] , \ram[101][8] , \ram[101][7] ,
         \ram[101][6] , \ram[101][5] , \ram[101][4] , \ram[101][3] ,
         \ram[101][2] , \ram[101][1] , \ram[101][0] , \ram[100][15] ,
         \ram[100][14] , \ram[100][13] , \ram[100][12] , \ram[100][11] ,
         \ram[100][10] , \ram[100][9] , \ram[100][8] , \ram[100][7] ,
         \ram[100][6] , \ram[100][5] , \ram[100][4] , \ram[100][3] ,
         \ram[100][2] , \ram[100][1] , \ram[100][0] , \ram[99][15] ,
         \ram[99][14] , \ram[99][13] , \ram[99][12] , \ram[99][11] ,
         \ram[99][10] , \ram[99][9] , \ram[99][8] , \ram[99][7] , \ram[99][6] ,
         \ram[99][5] , \ram[99][4] , \ram[99][3] , \ram[99][2] , \ram[99][1] ,
         \ram[99][0] , \ram[98][15] , \ram[98][14] , \ram[98][13] ,
         \ram[98][12] , \ram[98][11] , \ram[98][10] , \ram[98][9] ,
         \ram[98][8] , \ram[98][7] , \ram[98][6] , \ram[98][5] , \ram[98][4] ,
         \ram[98][3] , \ram[98][2] , \ram[98][1] , \ram[98][0] , \ram[97][15] ,
         \ram[97][14] , \ram[97][13] , \ram[97][12] , \ram[97][11] ,
         \ram[97][10] , \ram[97][9] , \ram[97][8] , \ram[97][7] , \ram[97][6] ,
         \ram[97][5] , \ram[97][4] , \ram[97][3] , \ram[97][2] , \ram[97][1] ,
         \ram[97][0] , \ram[96][15] , \ram[96][14] , \ram[96][13] ,
         \ram[96][12] , \ram[96][11] , \ram[96][10] , \ram[96][9] ,
         \ram[96][8] , \ram[96][7] , \ram[96][6] , \ram[96][5] , \ram[96][4] ,
         \ram[96][3] , \ram[96][2] , \ram[96][1] , \ram[96][0] , \ram[95][15] ,
         \ram[95][14] , \ram[95][13] , \ram[95][12] , \ram[95][11] ,
         \ram[95][10] , \ram[95][9] , \ram[95][8] , \ram[95][7] , \ram[95][6] ,
         \ram[95][5] , \ram[95][4] , \ram[95][3] , \ram[95][2] , \ram[95][1] ,
         \ram[95][0] , \ram[94][15] , \ram[94][14] , \ram[94][13] ,
         \ram[94][12] , \ram[94][11] , \ram[94][10] , \ram[94][9] ,
         \ram[94][8] , \ram[94][7] , \ram[94][6] , \ram[94][5] , \ram[94][4] ,
         \ram[94][3] , \ram[94][2] , \ram[94][1] , \ram[94][0] , \ram[93][15] ,
         \ram[93][14] , \ram[93][13] , \ram[93][12] , \ram[93][11] ,
         \ram[93][10] , \ram[93][9] , \ram[93][8] , \ram[93][7] , \ram[93][6] ,
         \ram[93][5] , \ram[93][4] , \ram[93][3] , \ram[93][2] , \ram[93][1] ,
         \ram[93][0] , \ram[92][15] , \ram[92][14] , \ram[92][13] ,
         \ram[92][12] , \ram[92][11] , \ram[92][10] , \ram[92][9] ,
         \ram[92][8] , \ram[92][7] , \ram[92][6] , \ram[92][5] , \ram[92][4] ,
         \ram[92][3] , \ram[92][2] , \ram[92][1] , \ram[92][0] , \ram[91][15] ,
         \ram[91][14] , \ram[91][13] , \ram[91][12] , \ram[91][11] ,
         \ram[91][10] , \ram[91][9] , \ram[91][8] , \ram[91][7] , \ram[91][6] ,
         \ram[91][5] , \ram[91][4] , \ram[91][3] , \ram[91][2] , \ram[91][1] ,
         \ram[91][0] , \ram[90][15] , \ram[90][14] , \ram[90][13] ,
         \ram[90][12] , \ram[90][11] , \ram[90][10] , \ram[90][9] ,
         \ram[90][8] , \ram[90][7] , \ram[90][6] , \ram[90][5] , \ram[90][4] ,
         \ram[90][3] , \ram[90][2] , \ram[90][1] , \ram[90][0] , \ram[89][15] ,
         \ram[89][14] , \ram[89][13] , \ram[89][12] , \ram[89][11] ,
         \ram[89][10] , \ram[89][9] , \ram[89][8] , \ram[89][7] , \ram[89][6] ,
         \ram[89][5] , \ram[89][4] , \ram[89][3] , \ram[89][2] , \ram[89][1] ,
         \ram[89][0] , \ram[88][15] , \ram[88][14] , \ram[88][13] ,
         \ram[88][12] , \ram[88][11] , \ram[88][10] , \ram[88][9] ,
         \ram[88][8] , \ram[88][7] , \ram[88][6] , \ram[88][5] , \ram[88][4] ,
         \ram[88][3] , \ram[88][2] , \ram[88][1] , \ram[88][0] , \ram[87][15] ,
         \ram[87][14] , \ram[87][13] , \ram[87][12] , \ram[87][11] ,
         \ram[87][10] , \ram[87][9] , \ram[87][8] , \ram[87][7] , \ram[87][6] ,
         \ram[87][5] , \ram[87][4] , \ram[87][3] , \ram[87][2] , \ram[87][1] ,
         \ram[87][0] , \ram[86][15] , \ram[86][14] , \ram[86][13] ,
         \ram[86][12] , \ram[86][11] , \ram[86][10] , \ram[86][9] ,
         \ram[86][8] , \ram[86][7] , \ram[86][6] , \ram[86][5] , \ram[86][4] ,
         \ram[86][3] , \ram[86][2] , \ram[86][1] , \ram[86][0] , \ram[85][15] ,
         \ram[85][14] , \ram[85][13] , \ram[85][12] , \ram[85][11] ,
         \ram[85][10] , \ram[85][9] , \ram[85][8] , \ram[85][7] , \ram[85][6] ,
         \ram[85][5] , \ram[85][4] , \ram[85][3] , \ram[85][2] , \ram[85][1] ,
         \ram[85][0] , \ram[84][15] , \ram[84][14] , \ram[84][13] ,
         \ram[84][12] , \ram[84][11] , \ram[84][10] , \ram[84][9] ,
         \ram[84][8] , \ram[84][7] , \ram[84][6] , \ram[84][5] , \ram[84][4] ,
         \ram[84][3] , \ram[84][2] , \ram[84][1] , \ram[84][0] , \ram[83][15] ,
         \ram[83][14] , \ram[83][13] , \ram[83][12] , \ram[83][11] ,
         \ram[83][10] , \ram[83][9] , \ram[83][8] , \ram[83][7] , \ram[83][6] ,
         \ram[83][5] , \ram[83][4] , \ram[83][3] , \ram[83][2] , \ram[83][1] ,
         \ram[83][0] , \ram[82][15] , \ram[82][14] , \ram[82][13] ,
         \ram[82][12] , \ram[82][11] , \ram[82][10] , \ram[82][9] ,
         \ram[82][8] , \ram[82][7] , \ram[82][6] , \ram[82][5] , \ram[82][4] ,
         \ram[82][3] , \ram[82][2] , \ram[82][1] , \ram[82][0] , \ram[81][15] ,
         \ram[81][14] , \ram[81][13] , \ram[81][12] , \ram[81][11] ,
         \ram[81][10] , \ram[81][9] , \ram[81][8] , \ram[81][7] , \ram[81][6] ,
         \ram[81][5] , \ram[81][4] , \ram[81][3] , \ram[81][2] , \ram[81][1] ,
         \ram[81][0] , \ram[80][15] , \ram[80][14] , \ram[80][13] ,
         \ram[80][12] , \ram[80][11] , \ram[80][10] , \ram[80][9] ,
         \ram[80][8] , \ram[80][7] , \ram[80][6] , \ram[80][5] , \ram[80][4] ,
         \ram[80][3] , \ram[80][2] , \ram[80][1] , \ram[80][0] , \ram[79][15] ,
         \ram[79][14] , \ram[79][13] , \ram[79][12] , \ram[79][11] ,
         \ram[79][10] , \ram[79][9] , \ram[79][8] , \ram[79][7] , \ram[79][6] ,
         \ram[79][5] , \ram[79][4] , \ram[79][3] , \ram[79][2] , \ram[79][1] ,
         \ram[79][0] , \ram[78][15] , \ram[78][14] , \ram[78][13] ,
         \ram[78][12] , \ram[78][11] , \ram[78][10] , \ram[78][9] ,
         \ram[78][8] , \ram[78][7] , \ram[78][6] , \ram[78][5] , \ram[78][4] ,
         \ram[78][3] , \ram[78][2] , \ram[78][1] , \ram[78][0] , \ram[77][15] ,
         \ram[77][14] , \ram[77][13] , \ram[77][12] , \ram[77][11] ,
         \ram[77][10] , \ram[77][9] , \ram[77][8] , \ram[77][7] , \ram[77][6] ,
         \ram[77][5] , \ram[77][4] , \ram[77][3] , \ram[77][2] , \ram[77][1] ,
         \ram[77][0] , \ram[76][15] , \ram[76][14] , \ram[76][13] ,
         \ram[76][12] , \ram[76][11] , \ram[76][10] , \ram[76][9] ,
         \ram[76][8] , \ram[76][7] , \ram[76][6] , \ram[76][5] , \ram[76][4] ,
         \ram[76][3] , \ram[76][2] , \ram[76][1] , \ram[76][0] , \ram[75][15] ,
         \ram[75][14] , \ram[75][13] , \ram[75][12] , \ram[75][11] ,
         \ram[75][10] , \ram[75][9] , \ram[75][8] , \ram[75][7] , \ram[75][6] ,
         \ram[75][5] , \ram[75][4] , \ram[75][3] , \ram[75][2] , \ram[75][1] ,
         \ram[75][0] , \ram[74][15] , \ram[74][14] , \ram[74][13] ,
         \ram[74][12] , \ram[74][11] , \ram[74][10] , \ram[74][9] ,
         \ram[74][8] , \ram[74][7] , \ram[74][6] , \ram[74][5] , \ram[74][4] ,
         \ram[74][3] , \ram[74][2] , \ram[74][1] , \ram[74][0] , \ram[73][15] ,
         \ram[73][14] , \ram[73][13] , \ram[73][12] , \ram[73][11] ,
         \ram[73][10] , \ram[73][9] , \ram[73][8] , \ram[73][7] , \ram[73][6] ,
         \ram[73][5] , \ram[73][4] , \ram[73][3] , \ram[73][2] , \ram[73][1] ,
         \ram[73][0] , \ram[72][15] , \ram[72][14] , \ram[72][13] ,
         \ram[72][12] , \ram[72][11] , \ram[72][10] , \ram[72][9] ,
         \ram[72][8] , \ram[72][7] , \ram[72][6] , \ram[72][5] , \ram[72][4] ,
         \ram[72][3] , \ram[72][2] , \ram[72][1] , \ram[72][0] , \ram[71][15] ,
         \ram[71][14] , \ram[71][13] , \ram[71][12] , \ram[71][11] ,
         \ram[71][10] , \ram[71][9] , \ram[71][8] , \ram[71][7] , \ram[71][6] ,
         \ram[71][5] , \ram[71][4] , \ram[71][3] , \ram[71][2] , \ram[71][1] ,
         \ram[71][0] , \ram[70][15] , \ram[70][14] , \ram[70][13] ,
         \ram[70][12] , \ram[70][11] , \ram[70][10] , \ram[70][9] ,
         \ram[70][8] , \ram[70][7] , \ram[70][6] , \ram[70][5] , \ram[70][4] ,
         \ram[70][3] , \ram[70][2] , \ram[70][1] , \ram[70][0] , \ram[69][15] ,
         \ram[69][14] , \ram[69][13] , \ram[69][12] , \ram[69][11] ,
         \ram[69][10] , \ram[69][9] , \ram[69][8] , \ram[69][7] , \ram[69][6] ,
         \ram[69][5] , \ram[69][4] , \ram[69][3] , \ram[69][2] , \ram[69][1] ,
         \ram[69][0] , \ram[68][15] , \ram[68][14] , \ram[68][13] ,
         \ram[68][12] , \ram[68][11] , \ram[68][10] , \ram[68][9] ,
         \ram[68][8] , \ram[68][7] , \ram[68][6] , \ram[68][5] , \ram[68][4] ,
         \ram[68][3] , \ram[68][2] , \ram[68][1] , \ram[68][0] , \ram[67][15] ,
         \ram[67][14] , \ram[67][13] , \ram[67][12] , \ram[67][11] ,
         \ram[67][10] , \ram[67][9] , \ram[67][8] , \ram[67][7] , \ram[67][6] ,
         \ram[67][5] , \ram[67][4] , \ram[67][3] , \ram[67][2] , \ram[67][1] ,
         \ram[67][0] , \ram[66][15] , \ram[66][14] , \ram[66][13] ,
         \ram[66][12] , \ram[66][11] , \ram[66][10] , \ram[66][9] ,
         \ram[66][8] , \ram[66][7] , \ram[66][6] , \ram[66][5] , \ram[66][4] ,
         \ram[66][3] , \ram[66][2] , \ram[66][1] , \ram[66][0] , \ram[65][15] ,
         \ram[65][14] , \ram[65][13] , \ram[65][12] , \ram[65][11] ,
         \ram[65][10] , \ram[65][9] , \ram[65][8] , \ram[65][7] , \ram[65][6] ,
         \ram[65][5] , \ram[65][4] , \ram[65][3] , \ram[65][2] , \ram[65][1] ,
         \ram[65][0] , \ram[64][15] , \ram[64][14] , \ram[64][13] ,
         \ram[64][12] , \ram[64][11] , \ram[64][10] , \ram[64][9] ,
         \ram[64][8] , \ram[64][7] , \ram[64][6] , \ram[64][5] , \ram[64][4] ,
         \ram[64][3] , \ram[64][2] , \ram[64][1] , \ram[64][0] , \ram[63][15] ,
         \ram[63][14] , \ram[63][13] , \ram[63][12] , \ram[63][11] ,
         \ram[63][10] , \ram[63][9] , \ram[63][8] , \ram[63][7] , \ram[63][6] ,
         \ram[63][5] , \ram[63][4] , \ram[63][3] , \ram[63][2] , \ram[63][1] ,
         \ram[63][0] , \ram[62][15] , \ram[62][14] , \ram[62][13] ,
         \ram[62][12] , \ram[62][11] , \ram[62][10] , \ram[62][9] ,
         \ram[62][8] , \ram[62][7] , \ram[62][6] , \ram[62][5] , \ram[62][4] ,
         \ram[62][3] , \ram[62][2] , \ram[62][1] , \ram[62][0] , \ram[61][15] ,
         \ram[61][14] , \ram[61][13] , \ram[61][12] , \ram[61][11] ,
         \ram[61][10] , \ram[61][9] , \ram[61][8] , \ram[61][7] , \ram[61][6] ,
         \ram[61][5] , \ram[61][4] , \ram[61][3] , \ram[61][2] , \ram[61][1] ,
         \ram[61][0] , \ram[60][15] , \ram[60][14] , \ram[60][13] ,
         \ram[60][12] , \ram[60][11] , \ram[60][10] , \ram[60][9] ,
         \ram[60][8] , \ram[60][7] , \ram[60][6] , \ram[60][5] , \ram[60][4] ,
         \ram[60][3] , \ram[60][2] , \ram[60][1] , \ram[60][0] , \ram[59][15] ,
         \ram[59][14] , \ram[59][13] , \ram[59][12] , \ram[59][11] ,
         \ram[59][10] , \ram[59][9] , \ram[59][8] , \ram[59][7] , \ram[59][6] ,
         \ram[59][5] , \ram[59][4] , \ram[59][3] , \ram[59][2] , \ram[59][1] ,
         \ram[59][0] , \ram[58][15] , \ram[58][14] , \ram[58][13] ,
         \ram[58][12] , \ram[58][11] , \ram[58][10] , \ram[58][9] ,
         \ram[58][8] , \ram[58][7] , \ram[58][6] , \ram[58][5] , \ram[58][4] ,
         \ram[58][3] , \ram[58][2] , \ram[58][1] , \ram[58][0] , \ram[57][15] ,
         \ram[57][14] , \ram[57][13] , \ram[57][12] , \ram[57][11] ,
         \ram[57][10] , \ram[57][9] , \ram[57][8] , \ram[57][7] , \ram[57][6] ,
         \ram[57][5] , \ram[57][4] , \ram[57][3] , \ram[57][2] , \ram[57][1] ,
         \ram[57][0] , \ram[56][15] , \ram[56][14] , \ram[56][13] ,
         \ram[56][12] , \ram[56][11] , \ram[56][10] , \ram[56][9] ,
         \ram[56][8] , \ram[56][7] , \ram[56][6] , \ram[56][5] , \ram[56][4] ,
         \ram[56][3] , \ram[56][2] , \ram[56][1] , \ram[56][0] , \ram[55][15] ,
         \ram[55][14] , \ram[55][13] , \ram[55][12] , \ram[55][11] ,
         \ram[55][10] , \ram[55][9] , \ram[55][8] , \ram[55][7] , \ram[55][6] ,
         \ram[55][5] , \ram[55][4] , \ram[55][3] , \ram[55][2] , \ram[55][1] ,
         \ram[55][0] , \ram[54][15] , \ram[54][14] , \ram[54][13] ,
         \ram[54][12] , \ram[54][11] , \ram[54][10] , \ram[54][9] ,
         \ram[54][8] , \ram[54][7] , \ram[54][6] , \ram[54][5] , \ram[54][4] ,
         \ram[54][3] , \ram[54][2] , \ram[54][1] , \ram[54][0] , \ram[53][15] ,
         \ram[53][14] , \ram[53][13] , \ram[53][12] , \ram[53][11] ,
         \ram[53][10] , \ram[53][9] , \ram[53][8] , \ram[53][7] , \ram[53][6] ,
         \ram[53][5] , \ram[53][4] , \ram[53][3] , \ram[53][2] , \ram[53][1] ,
         \ram[53][0] , \ram[52][15] , \ram[52][14] , \ram[52][13] ,
         \ram[52][12] , \ram[52][11] , \ram[52][10] , \ram[52][9] ,
         \ram[52][8] , \ram[52][7] , \ram[52][6] , \ram[52][5] , \ram[52][4] ,
         \ram[52][3] , \ram[52][2] , \ram[52][1] , \ram[52][0] , \ram[51][15] ,
         \ram[51][14] , \ram[51][13] , \ram[51][12] , \ram[51][11] ,
         \ram[51][10] , \ram[51][9] , \ram[51][8] , \ram[51][7] , \ram[51][6] ,
         \ram[51][5] , \ram[51][4] , \ram[51][3] , \ram[51][2] , \ram[51][1] ,
         \ram[51][0] , \ram[50][15] , \ram[50][14] , \ram[50][13] ,
         \ram[50][12] , \ram[50][11] , \ram[50][10] , \ram[50][9] ,
         \ram[50][8] , \ram[50][7] , \ram[50][6] , \ram[50][5] , \ram[50][4] ,
         \ram[50][3] , \ram[50][2] , \ram[50][1] , \ram[50][0] , \ram[49][15] ,
         \ram[49][14] , \ram[49][13] , \ram[49][12] , \ram[49][11] ,
         \ram[49][10] , \ram[49][9] , \ram[49][8] , \ram[49][7] , \ram[49][6] ,
         \ram[49][5] , \ram[49][4] , \ram[49][3] , \ram[49][2] , \ram[49][1] ,
         \ram[49][0] , \ram[48][15] , \ram[48][14] , \ram[48][13] ,
         \ram[48][12] , \ram[48][11] , \ram[48][10] , \ram[48][9] ,
         \ram[48][8] , \ram[48][7] , \ram[48][6] , \ram[48][5] , \ram[48][4] ,
         \ram[48][3] , \ram[48][2] , \ram[48][1] , \ram[48][0] , \ram[47][15] ,
         \ram[47][14] , \ram[47][13] , \ram[47][12] , \ram[47][11] ,
         \ram[47][10] , \ram[47][9] , \ram[47][8] , \ram[47][7] , \ram[47][6] ,
         \ram[47][5] , \ram[47][4] , \ram[47][3] , \ram[47][2] , \ram[47][1] ,
         \ram[47][0] , \ram[46][15] , \ram[46][14] , \ram[46][13] ,
         \ram[46][12] , \ram[46][11] , \ram[46][10] , \ram[46][9] ,
         \ram[46][8] , \ram[46][7] , \ram[46][6] , \ram[46][5] , \ram[46][4] ,
         \ram[46][3] , \ram[46][2] , \ram[46][1] , \ram[46][0] , \ram[45][15] ,
         \ram[45][14] , \ram[45][13] , \ram[45][12] , \ram[45][11] ,
         \ram[45][10] , \ram[45][9] , \ram[45][8] , \ram[45][7] , \ram[45][6] ,
         \ram[45][5] , \ram[45][4] , \ram[45][3] , \ram[45][2] , \ram[45][1] ,
         \ram[45][0] , \ram[44][15] , \ram[44][14] , \ram[44][13] ,
         \ram[44][12] , \ram[44][11] , \ram[44][10] , \ram[44][9] ,
         \ram[44][8] , \ram[44][7] , \ram[44][6] , \ram[44][5] , \ram[44][4] ,
         \ram[44][3] , \ram[44][2] , \ram[44][1] , \ram[44][0] , \ram[43][15] ,
         \ram[43][14] , \ram[43][13] , \ram[43][12] , \ram[43][11] ,
         \ram[43][10] , \ram[43][9] , \ram[43][8] , \ram[43][7] , \ram[43][6] ,
         \ram[43][5] , \ram[43][4] , \ram[43][3] , \ram[43][2] , \ram[43][1] ,
         \ram[43][0] , \ram[42][15] , \ram[42][14] , \ram[42][13] ,
         \ram[42][12] , \ram[42][11] , \ram[42][10] , \ram[42][9] ,
         \ram[42][8] , \ram[42][7] , \ram[42][6] , \ram[42][5] , \ram[42][4] ,
         \ram[42][3] , \ram[42][2] , \ram[42][1] , \ram[42][0] , \ram[41][15] ,
         \ram[41][14] , \ram[41][13] , \ram[41][12] , \ram[41][11] ,
         \ram[41][10] , \ram[41][9] , \ram[41][8] , \ram[41][7] , \ram[41][6] ,
         \ram[41][5] , \ram[41][4] , \ram[41][3] , \ram[41][2] , \ram[41][1] ,
         \ram[41][0] , \ram[40][15] , \ram[40][14] , \ram[40][13] ,
         \ram[40][12] , \ram[40][11] , \ram[40][10] , \ram[40][9] ,
         \ram[40][8] , \ram[40][7] , \ram[40][6] , \ram[40][5] , \ram[40][4] ,
         \ram[40][3] , \ram[40][2] , \ram[40][1] , \ram[40][0] , \ram[39][15] ,
         \ram[39][14] , \ram[39][13] , \ram[39][12] , \ram[39][11] ,
         \ram[39][10] , \ram[39][9] , \ram[39][8] , \ram[39][7] , \ram[39][6] ,
         \ram[39][5] , \ram[39][4] , \ram[39][3] , \ram[39][2] , \ram[39][1] ,
         \ram[39][0] , \ram[38][15] , \ram[38][14] , \ram[38][13] ,
         \ram[38][12] , \ram[38][11] , \ram[38][10] , \ram[38][9] ,
         \ram[38][8] , \ram[38][7] , \ram[38][6] , \ram[38][5] , \ram[38][4] ,
         \ram[38][3] , \ram[38][2] , \ram[38][1] , \ram[38][0] , \ram[37][15] ,
         \ram[37][14] , \ram[37][13] , \ram[37][12] , \ram[37][11] ,
         \ram[37][10] , \ram[37][9] , \ram[37][8] , \ram[37][7] , \ram[37][6] ,
         \ram[37][5] , \ram[37][4] , \ram[37][3] , \ram[37][2] , \ram[37][1] ,
         \ram[37][0] , \ram[36][15] , \ram[36][14] , \ram[36][13] ,
         \ram[36][12] , \ram[36][11] , \ram[36][10] , \ram[36][9] ,
         \ram[36][8] , \ram[36][7] , \ram[36][6] , \ram[36][5] , \ram[36][4] ,
         \ram[36][3] , \ram[36][2] , \ram[36][1] , \ram[36][0] , \ram[35][15] ,
         \ram[35][14] , \ram[35][13] , \ram[35][12] , \ram[35][11] ,
         \ram[35][10] , \ram[35][9] , \ram[35][8] , \ram[35][7] , \ram[35][6] ,
         \ram[35][5] , \ram[35][4] , \ram[35][3] , \ram[35][2] , \ram[35][1] ,
         \ram[35][0] , \ram[34][15] , \ram[34][14] , \ram[34][13] ,
         \ram[34][12] , \ram[34][11] , \ram[34][10] , \ram[34][9] ,
         \ram[34][8] , \ram[34][7] , \ram[34][6] , \ram[34][5] , \ram[34][4] ,
         \ram[34][3] , \ram[34][2] , \ram[34][1] , \ram[34][0] , \ram[33][15] ,
         \ram[33][14] , \ram[33][13] , \ram[33][12] , \ram[33][11] ,
         \ram[33][10] , \ram[33][9] , \ram[33][8] , \ram[33][7] , \ram[33][6] ,
         \ram[33][5] , \ram[33][4] , \ram[33][3] , \ram[33][2] , \ram[33][1] ,
         \ram[33][0] , \ram[32][15] , \ram[32][14] , \ram[32][13] ,
         \ram[32][12] , \ram[32][11] , \ram[32][10] , \ram[32][9] ,
         \ram[32][8] , \ram[32][7] , \ram[32][6] , \ram[32][5] , \ram[32][4] ,
         \ram[32][3] , \ram[32][2] , \ram[32][1] , \ram[32][0] , \ram[31][15] ,
         \ram[31][14] , \ram[31][13] , \ram[31][12] , \ram[31][11] ,
         \ram[31][10] , \ram[31][9] , \ram[31][8] , \ram[31][7] , \ram[31][6] ,
         \ram[31][5] , \ram[31][4] , \ram[31][3] , \ram[31][2] , \ram[31][1] ,
         \ram[31][0] , \ram[30][15] , \ram[30][14] , \ram[30][13] ,
         \ram[30][12] , \ram[30][11] , \ram[30][10] , \ram[30][9] ,
         \ram[30][8] , \ram[30][7] , \ram[30][6] , \ram[30][5] , \ram[30][4] ,
         \ram[30][3] , \ram[30][2] , \ram[30][1] , \ram[30][0] , \ram[29][15] ,
         \ram[29][14] , \ram[29][13] , \ram[29][12] , \ram[29][11] ,
         \ram[29][10] , \ram[29][9] , \ram[29][8] , \ram[29][7] , \ram[29][6] ,
         \ram[29][5] , \ram[29][4] , \ram[29][3] , \ram[29][2] , \ram[29][1] ,
         \ram[29][0] , \ram[28][15] , \ram[28][14] , \ram[28][13] ,
         \ram[28][12] , \ram[28][11] , \ram[28][10] , \ram[28][9] ,
         \ram[28][8] , \ram[28][7] , \ram[28][6] , \ram[28][5] , \ram[28][4] ,
         \ram[28][3] , \ram[28][2] , \ram[28][1] , \ram[28][0] , \ram[27][15] ,
         \ram[27][14] , \ram[27][13] , \ram[27][12] , \ram[27][11] ,
         \ram[27][10] , \ram[27][9] , \ram[27][8] , \ram[27][7] , \ram[27][6] ,
         \ram[27][5] , \ram[27][4] , \ram[27][3] , \ram[27][2] , \ram[27][1] ,
         \ram[27][0] , \ram[26][15] , \ram[26][14] , \ram[26][13] ,
         \ram[26][12] , \ram[26][11] , \ram[26][10] , \ram[26][9] ,
         \ram[26][8] , \ram[26][7] , \ram[26][6] , \ram[26][5] , \ram[26][4] ,
         \ram[26][3] , \ram[26][2] , \ram[26][1] , \ram[26][0] , \ram[25][15] ,
         \ram[25][14] , \ram[25][13] , \ram[25][12] , \ram[25][11] ,
         \ram[25][10] , \ram[25][9] , \ram[25][8] , \ram[25][7] , \ram[25][6] ,
         \ram[25][5] , \ram[25][4] , \ram[25][3] , \ram[25][2] , \ram[25][1] ,
         \ram[25][0] , \ram[24][15] , \ram[24][14] , \ram[24][13] ,
         \ram[24][12] , \ram[24][11] , \ram[24][10] , \ram[24][9] ,
         \ram[24][8] , \ram[24][7] , \ram[24][6] , \ram[24][5] , \ram[24][4] ,
         \ram[24][3] , \ram[24][2] , \ram[24][1] , \ram[24][0] , \ram[23][15] ,
         \ram[23][14] , \ram[23][13] , \ram[23][12] , \ram[23][11] ,
         \ram[23][10] , \ram[23][9] , \ram[23][8] , \ram[23][7] , \ram[23][6] ,
         \ram[23][5] , \ram[23][4] , \ram[23][3] , \ram[23][2] , \ram[23][1] ,
         \ram[23][0] , \ram[22][15] , \ram[22][14] , \ram[22][13] ,
         \ram[22][12] , \ram[22][11] , \ram[22][10] , \ram[22][9] ,
         \ram[22][8] , \ram[22][7] , \ram[22][6] , \ram[22][5] , \ram[22][4] ,
         \ram[22][3] , \ram[22][2] , \ram[22][1] , \ram[22][0] , \ram[21][15] ,
         \ram[21][14] , \ram[21][13] , \ram[21][12] , \ram[21][11] ,
         \ram[21][10] , \ram[21][9] , \ram[21][8] , \ram[21][7] , \ram[21][6] ,
         \ram[21][5] , \ram[21][4] , \ram[21][3] , \ram[21][2] , \ram[21][1] ,
         \ram[21][0] , \ram[20][15] , \ram[20][14] , \ram[20][13] ,
         \ram[20][12] , \ram[20][11] , \ram[20][10] , \ram[20][9] ,
         \ram[20][8] , \ram[20][7] , \ram[20][6] , \ram[20][5] , \ram[20][4] ,
         \ram[20][3] , \ram[20][2] , \ram[20][1] , \ram[20][0] , \ram[19][15] ,
         \ram[19][14] , \ram[19][13] , \ram[19][12] , \ram[19][11] ,
         \ram[19][10] , \ram[19][9] , \ram[19][8] , \ram[19][7] , \ram[19][6] ,
         \ram[19][5] , \ram[19][4] , \ram[19][3] , \ram[19][2] , \ram[19][1] ,
         \ram[19][0] , \ram[18][15] , \ram[18][14] , \ram[18][13] ,
         \ram[18][12] , \ram[18][11] , \ram[18][10] , \ram[18][9] ,
         \ram[18][8] , \ram[18][7] , \ram[18][6] , \ram[18][5] , \ram[18][4] ,
         \ram[18][3] , \ram[18][2] , \ram[18][1] , \ram[18][0] , \ram[17][15] ,
         \ram[17][14] , \ram[17][13] , \ram[17][12] , \ram[17][11] ,
         \ram[17][10] , \ram[17][9] , \ram[17][8] , \ram[17][7] , \ram[17][6] ,
         \ram[17][5] , \ram[17][4] , \ram[17][3] , \ram[17][2] , \ram[17][1] ,
         \ram[17][0] , \ram[16][15] , \ram[16][14] , \ram[16][13] ,
         \ram[16][12] , \ram[16][11] , \ram[16][10] , \ram[16][9] ,
         \ram[16][8] , \ram[16][7] , \ram[16][6] , \ram[16][5] , \ram[16][4] ,
         \ram[16][3] , \ram[16][2] , \ram[16][1] , \ram[16][0] , \ram[15][15] ,
         \ram[15][14] , \ram[15][13] , \ram[15][12] , \ram[15][11] ,
         \ram[15][10] , \ram[15][9] , \ram[15][8] , \ram[15][7] , \ram[15][6] ,
         \ram[15][5] , \ram[15][4] , \ram[15][3] , \ram[15][2] , \ram[15][1] ,
         \ram[15][0] , \ram[14][15] , \ram[14][14] , \ram[14][13] ,
         \ram[14][12] , \ram[14][11] , \ram[14][10] , \ram[14][9] ,
         \ram[14][8] , \ram[14][7] , \ram[14][6] , \ram[14][5] , \ram[14][4] ,
         \ram[14][3] , \ram[14][2] , \ram[14][1] , \ram[14][0] , \ram[13][15] ,
         \ram[13][14] , \ram[13][13] , \ram[13][12] , \ram[13][11] ,
         \ram[13][10] , \ram[13][9] , \ram[13][8] , \ram[13][7] , \ram[13][6] ,
         \ram[13][5] , \ram[13][4] , \ram[13][3] , \ram[13][2] , \ram[13][1] ,
         \ram[13][0] , \ram[12][15] , \ram[12][14] , \ram[12][13] ,
         \ram[12][12] , \ram[12][11] , \ram[12][10] , \ram[12][9] ,
         \ram[12][8] , \ram[12][7] , \ram[12][6] , \ram[12][5] , \ram[12][4] ,
         \ram[12][3] , \ram[12][2] , \ram[12][1] , \ram[12][0] , \ram[11][15] ,
         \ram[11][14] , \ram[11][13] , \ram[11][12] , \ram[11][11] ,
         \ram[11][10] , \ram[11][9] , \ram[11][8] , \ram[11][7] , \ram[11][6] ,
         \ram[11][5] , \ram[11][4] , \ram[11][3] , \ram[11][2] , \ram[11][1] ,
         \ram[11][0] , \ram[10][15] , \ram[10][14] , \ram[10][13] ,
         \ram[10][12] , \ram[10][11] , \ram[10][10] , \ram[10][9] ,
         \ram[10][8] , \ram[10][7] , \ram[10][6] , \ram[10][5] , \ram[10][4] ,
         \ram[10][3] , \ram[10][2] , \ram[10][1] , \ram[10][0] , \ram[9][15] ,
         \ram[9][14] , \ram[9][13] , \ram[9][12] , \ram[9][11] , \ram[9][10] ,
         \ram[9][9] , \ram[9][8] , \ram[9][7] , \ram[9][6] , \ram[9][5] ,
         \ram[9][4] , \ram[9][3] , \ram[9][2] , \ram[9][1] , \ram[9][0] ,
         \ram[8][15] , \ram[8][14] , \ram[8][13] , \ram[8][12] , \ram[8][11] ,
         \ram[8][10] , \ram[8][9] , \ram[8][8] , \ram[8][7] , \ram[8][6] ,
         \ram[8][5] , \ram[8][4] , \ram[8][3] , \ram[8][2] , \ram[8][1] ,
         \ram[8][0] , \ram[7][15] , \ram[7][14] , \ram[7][13] , \ram[7][12] ,
         \ram[7][11] , \ram[7][10] , \ram[7][9] , \ram[7][8] , \ram[7][7] ,
         \ram[7][6] , \ram[7][5] , \ram[7][4] , \ram[7][3] , \ram[7][2] ,
         \ram[7][1] , \ram[7][0] , \ram[6][15] , \ram[6][14] , \ram[6][13] ,
         \ram[6][12] , \ram[6][11] , \ram[6][10] , \ram[6][9] , \ram[6][8] ,
         \ram[6][7] , \ram[6][6] , \ram[6][5] , \ram[6][4] , \ram[6][3] ,
         \ram[6][2] , \ram[6][1] , \ram[6][0] , \ram[5][15] , \ram[5][14] ,
         \ram[5][13] , \ram[5][12] , \ram[5][11] , \ram[5][10] , \ram[5][9] ,
         \ram[5][8] , \ram[5][7] , \ram[5][6] , \ram[5][5] , \ram[5][4] ,
         \ram[5][3] , \ram[5][2] , \ram[5][1] , \ram[5][0] , \ram[4][15] ,
         \ram[4][14] , \ram[4][13] , \ram[4][12] , \ram[4][11] , \ram[4][10] ,
         \ram[4][9] , \ram[4][8] , \ram[4][7] , \ram[4][6] , \ram[4][5] ,
         \ram[4][4] , \ram[4][3] , \ram[4][2] , \ram[4][1] , \ram[4][0] ,
         \ram[3][15] , \ram[3][14] , \ram[3][13] , \ram[3][12] , \ram[3][11] ,
         \ram[3][10] , \ram[3][9] , \ram[3][8] , \ram[3][7] , \ram[3][6] ,
         \ram[3][5] , \ram[3][4] , \ram[3][3] , \ram[3][2] , \ram[3][1] ,
         \ram[3][0] , \ram[2][15] , \ram[2][14] , \ram[2][13] , \ram[2][12] ,
         \ram[2][11] , \ram[2][10] , \ram[2][9] , \ram[2][8] , \ram[2][7] ,
         \ram[2][6] , \ram[2][5] , \ram[2][4] , \ram[2][3] , \ram[2][2] ,
         \ram[2][1] , \ram[2][0] , \ram[1][15] , \ram[1][14] , \ram[1][13] ,
         \ram[1][12] , \ram[1][11] , \ram[1][10] , \ram[1][9] , \ram[1][8] ,
         \ram[1][7] , \ram[1][6] , \ram[1][5] , \ram[1][4] , \ram[1][3] ,
         \ram[1][2] , \ram[1][1] , \ram[1][0] , \ram[0][15] , \ram[0][14] ,
         \ram[0][13] , \ram[0][12] , \ram[0][11] , \ram[0][10] , \ram[0][9] ,
         \ram[0][8] , \ram[0][7] , \ram[0][6] , \ram[0][5] , \ram[0][4] ,
         \ram[0][3] , \ram[0][2] , \ram[0][1] , \ram[0][0] , n7, n8, n9, n10,
         n11, n27, n30, n33, n36, n39, n42, n45, n48, n51, n54, n57, n60, n63,
         n66, n69, n71, n72, n74, n77, n79, n81, n83, n85, n87, n89, n91, n93,
         n95, n97, n99, n101, n103, n105, n106, n108, n111, n113, n115, n117,
         n119, n121, n123, n125, n127, n129, n131, n133, n135, n137, n139,
         n140, n142, n145, n147, n149, n151, n153, n155, n157, n159, n161,
         n163, n165, n167, n169, n171, n173, n174, n176, n179, n181, n183,
         n185, n187, n189, n191, n193, n195, n197, n199, n201, n203, n205,
         n207, n208, n210, n213, n215, n217, n219, n221, n223, n225, n227,
         n229, n231, n233, n235, n237, n239, n241, n243, n246, n248, n250,
         n252, n254, n256, n258, n260, n262, n264, n266, n268, n270, n272,
         n274, n276, n279, n281, n283, n285, n287, n289, n291, n293, n295,
         n297, n299, n301, n303, n305, n307, n309, n312, n314, n316, n318,
         n320, n322, n324, n326, n328, n330, n332, n334, n336, n338, n340,
         n341, n343, n346, n348, n350, n352, n354, n356, n358, n360, n362,
         n364, n366, n368, n370, n372, n374, n376, n379, n381, n383, n385,
         n387, n389, n391, n393, n395, n397, n399, n401, n403, n405, n407,
         n409, n412, n414, n416, n418, n420, n422, n424, n426, n428, n430,
         n432, n434, n436, n438, n440, n442, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n474,
         n476, n479, n481, n483, n485, n487, n489, n491, n493, n495, n497,
         n499, n501, n503, n505, n507, n509, n512, n514, n516, n518, n520,
         n522, n524, n526, n528, n530, n532, n534, n536, n538, n540, n542,
         n544, n545, n547, n548, n550, n551, n553, n554, n556, n557, n559,
         n561, n563, n565, n566, n568, n570, n572, n574, n575, n577, n579,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n1, n2,
         n3, n4, n5, n6, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n28, n29, n31, n32, n34, n35, n37, n38, n40, n41,
         n43, n44, n46, n47, n49, n50, n52, n53, n55, n56, n58, n59, n61, n62,
         n64, n65, n67, n68, n70, n73, n75, n76, n78, n80, n82, n84, n86, n88,
         n90, n92, n94, n96, n98, n100, n102, n104, n107, n109, n110, n112,
         n114, n116, n118, n120, n122, n124, n126, n128, n130, n132, n134,
         n136, n138, n141, n143, n144, n146, n148, n150, n152, n154, n156,
         n158, n160, n162, n164, n166, n168, n170, n172, n175, n177, n178,
         n180, n182, n184, n186, n188, n190, n192, n194, n196, n198, n200,
         n202, n204, n206, n209, n211, n212, n214, n216, n218, n220, n222,
         n224, n226, n228, n230, n232, n234, n236, n238, n240, n242, n244,
         n245, n247, n249, n251, n253, n255, n257, n259, n261, n263, n265,
         n267, n269, n271, n273, n275, n277, n278, n280, n282, n284, n286,
         n288, n290, n292, n294, n296, n298, n300, n302, n304, n306, n308,
         n310, n311, n313, n315, n317, n319, n321, n323, n325, n327, n329,
         n331, n333, n335, n337, n339, n342, n344, n345, n347, n349, n351,
         n353, n355, n357, n359, n361, n363, n365, n367, n369, n371, n373,
         n375, n377, n378, n380, n382, n384, n386, n388, n390, n392, n394,
         n396, n398, n400, n402, n404, n406, n408, n410, n411, n413, n415,
         n417, n419, n421, n423, n425, n427, n429, n431, n433, n435, n437,
         n439, n441, n443, n444, n446, n448, n450, n452, n454, n456, n458,
         n460, n462, n464, n466, n468, n470, n472, n475, n477, n478, n480,
         n482, n484, n486, n488, n490, n492, n494, n496, n498, n500, n502,
         n504, n506, n508, n510, n511, n513, n515, n517, n519, n521, n523,
         n525, n527, n529, n531, n533, n535, n537, n539, n541, n543, n546,
         n549, n552, n555, n558, n560, n562, n564, n567, n569, n571, n573,
         n576, n578, n580, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017;
  assign N18 = mem_access_addr[0];
  assign N19 = mem_access_addr[1];
  assign N20 = mem_access_addr[2];
  assign N21 = mem_access_addr[3];
  assign N22 = mem_access_addr[4];
  assign N23 = mem_access_addr[5];
  assign N24 = mem_access_addr[6];
  assign N25 = mem_access_addr[7];

  DFFHQX1 \ram_reg[253][15]  ( .D(n4645), .CK(clk), .Q(\ram[253][15] ) );
  DFFHQX1 \ram_reg[253][14]  ( .D(n4644), .CK(clk), .Q(\ram[253][14] ) );
  DFFHQX1 \ram_reg[253][13]  ( .D(n4643), .CK(clk), .Q(\ram[253][13] ) );
  DFFHQX1 \ram_reg[253][12]  ( .D(n4642), .CK(clk), .Q(\ram[253][12] ) );
  DFFHQX1 \ram_reg[253][11]  ( .D(n4641), .CK(clk), .Q(\ram[253][11] ) );
  DFFHQX1 \ram_reg[253][10]  ( .D(n4640), .CK(clk), .Q(\ram[253][10] ) );
  DFFHQX1 \ram_reg[253][9]  ( .D(n4639), .CK(clk), .Q(\ram[253][9] ) );
  DFFHQX1 \ram_reg[253][8]  ( .D(n4638), .CK(clk), .Q(\ram[253][8] ) );
  DFFHQX1 \ram_reg[253][7]  ( .D(n4637), .CK(clk), .Q(\ram[253][7] ) );
  DFFHQX1 \ram_reg[253][6]  ( .D(n4636), .CK(clk), .Q(\ram[253][6] ) );
  DFFHQX1 \ram_reg[253][5]  ( .D(n4635), .CK(clk), .Q(\ram[253][5] ) );
  DFFHQX1 \ram_reg[253][4]  ( .D(n4634), .CK(clk), .Q(\ram[253][4] ) );
  DFFHQX1 \ram_reg[253][3]  ( .D(n4633), .CK(clk), .Q(\ram[253][3] ) );
  DFFHQX1 \ram_reg[253][2]  ( .D(n4632), .CK(clk), .Q(\ram[253][2] ) );
  DFFHQX1 \ram_reg[253][1]  ( .D(n4631), .CK(clk), .Q(\ram[253][1] ) );
  DFFHQX1 \ram_reg[253][0]  ( .D(n4630), .CK(clk), .Q(\ram[253][0] ) );
  DFFHQX1 \ram_reg[249][15]  ( .D(n4581), .CK(clk), .Q(\ram[249][15] ) );
  DFFHQX1 \ram_reg[249][14]  ( .D(n4580), .CK(clk), .Q(\ram[249][14] ) );
  DFFHQX1 \ram_reg[249][13]  ( .D(n4579), .CK(clk), .Q(\ram[249][13] ) );
  DFFHQX1 \ram_reg[249][12]  ( .D(n4578), .CK(clk), .Q(\ram[249][12] ) );
  DFFHQX1 \ram_reg[249][11]  ( .D(n4577), .CK(clk), .Q(\ram[249][11] ) );
  DFFHQX1 \ram_reg[249][10]  ( .D(n4576), .CK(clk), .Q(\ram[249][10] ) );
  DFFHQX1 \ram_reg[249][9]  ( .D(n4575), .CK(clk), .Q(\ram[249][9] ) );
  DFFHQX1 \ram_reg[249][8]  ( .D(n4574), .CK(clk), .Q(\ram[249][8] ) );
  DFFHQX1 \ram_reg[249][7]  ( .D(n4573), .CK(clk), .Q(\ram[249][7] ) );
  DFFHQX1 \ram_reg[249][6]  ( .D(n4572), .CK(clk), .Q(\ram[249][6] ) );
  DFFHQX1 \ram_reg[249][5]  ( .D(n4571), .CK(clk), .Q(\ram[249][5] ) );
  DFFHQX1 \ram_reg[249][4]  ( .D(n4570), .CK(clk), .Q(\ram[249][4] ) );
  DFFHQX1 \ram_reg[249][3]  ( .D(n4569), .CK(clk), .Q(\ram[249][3] ) );
  DFFHQX1 \ram_reg[249][2]  ( .D(n4568), .CK(clk), .Q(\ram[249][2] ) );
  DFFHQX1 \ram_reg[249][1]  ( .D(n4567), .CK(clk), .Q(\ram[249][1] ) );
  DFFHQX1 \ram_reg[249][0]  ( .D(n4566), .CK(clk), .Q(\ram[249][0] ) );
  DFFHQX1 \ram_reg[245][15]  ( .D(n4517), .CK(clk), .Q(\ram[245][15] ) );
  DFFHQX1 \ram_reg[245][14]  ( .D(n4516), .CK(clk), .Q(\ram[245][14] ) );
  DFFHQX1 \ram_reg[245][13]  ( .D(n4515), .CK(clk), .Q(\ram[245][13] ) );
  DFFHQX1 \ram_reg[245][12]  ( .D(n4514), .CK(clk), .Q(\ram[245][12] ) );
  DFFHQX1 \ram_reg[245][11]  ( .D(n4513), .CK(clk), .Q(\ram[245][11] ) );
  DFFHQX1 \ram_reg[245][10]  ( .D(n4512), .CK(clk), .Q(\ram[245][10] ) );
  DFFHQX1 \ram_reg[245][9]  ( .D(n4511), .CK(clk), .Q(\ram[245][9] ) );
  DFFHQX1 \ram_reg[245][8]  ( .D(n4510), .CK(clk), .Q(\ram[245][8] ) );
  DFFHQX1 \ram_reg[245][7]  ( .D(n4509), .CK(clk), .Q(\ram[245][7] ) );
  DFFHQX1 \ram_reg[245][6]  ( .D(n4508), .CK(clk), .Q(\ram[245][6] ) );
  DFFHQX1 \ram_reg[245][5]  ( .D(n4507), .CK(clk), .Q(\ram[245][5] ) );
  DFFHQX1 \ram_reg[245][4]  ( .D(n4506), .CK(clk), .Q(\ram[245][4] ) );
  DFFHQX1 \ram_reg[245][3]  ( .D(n4505), .CK(clk), .Q(\ram[245][3] ) );
  DFFHQX1 \ram_reg[245][2]  ( .D(n4504), .CK(clk), .Q(\ram[245][2] ) );
  DFFHQX1 \ram_reg[245][1]  ( .D(n4503), .CK(clk), .Q(\ram[245][1] ) );
  DFFHQX1 \ram_reg[245][0]  ( .D(n4502), .CK(clk), .Q(\ram[245][0] ) );
  DFFHQX1 \ram_reg[241][15]  ( .D(n4453), .CK(clk), .Q(\ram[241][15] ) );
  DFFHQX1 \ram_reg[241][14]  ( .D(n4452), .CK(clk), .Q(\ram[241][14] ) );
  DFFHQX1 \ram_reg[241][13]  ( .D(n4451), .CK(clk), .Q(\ram[241][13] ) );
  DFFHQX1 \ram_reg[241][12]  ( .D(n4450), .CK(clk), .Q(\ram[241][12] ) );
  DFFHQX1 \ram_reg[241][11]  ( .D(n4449), .CK(clk), .Q(\ram[241][11] ) );
  DFFHQX1 \ram_reg[241][10]  ( .D(n4448), .CK(clk), .Q(\ram[241][10] ) );
  DFFHQX1 \ram_reg[241][9]  ( .D(n4447), .CK(clk), .Q(\ram[241][9] ) );
  DFFHQX1 \ram_reg[241][8]  ( .D(n4446), .CK(clk), .Q(\ram[241][8] ) );
  DFFHQX1 \ram_reg[241][7]  ( .D(n4445), .CK(clk), .Q(\ram[241][7] ) );
  DFFHQX1 \ram_reg[241][6]  ( .D(n4444), .CK(clk), .Q(\ram[241][6] ) );
  DFFHQX1 \ram_reg[241][5]  ( .D(n4443), .CK(clk), .Q(\ram[241][5] ) );
  DFFHQX1 \ram_reg[241][4]  ( .D(n4442), .CK(clk), .Q(\ram[241][4] ) );
  DFFHQX1 \ram_reg[241][3]  ( .D(n4441), .CK(clk), .Q(\ram[241][3] ) );
  DFFHQX1 \ram_reg[241][2]  ( .D(n4440), .CK(clk), .Q(\ram[241][2] ) );
  DFFHQX1 \ram_reg[241][1]  ( .D(n4439), .CK(clk), .Q(\ram[241][1] ) );
  DFFHQX1 \ram_reg[241][0]  ( .D(n4438), .CK(clk), .Q(\ram[241][0] ) );
  DFFHQX1 \ram_reg[237][15]  ( .D(n4389), .CK(clk), .Q(\ram[237][15] ) );
  DFFHQX1 \ram_reg[237][14]  ( .D(n4388), .CK(clk), .Q(\ram[237][14] ) );
  DFFHQX1 \ram_reg[237][13]  ( .D(n4387), .CK(clk), .Q(\ram[237][13] ) );
  DFFHQX1 \ram_reg[237][12]  ( .D(n4386), .CK(clk), .Q(\ram[237][12] ) );
  DFFHQX1 \ram_reg[237][11]  ( .D(n4385), .CK(clk), .Q(\ram[237][11] ) );
  DFFHQX1 \ram_reg[237][10]  ( .D(n4384), .CK(clk), .Q(\ram[237][10] ) );
  DFFHQX1 \ram_reg[237][9]  ( .D(n4383), .CK(clk), .Q(\ram[237][9] ) );
  DFFHQX1 \ram_reg[237][8]  ( .D(n4382), .CK(clk), .Q(\ram[237][8] ) );
  DFFHQX1 \ram_reg[237][7]  ( .D(n4381), .CK(clk), .Q(\ram[237][7] ) );
  DFFHQX1 \ram_reg[237][6]  ( .D(n4380), .CK(clk), .Q(\ram[237][6] ) );
  DFFHQX1 \ram_reg[237][5]  ( .D(n4379), .CK(clk), .Q(\ram[237][5] ) );
  DFFHQX1 \ram_reg[237][4]  ( .D(n4378), .CK(clk), .Q(\ram[237][4] ) );
  DFFHQX1 \ram_reg[237][3]  ( .D(n4377), .CK(clk), .Q(\ram[237][3] ) );
  DFFHQX1 \ram_reg[237][2]  ( .D(n4376), .CK(clk), .Q(\ram[237][2] ) );
  DFFHQX1 \ram_reg[237][1]  ( .D(n4375), .CK(clk), .Q(\ram[237][1] ) );
  DFFHQX1 \ram_reg[237][0]  ( .D(n4374), .CK(clk), .Q(\ram[237][0] ) );
  DFFHQX1 \ram_reg[233][15]  ( .D(n4325), .CK(clk), .Q(\ram[233][15] ) );
  DFFHQX1 \ram_reg[233][14]  ( .D(n4324), .CK(clk), .Q(\ram[233][14] ) );
  DFFHQX1 \ram_reg[233][13]  ( .D(n4323), .CK(clk), .Q(\ram[233][13] ) );
  DFFHQX1 \ram_reg[233][12]  ( .D(n4322), .CK(clk), .Q(\ram[233][12] ) );
  DFFHQX1 \ram_reg[233][11]  ( .D(n4321), .CK(clk), .Q(\ram[233][11] ) );
  DFFHQX1 \ram_reg[233][10]  ( .D(n4320), .CK(clk), .Q(\ram[233][10] ) );
  DFFHQX1 \ram_reg[233][9]  ( .D(n4319), .CK(clk), .Q(\ram[233][9] ) );
  DFFHQX1 \ram_reg[233][8]  ( .D(n4318), .CK(clk), .Q(\ram[233][8] ) );
  DFFHQX1 \ram_reg[233][7]  ( .D(n4317), .CK(clk), .Q(\ram[233][7] ) );
  DFFHQX1 \ram_reg[233][6]  ( .D(n4316), .CK(clk), .Q(\ram[233][6] ) );
  DFFHQX1 \ram_reg[233][5]  ( .D(n4315), .CK(clk), .Q(\ram[233][5] ) );
  DFFHQX1 \ram_reg[233][4]  ( .D(n4314), .CK(clk), .Q(\ram[233][4] ) );
  DFFHQX1 \ram_reg[233][3]  ( .D(n4313), .CK(clk), .Q(\ram[233][3] ) );
  DFFHQX1 \ram_reg[233][2]  ( .D(n4312), .CK(clk), .Q(\ram[233][2] ) );
  DFFHQX1 \ram_reg[233][1]  ( .D(n4311), .CK(clk), .Q(\ram[233][1] ) );
  DFFHQX1 \ram_reg[233][0]  ( .D(n4310), .CK(clk), .Q(\ram[233][0] ) );
  DFFHQX1 \ram_reg[229][15]  ( .D(n4261), .CK(clk), .Q(\ram[229][15] ) );
  DFFHQX1 \ram_reg[229][14]  ( .D(n4260), .CK(clk), .Q(\ram[229][14] ) );
  DFFHQX1 \ram_reg[229][13]  ( .D(n4259), .CK(clk), .Q(\ram[229][13] ) );
  DFFHQX1 \ram_reg[229][12]  ( .D(n4258), .CK(clk), .Q(\ram[229][12] ) );
  DFFHQX1 \ram_reg[229][11]  ( .D(n4257), .CK(clk), .Q(\ram[229][11] ) );
  DFFHQX1 \ram_reg[229][10]  ( .D(n4256), .CK(clk), .Q(\ram[229][10] ) );
  DFFHQX1 \ram_reg[229][9]  ( .D(n4255), .CK(clk), .Q(\ram[229][9] ) );
  DFFHQX1 \ram_reg[229][8]  ( .D(n4254), .CK(clk), .Q(\ram[229][8] ) );
  DFFHQX1 \ram_reg[229][7]  ( .D(n4253), .CK(clk), .Q(\ram[229][7] ) );
  DFFHQX1 \ram_reg[229][6]  ( .D(n4252), .CK(clk), .Q(\ram[229][6] ) );
  DFFHQX1 \ram_reg[229][5]  ( .D(n4251), .CK(clk), .Q(\ram[229][5] ) );
  DFFHQX1 \ram_reg[229][4]  ( .D(n4250), .CK(clk), .Q(\ram[229][4] ) );
  DFFHQX1 \ram_reg[229][3]  ( .D(n4249), .CK(clk), .Q(\ram[229][3] ) );
  DFFHQX1 \ram_reg[229][2]  ( .D(n4248), .CK(clk), .Q(\ram[229][2] ) );
  DFFHQX1 \ram_reg[229][1]  ( .D(n4247), .CK(clk), .Q(\ram[229][1] ) );
  DFFHQX1 \ram_reg[229][0]  ( .D(n4246), .CK(clk), .Q(\ram[229][0] ) );
  DFFHQX1 \ram_reg[225][15]  ( .D(n4197), .CK(clk), .Q(\ram[225][15] ) );
  DFFHQX1 \ram_reg[225][14]  ( .D(n4196), .CK(clk), .Q(\ram[225][14] ) );
  DFFHQX1 \ram_reg[225][13]  ( .D(n4195), .CK(clk), .Q(\ram[225][13] ) );
  DFFHQX1 \ram_reg[225][12]  ( .D(n4194), .CK(clk), .Q(\ram[225][12] ) );
  DFFHQX1 \ram_reg[225][11]  ( .D(n4193), .CK(clk), .Q(\ram[225][11] ) );
  DFFHQX1 \ram_reg[225][10]  ( .D(n4192), .CK(clk), .Q(\ram[225][10] ) );
  DFFHQX1 \ram_reg[225][9]  ( .D(n4191), .CK(clk), .Q(\ram[225][9] ) );
  DFFHQX1 \ram_reg[225][8]  ( .D(n4190), .CK(clk), .Q(\ram[225][8] ) );
  DFFHQX1 \ram_reg[225][7]  ( .D(n4189), .CK(clk), .Q(\ram[225][7] ) );
  DFFHQX1 \ram_reg[225][6]  ( .D(n4188), .CK(clk), .Q(\ram[225][6] ) );
  DFFHQX1 \ram_reg[225][5]  ( .D(n4187), .CK(clk), .Q(\ram[225][5] ) );
  DFFHQX1 \ram_reg[225][4]  ( .D(n4186), .CK(clk), .Q(\ram[225][4] ) );
  DFFHQX1 \ram_reg[225][3]  ( .D(n4185), .CK(clk), .Q(\ram[225][3] ) );
  DFFHQX1 \ram_reg[225][2]  ( .D(n4184), .CK(clk), .Q(\ram[225][2] ) );
  DFFHQX1 \ram_reg[225][1]  ( .D(n4183), .CK(clk), .Q(\ram[225][1] ) );
  DFFHQX1 \ram_reg[225][0]  ( .D(n4182), .CK(clk), .Q(\ram[225][0] ) );
  DFFHQX1 \ram_reg[221][15]  ( .D(n4133), .CK(clk), .Q(\ram[221][15] ) );
  DFFHQX1 \ram_reg[221][14]  ( .D(n4132), .CK(clk), .Q(\ram[221][14] ) );
  DFFHQX1 \ram_reg[221][13]  ( .D(n4131), .CK(clk), .Q(\ram[221][13] ) );
  DFFHQX1 \ram_reg[221][12]  ( .D(n4130), .CK(clk), .Q(\ram[221][12] ) );
  DFFHQX1 \ram_reg[221][11]  ( .D(n4129), .CK(clk), .Q(\ram[221][11] ) );
  DFFHQX1 \ram_reg[221][10]  ( .D(n4128), .CK(clk), .Q(\ram[221][10] ) );
  DFFHQX1 \ram_reg[221][9]  ( .D(n4127), .CK(clk), .Q(\ram[221][9] ) );
  DFFHQX1 \ram_reg[221][8]  ( .D(n4126), .CK(clk), .Q(\ram[221][8] ) );
  DFFHQX1 \ram_reg[221][7]  ( .D(n4125), .CK(clk), .Q(\ram[221][7] ) );
  DFFHQX1 \ram_reg[221][6]  ( .D(n4124), .CK(clk), .Q(\ram[221][6] ) );
  DFFHQX1 \ram_reg[221][5]  ( .D(n4123), .CK(clk), .Q(\ram[221][5] ) );
  DFFHQX1 \ram_reg[221][4]  ( .D(n4122), .CK(clk), .Q(\ram[221][4] ) );
  DFFHQX1 \ram_reg[221][3]  ( .D(n4121), .CK(clk), .Q(\ram[221][3] ) );
  DFFHQX1 \ram_reg[221][2]  ( .D(n4120), .CK(clk), .Q(\ram[221][2] ) );
  DFFHQX1 \ram_reg[221][1]  ( .D(n4119), .CK(clk), .Q(\ram[221][1] ) );
  DFFHQX1 \ram_reg[221][0]  ( .D(n4118), .CK(clk), .Q(\ram[221][0] ) );
  DFFHQX1 \ram_reg[217][15]  ( .D(n4069), .CK(clk), .Q(\ram[217][15] ) );
  DFFHQX1 \ram_reg[217][14]  ( .D(n4068), .CK(clk), .Q(\ram[217][14] ) );
  DFFHQX1 \ram_reg[217][13]  ( .D(n4067), .CK(clk), .Q(\ram[217][13] ) );
  DFFHQX1 \ram_reg[217][12]  ( .D(n4066), .CK(clk), .Q(\ram[217][12] ) );
  DFFHQX1 \ram_reg[217][11]  ( .D(n4065), .CK(clk), .Q(\ram[217][11] ) );
  DFFHQX1 \ram_reg[217][10]  ( .D(n4064), .CK(clk), .Q(\ram[217][10] ) );
  DFFHQX1 \ram_reg[217][9]  ( .D(n4063), .CK(clk), .Q(\ram[217][9] ) );
  DFFHQX1 \ram_reg[217][8]  ( .D(n4062), .CK(clk), .Q(\ram[217][8] ) );
  DFFHQX1 \ram_reg[217][7]  ( .D(n4061), .CK(clk), .Q(\ram[217][7] ) );
  DFFHQX1 \ram_reg[217][6]  ( .D(n4060), .CK(clk), .Q(\ram[217][6] ) );
  DFFHQX1 \ram_reg[217][5]  ( .D(n4059), .CK(clk), .Q(\ram[217][5] ) );
  DFFHQX1 \ram_reg[217][4]  ( .D(n4058), .CK(clk), .Q(\ram[217][4] ) );
  DFFHQX1 \ram_reg[217][3]  ( .D(n4057), .CK(clk), .Q(\ram[217][3] ) );
  DFFHQX1 \ram_reg[217][2]  ( .D(n4056), .CK(clk), .Q(\ram[217][2] ) );
  DFFHQX1 \ram_reg[217][1]  ( .D(n4055), .CK(clk), .Q(\ram[217][1] ) );
  DFFHQX1 \ram_reg[217][0]  ( .D(n4054), .CK(clk), .Q(\ram[217][0] ) );
  DFFHQX1 \ram_reg[213][15]  ( .D(n4005), .CK(clk), .Q(\ram[213][15] ) );
  DFFHQX1 \ram_reg[213][14]  ( .D(n4004), .CK(clk), .Q(\ram[213][14] ) );
  DFFHQX1 \ram_reg[213][13]  ( .D(n4003), .CK(clk), .Q(\ram[213][13] ) );
  DFFHQX1 \ram_reg[213][12]  ( .D(n4002), .CK(clk), .Q(\ram[213][12] ) );
  DFFHQX1 \ram_reg[213][11]  ( .D(n4001), .CK(clk), .Q(\ram[213][11] ) );
  DFFHQX1 \ram_reg[213][10]  ( .D(n4000), .CK(clk), .Q(\ram[213][10] ) );
  DFFHQX1 \ram_reg[213][9]  ( .D(n3999), .CK(clk), .Q(\ram[213][9] ) );
  DFFHQX1 \ram_reg[213][8]  ( .D(n3998), .CK(clk), .Q(\ram[213][8] ) );
  DFFHQX1 \ram_reg[213][7]  ( .D(n3997), .CK(clk), .Q(\ram[213][7] ) );
  DFFHQX1 \ram_reg[213][6]  ( .D(n3996), .CK(clk), .Q(\ram[213][6] ) );
  DFFHQX1 \ram_reg[213][5]  ( .D(n3995), .CK(clk), .Q(\ram[213][5] ) );
  DFFHQX1 \ram_reg[213][4]  ( .D(n3994), .CK(clk), .Q(\ram[213][4] ) );
  DFFHQX1 \ram_reg[213][3]  ( .D(n3993), .CK(clk), .Q(\ram[213][3] ) );
  DFFHQX1 \ram_reg[213][2]  ( .D(n3992), .CK(clk), .Q(\ram[213][2] ) );
  DFFHQX1 \ram_reg[213][1]  ( .D(n3991), .CK(clk), .Q(\ram[213][1] ) );
  DFFHQX1 \ram_reg[213][0]  ( .D(n3990), .CK(clk), .Q(\ram[213][0] ) );
  DFFHQX1 \ram_reg[209][15]  ( .D(n3941), .CK(clk), .Q(\ram[209][15] ) );
  DFFHQX1 \ram_reg[209][14]  ( .D(n3940), .CK(clk), .Q(\ram[209][14] ) );
  DFFHQX1 \ram_reg[209][13]  ( .D(n3939), .CK(clk), .Q(\ram[209][13] ) );
  DFFHQX1 \ram_reg[209][12]  ( .D(n3938), .CK(clk), .Q(\ram[209][12] ) );
  DFFHQX1 \ram_reg[209][11]  ( .D(n3937), .CK(clk), .Q(\ram[209][11] ) );
  DFFHQX1 \ram_reg[209][10]  ( .D(n3936), .CK(clk), .Q(\ram[209][10] ) );
  DFFHQX1 \ram_reg[209][9]  ( .D(n3935), .CK(clk), .Q(\ram[209][9] ) );
  DFFHQX1 \ram_reg[209][8]  ( .D(n3934), .CK(clk), .Q(\ram[209][8] ) );
  DFFHQX1 \ram_reg[209][7]  ( .D(n3933), .CK(clk), .Q(\ram[209][7] ) );
  DFFHQX1 \ram_reg[209][6]  ( .D(n3932), .CK(clk), .Q(\ram[209][6] ) );
  DFFHQX1 \ram_reg[209][5]  ( .D(n3931), .CK(clk), .Q(\ram[209][5] ) );
  DFFHQX1 \ram_reg[209][4]  ( .D(n3930), .CK(clk), .Q(\ram[209][4] ) );
  DFFHQX1 \ram_reg[209][3]  ( .D(n3929), .CK(clk), .Q(\ram[209][3] ) );
  DFFHQX1 \ram_reg[209][2]  ( .D(n3928), .CK(clk), .Q(\ram[209][2] ) );
  DFFHQX1 \ram_reg[209][1]  ( .D(n3927), .CK(clk), .Q(\ram[209][1] ) );
  DFFHQX1 \ram_reg[209][0]  ( .D(n3926), .CK(clk), .Q(\ram[209][0] ) );
  DFFHQX1 \ram_reg[205][15]  ( .D(n3877), .CK(clk), .Q(\ram[205][15] ) );
  DFFHQX1 \ram_reg[205][14]  ( .D(n3876), .CK(clk), .Q(\ram[205][14] ) );
  DFFHQX1 \ram_reg[205][13]  ( .D(n3875), .CK(clk), .Q(\ram[205][13] ) );
  DFFHQX1 \ram_reg[205][12]  ( .D(n3874), .CK(clk), .Q(\ram[205][12] ) );
  DFFHQX1 \ram_reg[205][11]  ( .D(n3873), .CK(clk), .Q(\ram[205][11] ) );
  DFFHQX1 \ram_reg[205][10]  ( .D(n3872), .CK(clk), .Q(\ram[205][10] ) );
  DFFHQX1 \ram_reg[205][9]  ( .D(n3871), .CK(clk), .Q(\ram[205][9] ) );
  DFFHQX1 \ram_reg[205][8]  ( .D(n3870), .CK(clk), .Q(\ram[205][8] ) );
  DFFHQX1 \ram_reg[205][7]  ( .D(n3869), .CK(clk), .Q(\ram[205][7] ) );
  DFFHQX1 \ram_reg[205][6]  ( .D(n3868), .CK(clk), .Q(\ram[205][6] ) );
  DFFHQX1 \ram_reg[205][5]  ( .D(n3867), .CK(clk), .Q(\ram[205][5] ) );
  DFFHQX1 \ram_reg[205][4]  ( .D(n3866), .CK(clk), .Q(\ram[205][4] ) );
  DFFHQX1 \ram_reg[205][3]  ( .D(n3865), .CK(clk), .Q(\ram[205][3] ) );
  DFFHQX1 \ram_reg[205][2]  ( .D(n3864), .CK(clk), .Q(\ram[205][2] ) );
  DFFHQX1 \ram_reg[205][1]  ( .D(n3863), .CK(clk), .Q(\ram[205][1] ) );
  DFFHQX1 \ram_reg[205][0]  ( .D(n3862), .CK(clk), .Q(\ram[205][0] ) );
  DFFHQX1 \ram_reg[201][15]  ( .D(n3813), .CK(clk), .Q(\ram[201][15] ) );
  DFFHQX1 \ram_reg[201][14]  ( .D(n3812), .CK(clk), .Q(\ram[201][14] ) );
  DFFHQX1 \ram_reg[201][13]  ( .D(n3811), .CK(clk), .Q(\ram[201][13] ) );
  DFFHQX1 \ram_reg[201][12]  ( .D(n3810), .CK(clk), .Q(\ram[201][12] ) );
  DFFHQX1 \ram_reg[201][11]  ( .D(n3809), .CK(clk), .Q(\ram[201][11] ) );
  DFFHQX1 \ram_reg[201][10]  ( .D(n3808), .CK(clk), .Q(\ram[201][10] ) );
  DFFHQX1 \ram_reg[201][9]  ( .D(n3807), .CK(clk), .Q(\ram[201][9] ) );
  DFFHQX1 \ram_reg[201][8]  ( .D(n3806), .CK(clk), .Q(\ram[201][8] ) );
  DFFHQX1 \ram_reg[201][7]  ( .D(n3805), .CK(clk), .Q(\ram[201][7] ) );
  DFFHQX1 \ram_reg[201][6]  ( .D(n3804), .CK(clk), .Q(\ram[201][6] ) );
  DFFHQX1 \ram_reg[201][5]  ( .D(n3803), .CK(clk), .Q(\ram[201][5] ) );
  DFFHQX1 \ram_reg[201][4]  ( .D(n3802), .CK(clk), .Q(\ram[201][4] ) );
  DFFHQX1 \ram_reg[201][3]  ( .D(n3801), .CK(clk), .Q(\ram[201][3] ) );
  DFFHQX1 \ram_reg[201][2]  ( .D(n3800), .CK(clk), .Q(\ram[201][2] ) );
  DFFHQX1 \ram_reg[201][1]  ( .D(n3799), .CK(clk), .Q(\ram[201][1] ) );
  DFFHQX1 \ram_reg[201][0]  ( .D(n3798), .CK(clk), .Q(\ram[201][0] ) );
  DFFHQX1 \ram_reg[197][15]  ( .D(n3749), .CK(clk), .Q(\ram[197][15] ) );
  DFFHQX1 \ram_reg[197][14]  ( .D(n3748), .CK(clk), .Q(\ram[197][14] ) );
  DFFHQX1 \ram_reg[197][13]  ( .D(n3747), .CK(clk), .Q(\ram[197][13] ) );
  DFFHQX1 \ram_reg[197][12]  ( .D(n3746), .CK(clk), .Q(\ram[197][12] ) );
  DFFHQX1 \ram_reg[197][11]  ( .D(n3745), .CK(clk), .Q(\ram[197][11] ) );
  DFFHQX1 \ram_reg[197][10]  ( .D(n3744), .CK(clk), .Q(\ram[197][10] ) );
  DFFHQX1 \ram_reg[197][9]  ( .D(n3743), .CK(clk), .Q(\ram[197][9] ) );
  DFFHQX1 \ram_reg[197][8]  ( .D(n3742), .CK(clk), .Q(\ram[197][8] ) );
  DFFHQX1 \ram_reg[197][7]  ( .D(n3741), .CK(clk), .Q(\ram[197][7] ) );
  DFFHQX1 \ram_reg[197][6]  ( .D(n3740), .CK(clk), .Q(\ram[197][6] ) );
  DFFHQX1 \ram_reg[197][5]  ( .D(n3739), .CK(clk), .Q(\ram[197][5] ) );
  DFFHQX1 \ram_reg[197][4]  ( .D(n3738), .CK(clk), .Q(\ram[197][4] ) );
  DFFHQX1 \ram_reg[197][3]  ( .D(n3737), .CK(clk), .Q(\ram[197][3] ) );
  DFFHQX1 \ram_reg[197][2]  ( .D(n3736), .CK(clk), .Q(\ram[197][2] ) );
  DFFHQX1 \ram_reg[197][1]  ( .D(n3735), .CK(clk), .Q(\ram[197][1] ) );
  DFFHQX1 \ram_reg[197][0]  ( .D(n3734), .CK(clk), .Q(\ram[197][0] ) );
  DFFHQX1 \ram_reg[193][15]  ( .D(n3685), .CK(clk), .Q(\ram[193][15] ) );
  DFFHQX1 \ram_reg[193][14]  ( .D(n3684), .CK(clk), .Q(\ram[193][14] ) );
  DFFHQX1 \ram_reg[193][13]  ( .D(n3683), .CK(clk), .Q(\ram[193][13] ) );
  DFFHQX1 \ram_reg[193][12]  ( .D(n3682), .CK(clk), .Q(\ram[193][12] ) );
  DFFHQX1 \ram_reg[193][11]  ( .D(n3681), .CK(clk), .Q(\ram[193][11] ) );
  DFFHQX1 \ram_reg[193][10]  ( .D(n3680), .CK(clk), .Q(\ram[193][10] ) );
  DFFHQX1 \ram_reg[193][9]  ( .D(n3679), .CK(clk), .Q(\ram[193][9] ) );
  DFFHQX1 \ram_reg[193][8]  ( .D(n3678), .CK(clk), .Q(\ram[193][8] ) );
  DFFHQX1 \ram_reg[193][7]  ( .D(n3677), .CK(clk), .Q(\ram[193][7] ) );
  DFFHQX1 \ram_reg[193][6]  ( .D(n3676), .CK(clk), .Q(\ram[193][6] ) );
  DFFHQX1 \ram_reg[193][5]  ( .D(n3675), .CK(clk), .Q(\ram[193][5] ) );
  DFFHQX1 \ram_reg[193][4]  ( .D(n3674), .CK(clk), .Q(\ram[193][4] ) );
  DFFHQX1 \ram_reg[193][3]  ( .D(n3673), .CK(clk), .Q(\ram[193][3] ) );
  DFFHQX1 \ram_reg[193][2]  ( .D(n3672), .CK(clk), .Q(\ram[193][2] ) );
  DFFHQX1 \ram_reg[193][1]  ( .D(n3671), .CK(clk), .Q(\ram[193][1] ) );
  DFFHQX1 \ram_reg[193][0]  ( .D(n3670), .CK(clk), .Q(\ram[193][0] ) );
  DFFHQX1 \ram_reg[189][15]  ( .D(n3621), .CK(clk), .Q(\ram[189][15] ) );
  DFFHQX1 \ram_reg[189][14]  ( .D(n3620), .CK(clk), .Q(\ram[189][14] ) );
  DFFHQX1 \ram_reg[189][13]  ( .D(n3619), .CK(clk), .Q(\ram[189][13] ) );
  DFFHQX1 \ram_reg[189][12]  ( .D(n3618), .CK(clk), .Q(\ram[189][12] ) );
  DFFHQX1 \ram_reg[189][11]  ( .D(n3617), .CK(clk), .Q(\ram[189][11] ) );
  DFFHQX1 \ram_reg[189][10]  ( .D(n3616), .CK(clk), .Q(\ram[189][10] ) );
  DFFHQX1 \ram_reg[189][9]  ( .D(n3615), .CK(clk), .Q(\ram[189][9] ) );
  DFFHQX1 \ram_reg[189][8]  ( .D(n3614), .CK(clk), .Q(\ram[189][8] ) );
  DFFHQX1 \ram_reg[189][7]  ( .D(n3613), .CK(clk), .Q(\ram[189][7] ) );
  DFFHQX1 \ram_reg[189][6]  ( .D(n3612), .CK(clk), .Q(\ram[189][6] ) );
  DFFHQX1 \ram_reg[189][5]  ( .D(n3611), .CK(clk), .Q(\ram[189][5] ) );
  DFFHQX1 \ram_reg[189][4]  ( .D(n3610), .CK(clk), .Q(\ram[189][4] ) );
  DFFHQX1 \ram_reg[189][3]  ( .D(n3609), .CK(clk), .Q(\ram[189][3] ) );
  DFFHQX1 \ram_reg[189][2]  ( .D(n3608), .CK(clk), .Q(\ram[189][2] ) );
  DFFHQX1 \ram_reg[189][1]  ( .D(n3607), .CK(clk), .Q(\ram[189][1] ) );
  DFFHQX1 \ram_reg[189][0]  ( .D(n3606), .CK(clk), .Q(\ram[189][0] ) );
  DFFHQX1 \ram_reg[185][15]  ( .D(n3557), .CK(clk), .Q(\ram[185][15] ) );
  DFFHQX1 \ram_reg[185][14]  ( .D(n3556), .CK(clk), .Q(\ram[185][14] ) );
  DFFHQX1 \ram_reg[185][13]  ( .D(n3555), .CK(clk), .Q(\ram[185][13] ) );
  DFFHQX1 \ram_reg[185][12]  ( .D(n3554), .CK(clk), .Q(\ram[185][12] ) );
  DFFHQX1 \ram_reg[185][11]  ( .D(n3553), .CK(clk), .Q(\ram[185][11] ) );
  DFFHQX1 \ram_reg[185][10]  ( .D(n3552), .CK(clk), .Q(\ram[185][10] ) );
  DFFHQX1 \ram_reg[185][9]  ( .D(n3551), .CK(clk), .Q(\ram[185][9] ) );
  DFFHQX1 \ram_reg[185][8]  ( .D(n3550), .CK(clk), .Q(\ram[185][8] ) );
  DFFHQX1 \ram_reg[185][7]  ( .D(n3549), .CK(clk), .Q(\ram[185][7] ) );
  DFFHQX1 \ram_reg[185][6]  ( .D(n3548), .CK(clk), .Q(\ram[185][6] ) );
  DFFHQX1 \ram_reg[185][5]  ( .D(n3547), .CK(clk), .Q(\ram[185][5] ) );
  DFFHQX1 \ram_reg[185][4]  ( .D(n3546), .CK(clk), .Q(\ram[185][4] ) );
  DFFHQX1 \ram_reg[185][3]  ( .D(n3545), .CK(clk), .Q(\ram[185][3] ) );
  DFFHQX1 \ram_reg[185][2]  ( .D(n3544), .CK(clk), .Q(\ram[185][2] ) );
  DFFHQX1 \ram_reg[185][1]  ( .D(n3543), .CK(clk), .Q(\ram[185][1] ) );
  DFFHQX1 \ram_reg[185][0]  ( .D(n3542), .CK(clk), .Q(\ram[185][0] ) );
  DFFHQX1 \ram_reg[181][15]  ( .D(n3493), .CK(clk), .Q(\ram[181][15] ) );
  DFFHQX1 \ram_reg[181][14]  ( .D(n3492), .CK(clk), .Q(\ram[181][14] ) );
  DFFHQX1 \ram_reg[181][13]  ( .D(n3491), .CK(clk), .Q(\ram[181][13] ) );
  DFFHQX1 \ram_reg[181][12]  ( .D(n3490), .CK(clk), .Q(\ram[181][12] ) );
  DFFHQX1 \ram_reg[181][11]  ( .D(n3489), .CK(clk), .Q(\ram[181][11] ) );
  DFFHQX1 \ram_reg[181][10]  ( .D(n3488), .CK(clk), .Q(\ram[181][10] ) );
  DFFHQX1 \ram_reg[181][9]  ( .D(n3487), .CK(clk), .Q(\ram[181][9] ) );
  DFFHQX1 \ram_reg[181][8]  ( .D(n3486), .CK(clk), .Q(\ram[181][8] ) );
  DFFHQX1 \ram_reg[181][7]  ( .D(n3485), .CK(clk), .Q(\ram[181][7] ) );
  DFFHQX1 \ram_reg[181][6]  ( .D(n3484), .CK(clk), .Q(\ram[181][6] ) );
  DFFHQX1 \ram_reg[181][5]  ( .D(n3483), .CK(clk), .Q(\ram[181][5] ) );
  DFFHQX1 \ram_reg[181][4]  ( .D(n3482), .CK(clk), .Q(\ram[181][4] ) );
  DFFHQX1 \ram_reg[181][3]  ( .D(n3481), .CK(clk), .Q(\ram[181][3] ) );
  DFFHQX1 \ram_reg[181][2]  ( .D(n3480), .CK(clk), .Q(\ram[181][2] ) );
  DFFHQX1 \ram_reg[181][1]  ( .D(n3479), .CK(clk), .Q(\ram[181][1] ) );
  DFFHQX1 \ram_reg[181][0]  ( .D(n3478), .CK(clk), .Q(\ram[181][0] ) );
  DFFHQX1 \ram_reg[177][15]  ( .D(n3429), .CK(clk), .Q(\ram[177][15] ) );
  DFFHQX1 \ram_reg[177][14]  ( .D(n3428), .CK(clk), .Q(\ram[177][14] ) );
  DFFHQX1 \ram_reg[177][13]  ( .D(n3427), .CK(clk), .Q(\ram[177][13] ) );
  DFFHQX1 \ram_reg[177][12]  ( .D(n3426), .CK(clk), .Q(\ram[177][12] ) );
  DFFHQX1 \ram_reg[177][11]  ( .D(n3425), .CK(clk), .Q(\ram[177][11] ) );
  DFFHQX1 \ram_reg[177][10]  ( .D(n3424), .CK(clk), .Q(\ram[177][10] ) );
  DFFHQX1 \ram_reg[177][9]  ( .D(n3423), .CK(clk), .Q(\ram[177][9] ) );
  DFFHQX1 \ram_reg[177][8]  ( .D(n3422), .CK(clk), .Q(\ram[177][8] ) );
  DFFHQX1 \ram_reg[177][7]  ( .D(n3421), .CK(clk), .Q(\ram[177][7] ) );
  DFFHQX1 \ram_reg[177][6]  ( .D(n3420), .CK(clk), .Q(\ram[177][6] ) );
  DFFHQX1 \ram_reg[177][5]  ( .D(n3419), .CK(clk), .Q(\ram[177][5] ) );
  DFFHQX1 \ram_reg[177][4]  ( .D(n3418), .CK(clk), .Q(\ram[177][4] ) );
  DFFHQX1 \ram_reg[177][3]  ( .D(n3417), .CK(clk), .Q(\ram[177][3] ) );
  DFFHQX1 \ram_reg[177][2]  ( .D(n3416), .CK(clk), .Q(\ram[177][2] ) );
  DFFHQX1 \ram_reg[177][1]  ( .D(n3415), .CK(clk), .Q(\ram[177][1] ) );
  DFFHQX1 \ram_reg[177][0]  ( .D(n3414), .CK(clk), .Q(\ram[177][0] ) );
  DFFHQX1 \ram_reg[173][15]  ( .D(n3365), .CK(clk), .Q(\ram[173][15] ) );
  DFFHQX1 \ram_reg[173][14]  ( .D(n3364), .CK(clk), .Q(\ram[173][14] ) );
  DFFHQX1 \ram_reg[173][13]  ( .D(n3363), .CK(clk), .Q(\ram[173][13] ) );
  DFFHQX1 \ram_reg[173][12]  ( .D(n3362), .CK(clk), .Q(\ram[173][12] ) );
  DFFHQX1 \ram_reg[173][11]  ( .D(n3361), .CK(clk), .Q(\ram[173][11] ) );
  DFFHQX1 \ram_reg[173][10]  ( .D(n3360), .CK(clk), .Q(\ram[173][10] ) );
  DFFHQX1 \ram_reg[173][9]  ( .D(n3359), .CK(clk), .Q(\ram[173][9] ) );
  DFFHQX1 \ram_reg[173][8]  ( .D(n3358), .CK(clk), .Q(\ram[173][8] ) );
  DFFHQX1 \ram_reg[173][7]  ( .D(n3357), .CK(clk), .Q(\ram[173][7] ) );
  DFFHQX1 \ram_reg[173][6]  ( .D(n3356), .CK(clk), .Q(\ram[173][6] ) );
  DFFHQX1 \ram_reg[173][5]  ( .D(n3355), .CK(clk), .Q(\ram[173][5] ) );
  DFFHQX1 \ram_reg[173][4]  ( .D(n3354), .CK(clk), .Q(\ram[173][4] ) );
  DFFHQX1 \ram_reg[173][3]  ( .D(n3353), .CK(clk), .Q(\ram[173][3] ) );
  DFFHQX1 \ram_reg[173][2]  ( .D(n3352), .CK(clk), .Q(\ram[173][2] ) );
  DFFHQX1 \ram_reg[173][1]  ( .D(n3351), .CK(clk), .Q(\ram[173][1] ) );
  DFFHQX1 \ram_reg[173][0]  ( .D(n3350), .CK(clk), .Q(\ram[173][0] ) );
  DFFHQX1 \ram_reg[169][15]  ( .D(n3301), .CK(clk), .Q(\ram[169][15] ) );
  DFFHQX1 \ram_reg[169][14]  ( .D(n3300), .CK(clk), .Q(\ram[169][14] ) );
  DFFHQX1 \ram_reg[169][13]  ( .D(n3299), .CK(clk), .Q(\ram[169][13] ) );
  DFFHQX1 \ram_reg[169][12]  ( .D(n3298), .CK(clk), .Q(\ram[169][12] ) );
  DFFHQX1 \ram_reg[169][11]  ( .D(n3297), .CK(clk), .Q(\ram[169][11] ) );
  DFFHQX1 \ram_reg[169][10]  ( .D(n3296), .CK(clk), .Q(\ram[169][10] ) );
  DFFHQX1 \ram_reg[169][9]  ( .D(n3295), .CK(clk), .Q(\ram[169][9] ) );
  DFFHQX1 \ram_reg[169][8]  ( .D(n3294), .CK(clk), .Q(\ram[169][8] ) );
  DFFHQX1 \ram_reg[169][7]  ( .D(n3293), .CK(clk), .Q(\ram[169][7] ) );
  DFFHQX1 \ram_reg[169][6]  ( .D(n3292), .CK(clk), .Q(\ram[169][6] ) );
  DFFHQX1 \ram_reg[169][5]  ( .D(n3291), .CK(clk), .Q(\ram[169][5] ) );
  DFFHQX1 \ram_reg[169][4]  ( .D(n3290), .CK(clk), .Q(\ram[169][4] ) );
  DFFHQX1 \ram_reg[169][3]  ( .D(n3289), .CK(clk), .Q(\ram[169][3] ) );
  DFFHQX1 \ram_reg[169][2]  ( .D(n3288), .CK(clk), .Q(\ram[169][2] ) );
  DFFHQX1 \ram_reg[169][1]  ( .D(n3287), .CK(clk), .Q(\ram[169][1] ) );
  DFFHQX1 \ram_reg[169][0]  ( .D(n3286), .CK(clk), .Q(\ram[169][0] ) );
  DFFHQX1 \ram_reg[165][15]  ( .D(n3237), .CK(clk), .Q(\ram[165][15] ) );
  DFFHQX1 \ram_reg[165][14]  ( .D(n3236), .CK(clk), .Q(\ram[165][14] ) );
  DFFHQX1 \ram_reg[165][13]  ( .D(n3235), .CK(clk), .Q(\ram[165][13] ) );
  DFFHQX1 \ram_reg[165][12]  ( .D(n3234), .CK(clk), .Q(\ram[165][12] ) );
  DFFHQX1 \ram_reg[165][11]  ( .D(n3233), .CK(clk), .Q(\ram[165][11] ) );
  DFFHQX1 \ram_reg[165][10]  ( .D(n3232), .CK(clk), .Q(\ram[165][10] ) );
  DFFHQX1 \ram_reg[165][9]  ( .D(n3231), .CK(clk), .Q(\ram[165][9] ) );
  DFFHQX1 \ram_reg[165][8]  ( .D(n3230), .CK(clk), .Q(\ram[165][8] ) );
  DFFHQX1 \ram_reg[165][7]  ( .D(n3229), .CK(clk), .Q(\ram[165][7] ) );
  DFFHQX1 \ram_reg[165][6]  ( .D(n3228), .CK(clk), .Q(\ram[165][6] ) );
  DFFHQX1 \ram_reg[165][5]  ( .D(n3227), .CK(clk), .Q(\ram[165][5] ) );
  DFFHQX1 \ram_reg[165][4]  ( .D(n3226), .CK(clk), .Q(\ram[165][4] ) );
  DFFHQX1 \ram_reg[165][3]  ( .D(n3225), .CK(clk), .Q(\ram[165][3] ) );
  DFFHQX1 \ram_reg[165][2]  ( .D(n3224), .CK(clk), .Q(\ram[165][2] ) );
  DFFHQX1 \ram_reg[165][1]  ( .D(n3223), .CK(clk), .Q(\ram[165][1] ) );
  DFFHQX1 \ram_reg[165][0]  ( .D(n3222), .CK(clk), .Q(\ram[165][0] ) );
  DFFHQX1 \ram_reg[161][15]  ( .D(n3173), .CK(clk), .Q(\ram[161][15] ) );
  DFFHQX1 \ram_reg[161][14]  ( .D(n3172), .CK(clk), .Q(\ram[161][14] ) );
  DFFHQX1 \ram_reg[161][13]  ( .D(n3171), .CK(clk), .Q(\ram[161][13] ) );
  DFFHQX1 \ram_reg[161][12]  ( .D(n3170), .CK(clk), .Q(\ram[161][12] ) );
  DFFHQX1 \ram_reg[161][11]  ( .D(n3169), .CK(clk), .Q(\ram[161][11] ) );
  DFFHQX1 \ram_reg[161][10]  ( .D(n3168), .CK(clk), .Q(\ram[161][10] ) );
  DFFHQX1 \ram_reg[161][9]  ( .D(n3167), .CK(clk), .Q(\ram[161][9] ) );
  DFFHQX1 \ram_reg[161][8]  ( .D(n3166), .CK(clk), .Q(\ram[161][8] ) );
  DFFHQX1 \ram_reg[161][7]  ( .D(n3165), .CK(clk), .Q(\ram[161][7] ) );
  DFFHQX1 \ram_reg[161][6]  ( .D(n3164), .CK(clk), .Q(\ram[161][6] ) );
  DFFHQX1 \ram_reg[161][5]  ( .D(n3163), .CK(clk), .Q(\ram[161][5] ) );
  DFFHQX1 \ram_reg[161][4]  ( .D(n3162), .CK(clk), .Q(\ram[161][4] ) );
  DFFHQX1 \ram_reg[161][3]  ( .D(n3161), .CK(clk), .Q(\ram[161][3] ) );
  DFFHQX1 \ram_reg[161][2]  ( .D(n3160), .CK(clk), .Q(\ram[161][2] ) );
  DFFHQX1 \ram_reg[161][1]  ( .D(n3159), .CK(clk), .Q(\ram[161][1] ) );
  DFFHQX1 \ram_reg[161][0]  ( .D(n3158), .CK(clk), .Q(\ram[161][0] ) );
  DFFHQX1 \ram_reg[157][15]  ( .D(n3109), .CK(clk), .Q(\ram[157][15] ) );
  DFFHQX1 \ram_reg[157][14]  ( .D(n3108), .CK(clk), .Q(\ram[157][14] ) );
  DFFHQX1 \ram_reg[157][13]  ( .D(n3107), .CK(clk), .Q(\ram[157][13] ) );
  DFFHQX1 \ram_reg[157][12]  ( .D(n3106), .CK(clk), .Q(\ram[157][12] ) );
  DFFHQX1 \ram_reg[157][11]  ( .D(n3105), .CK(clk), .Q(\ram[157][11] ) );
  DFFHQX1 \ram_reg[157][10]  ( .D(n3104), .CK(clk), .Q(\ram[157][10] ) );
  DFFHQX1 \ram_reg[157][9]  ( .D(n3103), .CK(clk), .Q(\ram[157][9] ) );
  DFFHQX1 \ram_reg[157][8]  ( .D(n3102), .CK(clk), .Q(\ram[157][8] ) );
  DFFHQX1 \ram_reg[157][7]  ( .D(n3101), .CK(clk), .Q(\ram[157][7] ) );
  DFFHQX1 \ram_reg[157][6]  ( .D(n3100), .CK(clk), .Q(\ram[157][6] ) );
  DFFHQX1 \ram_reg[157][5]  ( .D(n3099), .CK(clk), .Q(\ram[157][5] ) );
  DFFHQX1 \ram_reg[157][4]  ( .D(n3098), .CK(clk), .Q(\ram[157][4] ) );
  DFFHQX1 \ram_reg[157][3]  ( .D(n3097), .CK(clk), .Q(\ram[157][3] ) );
  DFFHQX1 \ram_reg[157][2]  ( .D(n3096), .CK(clk), .Q(\ram[157][2] ) );
  DFFHQX1 \ram_reg[157][1]  ( .D(n3095), .CK(clk), .Q(\ram[157][1] ) );
  DFFHQX1 \ram_reg[157][0]  ( .D(n3094), .CK(clk), .Q(\ram[157][0] ) );
  DFFHQX1 \ram_reg[153][15]  ( .D(n3045), .CK(clk), .Q(\ram[153][15] ) );
  DFFHQX1 \ram_reg[153][14]  ( .D(n3044), .CK(clk), .Q(\ram[153][14] ) );
  DFFHQX1 \ram_reg[153][13]  ( .D(n3043), .CK(clk), .Q(\ram[153][13] ) );
  DFFHQX1 \ram_reg[153][12]  ( .D(n3042), .CK(clk), .Q(\ram[153][12] ) );
  DFFHQX1 \ram_reg[153][11]  ( .D(n3041), .CK(clk), .Q(\ram[153][11] ) );
  DFFHQX1 \ram_reg[153][10]  ( .D(n3040), .CK(clk), .Q(\ram[153][10] ) );
  DFFHQX1 \ram_reg[153][9]  ( .D(n3039), .CK(clk), .Q(\ram[153][9] ) );
  DFFHQX1 \ram_reg[153][8]  ( .D(n3038), .CK(clk), .Q(\ram[153][8] ) );
  DFFHQX1 \ram_reg[153][7]  ( .D(n3037), .CK(clk), .Q(\ram[153][7] ) );
  DFFHQX1 \ram_reg[153][6]  ( .D(n3036), .CK(clk), .Q(\ram[153][6] ) );
  DFFHQX1 \ram_reg[153][5]  ( .D(n3035), .CK(clk), .Q(\ram[153][5] ) );
  DFFHQX1 \ram_reg[153][4]  ( .D(n3034), .CK(clk), .Q(\ram[153][4] ) );
  DFFHQX1 \ram_reg[153][3]  ( .D(n3033), .CK(clk), .Q(\ram[153][3] ) );
  DFFHQX1 \ram_reg[153][2]  ( .D(n3032), .CK(clk), .Q(\ram[153][2] ) );
  DFFHQX1 \ram_reg[153][1]  ( .D(n3031), .CK(clk), .Q(\ram[153][1] ) );
  DFFHQX1 \ram_reg[153][0]  ( .D(n3030), .CK(clk), .Q(\ram[153][0] ) );
  DFFHQX1 \ram_reg[149][15]  ( .D(n2981), .CK(clk), .Q(\ram[149][15] ) );
  DFFHQX1 \ram_reg[149][14]  ( .D(n2980), .CK(clk), .Q(\ram[149][14] ) );
  DFFHQX1 \ram_reg[149][13]  ( .D(n2979), .CK(clk), .Q(\ram[149][13] ) );
  DFFHQX1 \ram_reg[149][12]  ( .D(n2978), .CK(clk), .Q(\ram[149][12] ) );
  DFFHQX1 \ram_reg[149][11]  ( .D(n2977), .CK(clk), .Q(\ram[149][11] ) );
  DFFHQX1 \ram_reg[149][10]  ( .D(n2976), .CK(clk), .Q(\ram[149][10] ) );
  DFFHQX1 \ram_reg[149][9]  ( .D(n2975), .CK(clk), .Q(\ram[149][9] ) );
  DFFHQX1 \ram_reg[149][8]  ( .D(n2974), .CK(clk), .Q(\ram[149][8] ) );
  DFFHQX1 \ram_reg[149][7]  ( .D(n2973), .CK(clk), .Q(\ram[149][7] ) );
  DFFHQX1 \ram_reg[149][6]  ( .D(n2972), .CK(clk), .Q(\ram[149][6] ) );
  DFFHQX1 \ram_reg[149][5]  ( .D(n2971), .CK(clk), .Q(\ram[149][5] ) );
  DFFHQX1 \ram_reg[149][4]  ( .D(n2970), .CK(clk), .Q(\ram[149][4] ) );
  DFFHQX1 \ram_reg[149][3]  ( .D(n2969), .CK(clk), .Q(\ram[149][3] ) );
  DFFHQX1 \ram_reg[149][2]  ( .D(n2968), .CK(clk), .Q(\ram[149][2] ) );
  DFFHQX1 \ram_reg[149][1]  ( .D(n2967), .CK(clk), .Q(\ram[149][1] ) );
  DFFHQX1 \ram_reg[149][0]  ( .D(n2966), .CK(clk), .Q(\ram[149][0] ) );
  DFFHQX1 \ram_reg[145][15]  ( .D(n2917), .CK(clk), .Q(\ram[145][15] ) );
  DFFHQX1 \ram_reg[145][14]  ( .D(n2916), .CK(clk), .Q(\ram[145][14] ) );
  DFFHQX1 \ram_reg[145][13]  ( .D(n2915), .CK(clk), .Q(\ram[145][13] ) );
  DFFHQX1 \ram_reg[145][12]  ( .D(n2914), .CK(clk), .Q(\ram[145][12] ) );
  DFFHQX1 \ram_reg[145][11]  ( .D(n2913), .CK(clk), .Q(\ram[145][11] ) );
  DFFHQX1 \ram_reg[145][10]  ( .D(n2912), .CK(clk), .Q(\ram[145][10] ) );
  DFFHQX1 \ram_reg[145][9]  ( .D(n2911), .CK(clk), .Q(\ram[145][9] ) );
  DFFHQX1 \ram_reg[145][8]  ( .D(n2910), .CK(clk), .Q(\ram[145][8] ) );
  DFFHQX1 \ram_reg[145][7]  ( .D(n2909), .CK(clk), .Q(\ram[145][7] ) );
  DFFHQX1 \ram_reg[145][6]  ( .D(n2908), .CK(clk), .Q(\ram[145][6] ) );
  DFFHQX1 \ram_reg[145][5]  ( .D(n2907), .CK(clk), .Q(\ram[145][5] ) );
  DFFHQX1 \ram_reg[145][4]  ( .D(n2906), .CK(clk), .Q(\ram[145][4] ) );
  DFFHQX1 \ram_reg[145][3]  ( .D(n2905), .CK(clk), .Q(\ram[145][3] ) );
  DFFHQX1 \ram_reg[145][2]  ( .D(n2904), .CK(clk), .Q(\ram[145][2] ) );
  DFFHQX1 \ram_reg[145][1]  ( .D(n2903), .CK(clk), .Q(\ram[145][1] ) );
  DFFHQX1 \ram_reg[145][0]  ( .D(n2902), .CK(clk), .Q(\ram[145][0] ) );
  DFFHQX1 \ram_reg[141][15]  ( .D(n2853), .CK(clk), .Q(\ram[141][15] ) );
  DFFHQX1 \ram_reg[141][14]  ( .D(n2852), .CK(clk), .Q(\ram[141][14] ) );
  DFFHQX1 \ram_reg[141][13]  ( .D(n2851), .CK(clk), .Q(\ram[141][13] ) );
  DFFHQX1 \ram_reg[141][12]  ( .D(n2850), .CK(clk), .Q(\ram[141][12] ) );
  DFFHQX1 \ram_reg[141][11]  ( .D(n2849), .CK(clk), .Q(\ram[141][11] ) );
  DFFHQX1 \ram_reg[141][10]  ( .D(n2848), .CK(clk), .Q(\ram[141][10] ) );
  DFFHQX1 \ram_reg[141][9]  ( .D(n2847), .CK(clk), .Q(\ram[141][9] ) );
  DFFHQX1 \ram_reg[141][8]  ( .D(n2846), .CK(clk), .Q(\ram[141][8] ) );
  DFFHQX1 \ram_reg[141][7]  ( .D(n2845), .CK(clk), .Q(\ram[141][7] ) );
  DFFHQX1 \ram_reg[141][6]  ( .D(n2844), .CK(clk), .Q(\ram[141][6] ) );
  DFFHQX1 \ram_reg[141][5]  ( .D(n2843), .CK(clk), .Q(\ram[141][5] ) );
  DFFHQX1 \ram_reg[141][4]  ( .D(n2842), .CK(clk), .Q(\ram[141][4] ) );
  DFFHQX1 \ram_reg[141][3]  ( .D(n2841), .CK(clk), .Q(\ram[141][3] ) );
  DFFHQX1 \ram_reg[141][2]  ( .D(n2840), .CK(clk), .Q(\ram[141][2] ) );
  DFFHQX1 \ram_reg[141][1]  ( .D(n2839), .CK(clk), .Q(\ram[141][1] ) );
  DFFHQX1 \ram_reg[141][0]  ( .D(n2838), .CK(clk), .Q(\ram[141][0] ) );
  DFFHQX1 \ram_reg[137][15]  ( .D(n2789), .CK(clk), .Q(\ram[137][15] ) );
  DFFHQX1 \ram_reg[137][14]  ( .D(n2788), .CK(clk), .Q(\ram[137][14] ) );
  DFFHQX1 \ram_reg[137][13]  ( .D(n2787), .CK(clk), .Q(\ram[137][13] ) );
  DFFHQX1 \ram_reg[137][12]  ( .D(n2786), .CK(clk), .Q(\ram[137][12] ) );
  DFFHQX1 \ram_reg[137][11]  ( .D(n2785), .CK(clk), .Q(\ram[137][11] ) );
  DFFHQX1 \ram_reg[137][10]  ( .D(n2784), .CK(clk), .Q(\ram[137][10] ) );
  DFFHQX1 \ram_reg[137][9]  ( .D(n2783), .CK(clk), .Q(\ram[137][9] ) );
  DFFHQX1 \ram_reg[137][8]  ( .D(n2782), .CK(clk), .Q(\ram[137][8] ) );
  DFFHQX1 \ram_reg[137][7]  ( .D(n2781), .CK(clk), .Q(\ram[137][7] ) );
  DFFHQX1 \ram_reg[137][6]  ( .D(n2780), .CK(clk), .Q(\ram[137][6] ) );
  DFFHQX1 \ram_reg[137][5]  ( .D(n2779), .CK(clk), .Q(\ram[137][5] ) );
  DFFHQX1 \ram_reg[137][4]  ( .D(n2778), .CK(clk), .Q(\ram[137][4] ) );
  DFFHQX1 \ram_reg[137][3]  ( .D(n2777), .CK(clk), .Q(\ram[137][3] ) );
  DFFHQX1 \ram_reg[137][2]  ( .D(n2776), .CK(clk), .Q(\ram[137][2] ) );
  DFFHQX1 \ram_reg[137][1]  ( .D(n2775), .CK(clk), .Q(\ram[137][1] ) );
  DFFHQX1 \ram_reg[137][0]  ( .D(n2774), .CK(clk), .Q(\ram[137][0] ) );
  DFFHQX1 \ram_reg[133][15]  ( .D(n2725), .CK(clk), .Q(\ram[133][15] ) );
  DFFHQX1 \ram_reg[133][14]  ( .D(n2724), .CK(clk), .Q(\ram[133][14] ) );
  DFFHQX1 \ram_reg[133][13]  ( .D(n2723), .CK(clk), .Q(\ram[133][13] ) );
  DFFHQX1 \ram_reg[133][12]  ( .D(n2722), .CK(clk), .Q(\ram[133][12] ) );
  DFFHQX1 \ram_reg[133][11]  ( .D(n2721), .CK(clk), .Q(\ram[133][11] ) );
  DFFHQX1 \ram_reg[133][10]  ( .D(n2720), .CK(clk), .Q(\ram[133][10] ) );
  DFFHQX1 \ram_reg[133][9]  ( .D(n2719), .CK(clk), .Q(\ram[133][9] ) );
  DFFHQX1 \ram_reg[133][8]  ( .D(n2718), .CK(clk), .Q(\ram[133][8] ) );
  DFFHQX1 \ram_reg[133][7]  ( .D(n2717), .CK(clk), .Q(\ram[133][7] ) );
  DFFHQX1 \ram_reg[133][6]  ( .D(n2716), .CK(clk), .Q(\ram[133][6] ) );
  DFFHQX1 \ram_reg[133][5]  ( .D(n2715), .CK(clk), .Q(\ram[133][5] ) );
  DFFHQX1 \ram_reg[133][4]  ( .D(n2714), .CK(clk), .Q(\ram[133][4] ) );
  DFFHQX1 \ram_reg[133][3]  ( .D(n2713), .CK(clk), .Q(\ram[133][3] ) );
  DFFHQX1 \ram_reg[133][2]  ( .D(n2712), .CK(clk), .Q(\ram[133][2] ) );
  DFFHQX1 \ram_reg[133][1]  ( .D(n2711), .CK(clk), .Q(\ram[133][1] ) );
  DFFHQX1 \ram_reg[133][0]  ( .D(n2710), .CK(clk), .Q(\ram[133][0] ) );
  DFFHQX1 \ram_reg[129][15]  ( .D(n2661), .CK(clk), .Q(\ram[129][15] ) );
  DFFHQX1 \ram_reg[129][14]  ( .D(n2660), .CK(clk), .Q(\ram[129][14] ) );
  DFFHQX1 \ram_reg[129][13]  ( .D(n2659), .CK(clk), .Q(\ram[129][13] ) );
  DFFHQX1 \ram_reg[129][12]  ( .D(n2658), .CK(clk), .Q(\ram[129][12] ) );
  DFFHQX1 \ram_reg[129][11]  ( .D(n2657), .CK(clk), .Q(\ram[129][11] ) );
  DFFHQX1 \ram_reg[129][10]  ( .D(n2656), .CK(clk), .Q(\ram[129][10] ) );
  DFFHQX1 \ram_reg[129][9]  ( .D(n2655), .CK(clk), .Q(\ram[129][9] ) );
  DFFHQX1 \ram_reg[129][8]  ( .D(n2654), .CK(clk), .Q(\ram[129][8] ) );
  DFFHQX1 \ram_reg[129][7]  ( .D(n2653), .CK(clk), .Q(\ram[129][7] ) );
  DFFHQX1 \ram_reg[129][6]  ( .D(n2652), .CK(clk), .Q(\ram[129][6] ) );
  DFFHQX1 \ram_reg[129][5]  ( .D(n2651), .CK(clk), .Q(\ram[129][5] ) );
  DFFHQX1 \ram_reg[129][4]  ( .D(n2650), .CK(clk), .Q(\ram[129][4] ) );
  DFFHQX1 \ram_reg[129][3]  ( .D(n2649), .CK(clk), .Q(\ram[129][3] ) );
  DFFHQX1 \ram_reg[129][2]  ( .D(n2648), .CK(clk), .Q(\ram[129][2] ) );
  DFFHQX1 \ram_reg[129][1]  ( .D(n2647), .CK(clk), .Q(\ram[129][1] ) );
  DFFHQX1 \ram_reg[129][0]  ( .D(n2646), .CK(clk), .Q(\ram[129][0] ) );
  DFFHQX1 \ram_reg[125][15]  ( .D(n2597), .CK(clk), .Q(\ram[125][15] ) );
  DFFHQX1 \ram_reg[125][14]  ( .D(n2596), .CK(clk), .Q(\ram[125][14] ) );
  DFFHQX1 \ram_reg[125][13]  ( .D(n2595), .CK(clk), .Q(\ram[125][13] ) );
  DFFHQX1 \ram_reg[125][12]  ( .D(n2594), .CK(clk), .Q(\ram[125][12] ) );
  DFFHQX1 \ram_reg[125][11]  ( .D(n2593), .CK(clk), .Q(\ram[125][11] ) );
  DFFHQX1 \ram_reg[125][10]  ( .D(n2592), .CK(clk), .Q(\ram[125][10] ) );
  DFFHQX1 \ram_reg[125][9]  ( .D(n2591), .CK(clk), .Q(\ram[125][9] ) );
  DFFHQX1 \ram_reg[125][8]  ( .D(n2590), .CK(clk), .Q(\ram[125][8] ) );
  DFFHQX1 \ram_reg[125][7]  ( .D(n2589), .CK(clk), .Q(\ram[125][7] ) );
  DFFHQX1 \ram_reg[125][6]  ( .D(n2588), .CK(clk), .Q(\ram[125][6] ) );
  DFFHQX1 \ram_reg[125][5]  ( .D(n2587), .CK(clk), .Q(\ram[125][5] ) );
  DFFHQX1 \ram_reg[125][4]  ( .D(n2586), .CK(clk), .Q(\ram[125][4] ) );
  DFFHQX1 \ram_reg[125][3]  ( .D(n2585), .CK(clk), .Q(\ram[125][3] ) );
  DFFHQX1 \ram_reg[125][2]  ( .D(n2584), .CK(clk), .Q(\ram[125][2] ) );
  DFFHQX1 \ram_reg[125][1]  ( .D(n2583), .CK(clk), .Q(\ram[125][1] ) );
  DFFHQX1 \ram_reg[125][0]  ( .D(n2582), .CK(clk), .Q(\ram[125][0] ) );
  DFFHQX1 \ram_reg[121][15]  ( .D(n2533), .CK(clk), .Q(\ram[121][15] ) );
  DFFHQX1 \ram_reg[121][14]  ( .D(n2532), .CK(clk), .Q(\ram[121][14] ) );
  DFFHQX1 \ram_reg[121][13]  ( .D(n2531), .CK(clk), .Q(\ram[121][13] ) );
  DFFHQX1 \ram_reg[121][12]  ( .D(n2530), .CK(clk), .Q(\ram[121][12] ) );
  DFFHQX1 \ram_reg[121][11]  ( .D(n2529), .CK(clk), .Q(\ram[121][11] ) );
  DFFHQX1 \ram_reg[121][10]  ( .D(n2528), .CK(clk), .Q(\ram[121][10] ) );
  DFFHQX1 \ram_reg[121][9]  ( .D(n2527), .CK(clk), .Q(\ram[121][9] ) );
  DFFHQX1 \ram_reg[121][8]  ( .D(n2526), .CK(clk), .Q(\ram[121][8] ) );
  DFFHQX1 \ram_reg[121][7]  ( .D(n2525), .CK(clk), .Q(\ram[121][7] ) );
  DFFHQX1 \ram_reg[121][6]  ( .D(n2524), .CK(clk), .Q(\ram[121][6] ) );
  DFFHQX1 \ram_reg[121][5]  ( .D(n2523), .CK(clk), .Q(\ram[121][5] ) );
  DFFHQX1 \ram_reg[121][4]  ( .D(n2522), .CK(clk), .Q(\ram[121][4] ) );
  DFFHQX1 \ram_reg[121][3]  ( .D(n2521), .CK(clk), .Q(\ram[121][3] ) );
  DFFHQX1 \ram_reg[121][2]  ( .D(n2520), .CK(clk), .Q(\ram[121][2] ) );
  DFFHQX1 \ram_reg[121][1]  ( .D(n2519), .CK(clk), .Q(\ram[121][1] ) );
  DFFHQX1 \ram_reg[121][0]  ( .D(n2518), .CK(clk), .Q(\ram[121][0] ) );
  DFFHQX1 \ram_reg[117][15]  ( .D(n2469), .CK(clk), .Q(\ram[117][15] ) );
  DFFHQX1 \ram_reg[117][14]  ( .D(n2468), .CK(clk), .Q(\ram[117][14] ) );
  DFFHQX1 \ram_reg[117][13]  ( .D(n2467), .CK(clk), .Q(\ram[117][13] ) );
  DFFHQX1 \ram_reg[117][12]  ( .D(n2466), .CK(clk), .Q(\ram[117][12] ) );
  DFFHQX1 \ram_reg[117][11]  ( .D(n2465), .CK(clk), .Q(\ram[117][11] ) );
  DFFHQX1 \ram_reg[117][10]  ( .D(n2464), .CK(clk), .Q(\ram[117][10] ) );
  DFFHQX1 \ram_reg[117][9]  ( .D(n2463), .CK(clk), .Q(\ram[117][9] ) );
  DFFHQX1 \ram_reg[117][8]  ( .D(n2462), .CK(clk), .Q(\ram[117][8] ) );
  DFFHQX1 \ram_reg[117][7]  ( .D(n2461), .CK(clk), .Q(\ram[117][7] ) );
  DFFHQX1 \ram_reg[117][6]  ( .D(n2460), .CK(clk), .Q(\ram[117][6] ) );
  DFFHQX1 \ram_reg[117][5]  ( .D(n2459), .CK(clk), .Q(\ram[117][5] ) );
  DFFHQX1 \ram_reg[117][4]  ( .D(n2458), .CK(clk), .Q(\ram[117][4] ) );
  DFFHQX1 \ram_reg[117][3]  ( .D(n2457), .CK(clk), .Q(\ram[117][3] ) );
  DFFHQX1 \ram_reg[117][2]  ( .D(n2456), .CK(clk), .Q(\ram[117][2] ) );
  DFFHQX1 \ram_reg[117][1]  ( .D(n2455), .CK(clk), .Q(\ram[117][1] ) );
  DFFHQX1 \ram_reg[117][0]  ( .D(n2454), .CK(clk), .Q(\ram[117][0] ) );
  DFFHQX1 \ram_reg[113][15]  ( .D(n2405), .CK(clk), .Q(\ram[113][15] ) );
  DFFHQX1 \ram_reg[113][14]  ( .D(n2404), .CK(clk), .Q(\ram[113][14] ) );
  DFFHQX1 \ram_reg[113][13]  ( .D(n2403), .CK(clk), .Q(\ram[113][13] ) );
  DFFHQX1 \ram_reg[113][12]  ( .D(n2402), .CK(clk), .Q(\ram[113][12] ) );
  DFFHQX1 \ram_reg[113][11]  ( .D(n2401), .CK(clk), .Q(\ram[113][11] ) );
  DFFHQX1 \ram_reg[113][10]  ( .D(n2400), .CK(clk), .Q(\ram[113][10] ) );
  DFFHQX1 \ram_reg[113][9]  ( .D(n2399), .CK(clk), .Q(\ram[113][9] ) );
  DFFHQX1 \ram_reg[113][8]  ( .D(n2398), .CK(clk), .Q(\ram[113][8] ) );
  DFFHQX1 \ram_reg[113][7]  ( .D(n2397), .CK(clk), .Q(\ram[113][7] ) );
  DFFHQX1 \ram_reg[113][6]  ( .D(n2396), .CK(clk), .Q(\ram[113][6] ) );
  DFFHQX1 \ram_reg[113][5]  ( .D(n2395), .CK(clk), .Q(\ram[113][5] ) );
  DFFHQX1 \ram_reg[113][4]  ( .D(n2394), .CK(clk), .Q(\ram[113][4] ) );
  DFFHQX1 \ram_reg[113][3]  ( .D(n2393), .CK(clk), .Q(\ram[113][3] ) );
  DFFHQX1 \ram_reg[113][2]  ( .D(n2392), .CK(clk), .Q(\ram[113][2] ) );
  DFFHQX1 \ram_reg[113][1]  ( .D(n2391), .CK(clk), .Q(\ram[113][1] ) );
  DFFHQX1 \ram_reg[113][0]  ( .D(n2390), .CK(clk), .Q(\ram[113][0] ) );
  DFFHQX1 \ram_reg[109][15]  ( .D(n2341), .CK(clk), .Q(\ram[109][15] ) );
  DFFHQX1 \ram_reg[109][14]  ( .D(n2340), .CK(clk), .Q(\ram[109][14] ) );
  DFFHQX1 \ram_reg[109][13]  ( .D(n2339), .CK(clk), .Q(\ram[109][13] ) );
  DFFHQX1 \ram_reg[109][12]  ( .D(n2338), .CK(clk), .Q(\ram[109][12] ) );
  DFFHQX1 \ram_reg[109][11]  ( .D(n2337), .CK(clk), .Q(\ram[109][11] ) );
  DFFHQX1 \ram_reg[109][10]  ( .D(n2336), .CK(clk), .Q(\ram[109][10] ) );
  DFFHQX1 \ram_reg[109][9]  ( .D(n2335), .CK(clk), .Q(\ram[109][9] ) );
  DFFHQX1 \ram_reg[109][8]  ( .D(n2334), .CK(clk), .Q(\ram[109][8] ) );
  DFFHQX1 \ram_reg[109][7]  ( .D(n2333), .CK(clk), .Q(\ram[109][7] ) );
  DFFHQX1 \ram_reg[109][6]  ( .D(n2332), .CK(clk), .Q(\ram[109][6] ) );
  DFFHQX1 \ram_reg[109][5]  ( .D(n2331), .CK(clk), .Q(\ram[109][5] ) );
  DFFHQX1 \ram_reg[109][4]  ( .D(n2330), .CK(clk), .Q(\ram[109][4] ) );
  DFFHQX1 \ram_reg[109][3]  ( .D(n2329), .CK(clk), .Q(\ram[109][3] ) );
  DFFHQX1 \ram_reg[109][2]  ( .D(n2328), .CK(clk), .Q(\ram[109][2] ) );
  DFFHQX1 \ram_reg[109][1]  ( .D(n2327), .CK(clk), .Q(\ram[109][1] ) );
  DFFHQX1 \ram_reg[109][0]  ( .D(n2326), .CK(clk), .Q(\ram[109][0] ) );
  DFFHQX1 \ram_reg[105][15]  ( .D(n2277), .CK(clk), .Q(\ram[105][15] ) );
  DFFHQX1 \ram_reg[105][14]  ( .D(n2276), .CK(clk), .Q(\ram[105][14] ) );
  DFFHQX1 \ram_reg[105][13]  ( .D(n2275), .CK(clk), .Q(\ram[105][13] ) );
  DFFHQX1 \ram_reg[105][12]  ( .D(n2274), .CK(clk), .Q(\ram[105][12] ) );
  DFFHQX1 \ram_reg[105][11]  ( .D(n2273), .CK(clk), .Q(\ram[105][11] ) );
  DFFHQX1 \ram_reg[105][10]  ( .D(n2272), .CK(clk), .Q(\ram[105][10] ) );
  DFFHQX1 \ram_reg[105][9]  ( .D(n2271), .CK(clk), .Q(\ram[105][9] ) );
  DFFHQX1 \ram_reg[105][8]  ( .D(n2270), .CK(clk), .Q(\ram[105][8] ) );
  DFFHQX1 \ram_reg[105][7]  ( .D(n2269), .CK(clk), .Q(\ram[105][7] ) );
  DFFHQX1 \ram_reg[105][6]  ( .D(n2268), .CK(clk), .Q(\ram[105][6] ) );
  DFFHQX1 \ram_reg[105][5]  ( .D(n2267), .CK(clk), .Q(\ram[105][5] ) );
  DFFHQX1 \ram_reg[105][4]  ( .D(n2266), .CK(clk), .Q(\ram[105][4] ) );
  DFFHQX1 \ram_reg[105][3]  ( .D(n2265), .CK(clk), .Q(\ram[105][3] ) );
  DFFHQX1 \ram_reg[105][2]  ( .D(n2264), .CK(clk), .Q(\ram[105][2] ) );
  DFFHQX1 \ram_reg[105][1]  ( .D(n2263), .CK(clk), .Q(\ram[105][1] ) );
  DFFHQX1 \ram_reg[105][0]  ( .D(n2262), .CK(clk), .Q(\ram[105][0] ) );
  DFFHQX1 \ram_reg[101][15]  ( .D(n2213), .CK(clk), .Q(\ram[101][15] ) );
  DFFHQX1 \ram_reg[101][14]  ( .D(n2212), .CK(clk), .Q(\ram[101][14] ) );
  DFFHQX1 \ram_reg[101][13]  ( .D(n2211), .CK(clk), .Q(\ram[101][13] ) );
  DFFHQX1 \ram_reg[101][12]  ( .D(n2210), .CK(clk), .Q(\ram[101][12] ) );
  DFFHQX1 \ram_reg[101][11]  ( .D(n2209), .CK(clk), .Q(\ram[101][11] ) );
  DFFHQX1 \ram_reg[101][10]  ( .D(n2208), .CK(clk), .Q(\ram[101][10] ) );
  DFFHQX1 \ram_reg[101][9]  ( .D(n2207), .CK(clk), .Q(\ram[101][9] ) );
  DFFHQX1 \ram_reg[101][8]  ( .D(n2206), .CK(clk), .Q(\ram[101][8] ) );
  DFFHQX1 \ram_reg[101][7]  ( .D(n2205), .CK(clk), .Q(\ram[101][7] ) );
  DFFHQX1 \ram_reg[101][6]  ( .D(n2204), .CK(clk), .Q(\ram[101][6] ) );
  DFFHQX1 \ram_reg[101][5]  ( .D(n2203), .CK(clk), .Q(\ram[101][5] ) );
  DFFHQX1 \ram_reg[101][4]  ( .D(n2202), .CK(clk), .Q(\ram[101][4] ) );
  DFFHQX1 \ram_reg[101][3]  ( .D(n2201), .CK(clk), .Q(\ram[101][3] ) );
  DFFHQX1 \ram_reg[101][2]  ( .D(n2200), .CK(clk), .Q(\ram[101][2] ) );
  DFFHQX1 \ram_reg[101][1]  ( .D(n2199), .CK(clk), .Q(\ram[101][1] ) );
  DFFHQX1 \ram_reg[101][0]  ( .D(n2198), .CK(clk), .Q(\ram[101][0] ) );
  DFFHQX1 \ram_reg[97][15]  ( .D(n2149), .CK(clk), .Q(\ram[97][15] ) );
  DFFHQX1 \ram_reg[97][14]  ( .D(n2148), .CK(clk), .Q(\ram[97][14] ) );
  DFFHQX1 \ram_reg[97][13]  ( .D(n2147), .CK(clk), .Q(\ram[97][13] ) );
  DFFHQX1 \ram_reg[97][12]  ( .D(n2146), .CK(clk), .Q(\ram[97][12] ) );
  DFFHQX1 \ram_reg[97][11]  ( .D(n2145), .CK(clk), .Q(\ram[97][11] ) );
  DFFHQX1 \ram_reg[97][10]  ( .D(n2144), .CK(clk), .Q(\ram[97][10] ) );
  DFFHQX1 \ram_reg[97][9]  ( .D(n2143), .CK(clk), .Q(\ram[97][9] ) );
  DFFHQX1 \ram_reg[97][8]  ( .D(n2142), .CK(clk), .Q(\ram[97][8] ) );
  DFFHQX1 \ram_reg[97][7]  ( .D(n2141), .CK(clk), .Q(\ram[97][7] ) );
  DFFHQX1 \ram_reg[97][6]  ( .D(n2140), .CK(clk), .Q(\ram[97][6] ) );
  DFFHQX1 \ram_reg[97][5]  ( .D(n2139), .CK(clk), .Q(\ram[97][5] ) );
  DFFHQX1 \ram_reg[97][4]  ( .D(n2138), .CK(clk), .Q(\ram[97][4] ) );
  DFFHQX1 \ram_reg[97][3]  ( .D(n2137), .CK(clk), .Q(\ram[97][3] ) );
  DFFHQX1 \ram_reg[97][2]  ( .D(n2136), .CK(clk), .Q(\ram[97][2] ) );
  DFFHQX1 \ram_reg[97][1]  ( .D(n2135), .CK(clk), .Q(\ram[97][1] ) );
  DFFHQX1 \ram_reg[97][0]  ( .D(n2134), .CK(clk), .Q(\ram[97][0] ) );
  DFFHQX1 \ram_reg[93][15]  ( .D(n2085), .CK(clk), .Q(\ram[93][15] ) );
  DFFHQX1 \ram_reg[93][14]  ( .D(n2084), .CK(clk), .Q(\ram[93][14] ) );
  DFFHQX1 \ram_reg[93][13]  ( .D(n2083), .CK(clk), .Q(\ram[93][13] ) );
  DFFHQX1 \ram_reg[93][12]  ( .D(n2082), .CK(clk), .Q(\ram[93][12] ) );
  DFFHQX1 \ram_reg[93][11]  ( .D(n2081), .CK(clk), .Q(\ram[93][11] ) );
  DFFHQX1 \ram_reg[93][10]  ( .D(n2080), .CK(clk), .Q(\ram[93][10] ) );
  DFFHQX1 \ram_reg[93][9]  ( .D(n2079), .CK(clk), .Q(\ram[93][9] ) );
  DFFHQX1 \ram_reg[93][8]  ( .D(n2078), .CK(clk), .Q(\ram[93][8] ) );
  DFFHQX1 \ram_reg[93][7]  ( .D(n2077), .CK(clk), .Q(\ram[93][7] ) );
  DFFHQX1 \ram_reg[93][6]  ( .D(n2076), .CK(clk), .Q(\ram[93][6] ) );
  DFFHQX1 \ram_reg[93][5]  ( .D(n2075), .CK(clk), .Q(\ram[93][5] ) );
  DFFHQX1 \ram_reg[93][4]  ( .D(n2074), .CK(clk), .Q(\ram[93][4] ) );
  DFFHQX1 \ram_reg[93][3]  ( .D(n2073), .CK(clk), .Q(\ram[93][3] ) );
  DFFHQX1 \ram_reg[93][2]  ( .D(n2072), .CK(clk), .Q(\ram[93][2] ) );
  DFFHQX1 \ram_reg[93][1]  ( .D(n2071), .CK(clk), .Q(\ram[93][1] ) );
  DFFHQX1 \ram_reg[93][0]  ( .D(n2070), .CK(clk), .Q(\ram[93][0] ) );
  DFFHQX1 \ram_reg[89][15]  ( .D(n2021), .CK(clk), .Q(\ram[89][15] ) );
  DFFHQX1 \ram_reg[89][14]  ( .D(n2020), .CK(clk), .Q(\ram[89][14] ) );
  DFFHQX1 \ram_reg[89][13]  ( .D(n2019), .CK(clk), .Q(\ram[89][13] ) );
  DFFHQX1 \ram_reg[89][12]  ( .D(n2018), .CK(clk), .Q(\ram[89][12] ) );
  DFFHQX1 \ram_reg[89][11]  ( .D(n2017), .CK(clk), .Q(\ram[89][11] ) );
  DFFHQX1 \ram_reg[89][10]  ( .D(n2016), .CK(clk), .Q(\ram[89][10] ) );
  DFFHQX1 \ram_reg[89][9]  ( .D(n2015), .CK(clk), .Q(\ram[89][9] ) );
  DFFHQX1 \ram_reg[89][8]  ( .D(n2014), .CK(clk), .Q(\ram[89][8] ) );
  DFFHQX1 \ram_reg[89][7]  ( .D(n2013), .CK(clk), .Q(\ram[89][7] ) );
  DFFHQX1 \ram_reg[89][6]  ( .D(n2012), .CK(clk), .Q(\ram[89][6] ) );
  DFFHQX1 \ram_reg[89][5]  ( .D(n2011), .CK(clk), .Q(\ram[89][5] ) );
  DFFHQX1 \ram_reg[89][4]  ( .D(n2010), .CK(clk), .Q(\ram[89][4] ) );
  DFFHQX1 \ram_reg[89][3]  ( .D(n2009), .CK(clk), .Q(\ram[89][3] ) );
  DFFHQX1 \ram_reg[89][2]  ( .D(n2008), .CK(clk), .Q(\ram[89][2] ) );
  DFFHQX1 \ram_reg[89][1]  ( .D(n2007), .CK(clk), .Q(\ram[89][1] ) );
  DFFHQX1 \ram_reg[89][0]  ( .D(n2006), .CK(clk), .Q(\ram[89][0] ) );
  DFFHQX1 \ram_reg[85][15]  ( .D(n1957), .CK(clk), .Q(\ram[85][15] ) );
  DFFHQX1 \ram_reg[85][14]  ( .D(n1956), .CK(clk), .Q(\ram[85][14] ) );
  DFFHQX1 \ram_reg[85][13]  ( .D(n1955), .CK(clk), .Q(\ram[85][13] ) );
  DFFHQX1 \ram_reg[85][12]  ( .D(n1954), .CK(clk), .Q(\ram[85][12] ) );
  DFFHQX1 \ram_reg[85][11]  ( .D(n1953), .CK(clk), .Q(\ram[85][11] ) );
  DFFHQX1 \ram_reg[85][10]  ( .D(n1952), .CK(clk), .Q(\ram[85][10] ) );
  DFFHQX1 \ram_reg[85][9]  ( .D(n1951), .CK(clk), .Q(\ram[85][9] ) );
  DFFHQX1 \ram_reg[85][8]  ( .D(n1950), .CK(clk), .Q(\ram[85][8] ) );
  DFFHQX1 \ram_reg[85][7]  ( .D(n1949), .CK(clk), .Q(\ram[85][7] ) );
  DFFHQX1 \ram_reg[85][6]  ( .D(n1948), .CK(clk), .Q(\ram[85][6] ) );
  DFFHQX1 \ram_reg[85][5]  ( .D(n1947), .CK(clk), .Q(\ram[85][5] ) );
  DFFHQX1 \ram_reg[85][4]  ( .D(n1946), .CK(clk), .Q(\ram[85][4] ) );
  DFFHQX1 \ram_reg[85][3]  ( .D(n1945), .CK(clk), .Q(\ram[85][3] ) );
  DFFHQX1 \ram_reg[85][2]  ( .D(n1944), .CK(clk), .Q(\ram[85][2] ) );
  DFFHQX1 \ram_reg[85][1]  ( .D(n1943), .CK(clk), .Q(\ram[85][1] ) );
  DFFHQX1 \ram_reg[85][0]  ( .D(n1942), .CK(clk), .Q(\ram[85][0] ) );
  DFFHQX1 \ram_reg[81][15]  ( .D(n1893), .CK(clk), .Q(\ram[81][15] ) );
  DFFHQX1 \ram_reg[81][14]  ( .D(n1892), .CK(clk), .Q(\ram[81][14] ) );
  DFFHQX1 \ram_reg[81][13]  ( .D(n1891), .CK(clk), .Q(\ram[81][13] ) );
  DFFHQX1 \ram_reg[81][12]  ( .D(n1890), .CK(clk), .Q(\ram[81][12] ) );
  DFFHQX1 \ram_reg[81][11]  ( .D(n1889), .CK(clk), .Q(\ram[81][11] ) );
  DFFHQX1 \ram_reg[81][10]  ( .D(n1888), .CK(clk), .Q(\ram[81][10] ) );
  DFFHQX1 \ram_reg[81][9]  ( .D(n1887), .CK(clk), .Q(\ram[81][9] ) );
  DFFHQX1 \ram_reg[81][8]  ( .D(n1886), .CK(clk), .Q(\ram[81][8] ) );
  DFFHQX1 \ram_reg[81][7]  ( .D(n1885), .CK(clk), .Q(\ram[81][7] ) );
  DFFHQX1 \ram_reg[81][6]  ( .D(n1884), .CK(clk), .Q(\ram[81][6] ) );
  DFFHQX1 \ram_reg[81][5]  ( .D(n1883), .CK(clk), .Q(\ram[81][5] ) );
  DFFHQX1 \ram_reg[81][4]  ( .D(n1882), .CK(clk), .Q(\ram[81][4] ) );
  DFFHQX1 \ram_reg[81][3]  ( .D(n1881), .CK(clk), .Q(\ram[81][3] ) );
  DFFHQX1 \ram_reg[81][2]  ( .D(n1880), .CK(clk), .Q(\ram[81][2] ) );
  DFFHQX1 \ram_reg[81][1]  ( .D(n1879), .CK(clk), .Q(\ram[81][1] ) );
  DFFHQX1 \ram_reg[81][0]  ( .D(n1878), .CK(clk), .Q(\ram[81][0] ) );
  DFFHQX1 \ram_reg[77][15]  ( .D(n1829), .CK(clk), .Q(\ram[77][15] ) );
  DFFHQX1 \ram_reg[77][14]  ( .D(n1828), .CK(clk), .Q(\ram[77][14] ) );
  DFFHQX1 \ram_reg[77][13]  ( .D(n1827), .CK(clk), .Q(\ram[77][13] ) );
  DFFHQX1 \ram_reg[77][12]  ( .D(n1826), .CK(clk), .Q(\ram[77][12] ) );
  DFFHQX1 \ram_reg[77][11]  ( .D(n1825), .CK(clk), .Q(\ram[77][11] ) );
  DFFHQX1 \ram_reg[77][10]  ( .D(n1824), .CK(clk), .Q(\ram[77][10] ) );
  DFFHQX1 \ram_reg[77][9]  ( .D(n1823), .CK(clk), .Q(\ram[77][9] ) );
  DFFHQX1 \ram_reg[77][8]  ( .D(n1822), .CK(clk), .Q(\ram[77][8] ) );
  DFFHQX1 \ram_reg[77][7]  ( .D(n1821), .CK(clk), .Q(\ram[77][7] ) );
  DFFHQX1 \ram_reg[77][6]  ( .D(n1820), .CK(clk), .Q(\ram[77][6] ) );
  DFFHQX1 \ram_reg[77][5]  ( .D(n1819), .CK(clk), .Q(\ram[77][5] ) );
  DFFHQX1 \ram_reg[77][4]  ( .D(n1818), .CK(clk), .Q(\ram[77][4] ) );
  DFFHQX1 \ram_reg[77][3]  ( .D(n1817), .CK(clk), .Q(\ram[77][3] ) );
  DFFHQX1 \ram_reg[77][2]  ( .D(n1816), .CK(clk), .Q(\ram[77][2] ) );
  DFFHQX1 \ram_reg[77][1]  ( .D(n1815), .CK(clk), .Q(\ram[77][1] ) );
  DFFHQX1 \ram_reg[77][0]  ( .D(n1814), .CK(clk), .Q(\ram[77][0] ) );
  DFFHQX1 \ram_reg[73][15]  ( .D(n1765), .CK(clk), .Q(\ram[73][15] ) );
  DFFHQX1 \ram_reg[73][14]  ( .D(n1764), .CK(clk), .Q(\ram[73][14] ) );
  DFFHQX1 \ram_reg[73][13]  ( .D(n1763), .CK(clk), .Q(\ram[73][13] ) );
  DFFHQX1 \ram_reg[73][12]  ( .D(n1762), .CK(clk), .Q(\ram[73][12] ) );
  DFFHQX1 \ram_reg[73][11]  ( .D(n1761), .CK(clk), .Q(\ram[73][11] ) );
  DFFHQX1 \ram_reg[73][10]  ( .D(n1760), .CK(clk), .Q(\ram[73][10] ) );
  DFFHQX1 \ram_reg[73][9]  ( .D(n1759), .CK(clk), .Q(\ram[73][9] ) );
  DFFHQX1 \ram_reg[73][8]  ( .D(n1758), .CK(clk), .Q(\ram[73][8] ) );
  DFFHQX1 \ram_reg[73][7]  ( .D(n1757), .CK(clk), .Q(\ram[73][7] ) );
  DFFHQX1 \ram_reg[73][6]  ( .D(n1756), .CK(clk), .Q(\ram[73][6] ) );
  DFFHQX1 \ram_reg[73][5]  ( .D(n1755), .CK(clk), .Q(\ram[73][5] ) );
  DFFHQX1 \ram_reg[73][4]  ( .D(n1754), .CK(clk), .Q(\ram[73][4] ) );
  DFFHQX1 \ram_reg[73][3]  ( .D(n1753), .CK(clk), .Q(\ram[73][3] ) );
  DFFHQX1 \ram_reg[73][2]  ( .D(n1752), .CK(clk), .Q(\ram[73][2] ) );
  DFFHQX1 \ram_reg[73][1]  ( .D(n1751), .CK(clk), .Q(\ram[73][1] ) );
  DFFHQX1 \ram_reg[73][0]  ( .D(n1750), .CK(clk), .Q(\ram[73][0] ) );
  DFFHQX1 \ram_reg[69][15]  ( .D(n1701), .CK(clk), .Q(\ram[69][15] ) );
  DFFHQX1 \ram_reg[69][14]  ( .D(n1700), .CK(clk), .Q(\ram[69][14] ) );
  DFFHQX1 \ram_reg[69][13]  ( .D(n1699), .CK(clk), .Q(\ram[69][13] ) );
  DFFHQX1 \ram_reg[69][12]  ( .D(n1698), .CK(clk), .Q(\ram[69][12] ) );
  DFFHQX1 \ram_reg[69][11]  ( .D(n1697), .CK(clk), .Q(\ram[69][11] ) );
  DFFHQX1 \ram_reg[69][10]  ( .D(n1696), .CK(clk), .Q(\ram[69][10] ) );
  DFFHQX1 \ram_reg[69][9]  ( .D(n1695), .CK(clk), .Q(\ram[69][9] ) );
  DFFHQX1 \ram_reg[69][8]  ( .D(n1694), .CK(clk), .Q(\ram[69][8] ) );
  DFFHQX1 \ram_reg[69][7]  ( .D(n1693), .CK(clk), .Q(\ram[69][7] ) );
  DFFHQX1 \ram_reg[69][6]  ( .D(n1692), .CK(clk), .Q(\ram[69][6] ) );
  DFFHQX1 \ram_reg[69][5]  ( .D(n1691), .CK(clk), .Q(\ram[69][5] ) );
  DFFHQX1 \ram_reg[69][4]  ( .D(n1690), .CK(clk), .Q(\ram[69][4] ) );
  DFFHQX1 \ram_reg[69][3]  ( .D(n1689), .CK(clk), .Q(\ram[69][3] ) );
  DFFHQX1 \ram_reg[69][2]  ( .D(n1688), .CK(clk), .Q(\ram[69][2] ) );
  DFFHQX1 \ram_reg[69][1]  ( .D(n1687), .CK(clk), .Q(\ram[69][1] ) );
  DFFHQX1 \ram_reg[69][0]  ( .D(n1686), .CK(clk), .Q(\ram[69][0] ) );
  DFFHQX1 \ram_reg[65][15]  ( .D(n1637), .CK(clk), .Q(\ram[65][15] ) );
  DFFHQX1 \ram_reg[65][14]  ( .D(n1636), .CK(clk), .Q(\ram[65][14] ) );
  DFFHQX1 \ram_reg[65][13]  ( .D(n1635), .CK(clk), .Q(\ram[65][13] ) );
  DFFHQX1 \ram_reg[65][12]  ( .D(n1634), .CK(clk), .Q(\ram[65][12] ) );
  DFFHQX1 \ram_reg[65][11]  ( .D(n1633), .CK(clk), .Q(\ram[65][11] ) );
  DFFHQX1 \ram_reg[65][10]  ( .D(n1632), .CK(clk), .Q(\ram[65][10] ) );
  DFFHQX1 \ram_reg[65][9]  ( .D(n1631), .CK(clk), .Q(\ram[65][9] ) );
  DFFHQX1 \ram_reg[65][8]  ( .D(n1630), .CK(clk), .Q(\ram[65][8] ) );
  DFFHQX1 \ram_reg[65][7]  ( .D(n1629), .CK(clk), .Q(\ram[65][7] ) );
  DFFHQX1 \ram_reg[65][6]  ( .D(n1628), .CK(clk), .Q(\ram[65][6] ) );
  DFFHQX1 \ram_reg[65][5]  ( .D(n1627), .CK(clk), .Q(\ram[65][5] ) );
  DFFHQX1 \ram_reg[65][4]  ( .D(n1626), .CK(clk), .Q(\ram[65][4] ) );
  DFFHQX1 \ram_reg[65][3]  ( .D(n1625), .CK(clk), .Q(\ram[65][3] ) );
  DFFHQX1 \ram_reg[65][2]  ( .D(n1624), .CK(clk), .Q(\ram[65][2] ) );
  DFFHQX1 \ram_reg[65][1]  ( .D(n1623), .CK(clk), .Q(\ram[65][1] ) );
  DFFHQX1 \ram_reg[65][0]  ( .D(n1622), .CK(clk), .Q(\ram[65][0] ) );
  DFFHQX1 \ram_reg[61][15]  ( .D(n1573), .CK(clk), .Q(\ram[61][15] ) );
  DFFHQX1 \ram_reg[61][14]  ( .D(n1572), .CK(clk), .Q(\ram[61][14] ) );
  DFFHQX1 \ram_reg[61][13]  ( .D(n1571), .CK(clk), .Q(\ram[61][13] ) );
  DFFHQX1 \ram_reg[61][12]  ( .D(n1570), .CK(clk), .Q(\ram[61][12] ) );
  DFFHQX1 \ram_reg[61][11]  ( .D(n1569), .CK(clk), .Q(\ram[61][11] ) );
  DFFHQX1 \ram_reg[61][10]  ( .D(n1568), .CK(clk), .Q(\ram[61][10] ) );
  DFFHQX1 \ram_reg[61][9]  ( .D(n1567), .CK(clk), .Q(\ram[61][9] ) );
  DFFHQX1 \ram_reg[61][8]  ( .D(n1566), .CK(clk), .Q(\ram[61][8] ) );
  DFFHQX1 \ram_reg[61][7]  ( .D(n1565), .CK(clk), .Q(\ram[61][7] ) );
  DFFHQX1 \ram_reg[61][6]  ( .D(n1564), .CK(clk), .Q(\ram[61][6] ) );
  DFFHQX1 \ram_reg[61][5]  ( .D(n1563), .CK(clk), .Q(\ram[61][5] ) );
  DFFHQX1 \ram_reg[61][4]  ( .D(n1562), .CK(clk), .Q(\ram[61][4] ) );
  DFFHQX1 \ram_reg[61][3]  ( .D(n1561), .CK(clk), .Q(\ram[61][3] ) );
  DFFHQX1 \ram_reg[61][2]  ( .D(n1560), .CK(clk), .Q(\ram[61][2] ) );
  DFFHQX1 \ram_reg[61][1]  ( .D(n1559), .CK(clk), .Q(\ram[61][1] ) );
  DFFHQX1 \ram_reg[61][0]  ( .D(n1558), .CK(clk), .Q(\ram[61][0] ) );
  DFFHQX1 \ram_reg[57][15]  ( .D(n1509), .CK(clk), .Q(\ram[57][15] ) );
  DFFHQX1 \ram_reg[57][14]  ( .D(n1508), .CK(clk), .Q(\ram[57][14] ) );
  DFFHQX1 \ram_reg[57][13]  ( .D(n1507), .CK(clk), .Q(\ram[57][13] ) );
  DFFHQX1 \ram_reg[57][12]  ( .D(n1506), .CK(clk), .Q(\ram[57][12] ) );
  DFFHQX1 \ram_reg[57][11]  ( .D(n1505), .CK(clk), .Q(\ram[57][11] ) );
  DFFHQX1 \ram_reg[57][10]  ( .D(n1504), .CK(clk), .Q(\ram[57][10] ) );
  DFFHQX1 \ram_reg[57][9]  ( .D(n1503), .CK(clk), .Q(\ram[57][9] ) );
  DFFHQX1 \ram_reg[57][8]  ( .D(n1502), .CK(clk), .Q(\ram[57][8] ) );
  DFFHQX1 \ram_reg[57][7]  ( .D(n1501), .CK(clk), .Q(\ram[57][7] ) );
  DFFHQX1 \ram_reg[57][6]  ( .D(n1500), .CK(clk), .Q(\ram[57][6] ) );
  DFFHQX1 \ram_reg[57][5]  ( .D(n1499), .CK(clk), .Q(\ram[57][5] ) );
  DFFHQX1 \ram_reg[57][4]  ( .D(n1498), .CK(clk), .Q(\ram[57][4] ) );
  DFFHQX1 \ram_reg[57][3]  ( .D(n1497), .CK(clk), .Q(\ram[57][3] ) );
  DFFHQX1 \ram_reg[57][2]  ( .D(n1496), .CK(clk), .Q(\ram[57][2] ) );
  DFFHQX1 \ram_reg[57][1]  ( .D(n1495), .CK(clk), .Q(\ram[57][1] ) );
  DFFHQX1 \ram_reg[57][0]  ( .D(n1494), .CK(clk), .Q(\ram[57][0] ) );
  DFFHQX1 \ram_reg[53][15]  ( .D(n1445), .CK(clk), .Q(\ram[53][15] ) );
  DFFHQX1 \ram_reg[53][14]  ( .D(n1444), .CK(clk), .Q(\ram[53][14] ) );
  DFFHQX1 \ram_reg[53][13]  ( .D(n1443), .CK(clk), .Q(\ram[53][13] ) );
  DFFHQX1 \ram_reg[53][12]  ( .D(n1442), .CK(clk), .Q(\ram[53][12] ) );
  DFFHQX1 \ram_reg[53][11]  ( .D(n1441), .CK(clk), .Q(\ram[53][11] ) );
  DFFHQX1 \ram_reg[53][10]  ( .D(n1440), .CK(clk), .Q(\ram[53][10] ) );
  DFFHQX1 \ram_reg[53][9]  ( .D(n1439), .CK(clk), .Q(\ram[53][9] ) );
  DFFHQX1 \ram_reg[53][8]  ( .D(n1438), .CK(clk), .Q(\ram[53][8] ) );
  DFFHQX1 \ram_reg[53][7]  ( .D(n1437), .CK(clk), .Q(\ram[53][7] ) );
  DFFHQX1 \ram_reg[53][6]  ( .D(n1436), .CK(clk), .Q(\ram[53][6] ) );
  DFFHQX1 \ram_reg[53][5]  ( .D(n1435), .CK(clk), .Q(\ram[53][5] ) );
  DFFHQX1 \ram_reg[53][4]  ( .D(n1434), .CK(clk), .Q(\ram[53][4] ) );
  DFFHQX1 \ram_reg[53][3]  ( .D(n1433), .CK(clk), .Q(\ram[53][3] ) );
  DFFHQX1 \ram_reg[53][2]  ( .D(n1432), .CK(clk), .Q(\ram[53][2] ) );
  DFFHQX1 \ram_reg[53][1]  ( .D(n1431), .CK(clk), .Q(\ram[53][1] ) );
  DFFHQX1 \ram_reg[53][0]  ( .D(n1430), .CK(clk), .Q(\ram[53][0] ) );
  DFFHQX1 \ram_reg[49][15]  ( .D(n1381), .CK(clk), .Q(\ram[49][15] ) );
  DFFHQX1 \ram_reg[49][14]  ( .D(n1380), .CK(clk), .Q(\ram[49][14] ) );
  DFFHQX1 \ram_reg[49][13]  ( .D(n1379), .CK(clk), .Q(\ram[49][13] ) );
  DFFHQX1 \ram_reg[49][12]  ( .D(n1378), .CK(clk), .Q(\ram[49][12] ) );
  DFFHQX1 \ram_reg[49][11]  ( .D(n1377), .CK(clk), .Q(\ram[49][11] ) );
  DFFHQX1 \ram_reg[49][10]  ( .D(n1376), .CK(clk), .Q(\ram[49][10] ) );
  DFFHQX1 \ram_reg[49][9]  ( .D(n1375), .CK(clk), .Q(\ram[49][9] ) );
  DFFHQX1 \ram_reg[49][8]  ( .D(n1374), .CK(clk), .Q(\ram[49][8] ) );
  DFFHQX1 \ram_reg[49][7]  ( .D(n1373), .CK(clk), .Q(\ram[49][7] ) );
  DFFHQX1 \ram_reg[49][6]  ( .D(n1372), .CK(clk), .Q(\ram[49][6] ) );
  DFFHQX1 \ram_reg[49][5]  ( .D(n1371), .CK(clk), .Q(\ram[49][5] ) );
  DFFHQX1 \ram_reg[49][4]  ( .D(n1370), .CK(clk), .Q(\ram[49][4] ) );
  DFFHQX1 \ram_reg[49][3]  ( .D(n1369), .CK(clk), .Q(\ram[49][3] ) );
  DFFHQX1 \ram_reg[49][2]  ( .D(n1368), .CK(clk), .Q(\ram[49][2] ) );
  DFFHQX1 \ram_reg[49][1]  ( .D(n1367), .CK(clk), .Q(\ram[49][1] ) );
  DFFHQX1 \ram_reg[49][0]  ( .D(n1366), .CK(clk), .Q(\ram[49][0] ) );
  DFFHQX1 \ram_reg[45][15]  ( .D(n1317), .CK(clk), .Q(\ram[45][15] ) );
  DFFHQX1 \ram_reg[45][14]  ( .D(n1316), .CK(clk), .Q(\ram[45][14] ) );
  DFFHQX1 \ram_reg[45][13]  ( .D(n1315), .CK(clk), .Q(\ram[45][13] ) );
  DFFHQX1 \ram_reg[45][12]  ( .D(n1314), .CK(clk), .Q(\ram[45][12] ) );
  DFFHQX1 \ram_reg[45][11]  ( .D(n1313), .CK(clk), .Q(\ram[45][11] ) );
  DFFHQX1 \ram_reg[45][10]  ( .D(n1312), .CK(clk), .Q(\ram[45][10] ) );
  DFFHQX1 \ram_reg[45][9]  ( .D(n1311), .CK(clk), .Q(\ram[45][9] ) );
  DFFHQX1 \ram_reg[45][8]  ( .D(n1310), .CK(clk), .Q(\ram[45][8] ) );
  DFFHQX1 \ram_reg[45][7]  ( .D(n1309), .CK(clk), .Q(\ram[45][7] ) );
  DFFHQX1 \ram_reg[45][6]  ( .D(n1308), .CK(clk), .Q(\ram[45][6] ) );
  DFFHQX1 \ram_reg[45][5]  ( .D(n1307), .CK(clk), .Q(\ram[45][5] ) );
  DFFHQX1 \ram_reg[45][4]  ( .D(n1306), .CK(clk), .Q(\ram[45][4] ) );
  DFFHQX1 \ram_reg[45][3]  ( .D(n1305), .CK(clk), .Q(\ram[45][3] ) );
  DFFHQX1 \ram_reg[45][2]  ( .D(n1304), .CK(clk), .Q(\ram[45][2] ) );
  DFFHQX1 \ram_reg[45][1]  ( .D(n1303), .CK(clk), .Q(\ram[45][1] ) );
  DFFHQX1 \ram_reg[45][0]  ( .D(n1302), .CK(clk), .Q(\ram[45][0] ) );
  DFFHQX1 \ram_reg[41][15]  ( .D(n1253), .CK(clk), .Q(\ram[41][15] ) );
  DFFHQX1 \ram_reg[41][14]  ( .D(n1252), .CK(clk), .Q(\ram[41][14] ) );
  DFFHQX1 \ram_reg[41][13]  ( .D(n1251), .CK(clk), .Q(\ram[41][13] ) );
  DFFHQX1 \ram_reg[41][12]  ( .D(n1250), .CK(clk), .Q(\ram[41][12] ) );
  DFFHQX1 \ram_reg[41][11]  ( .D(n1249), .CK(clk), .Q(\ram[41][11] ) );
  DFFHQX1 \ram_reg[41][10]  ( .D(n1248), .CK(clk), .Q(\ram[41][10] ) );
  DFFHQX1 \ram_reg[41][9]  ( .D(n1247), .CK(clk), .Q(\ram[41][9] ) );
  DFFHQX1 \ram_reg[41][8]  ( .D(n1246), .CK(clk), .Q(\ram[41][8] ) );
  DFFHQX1 \ram_reg[41][7]  ( .D(n1245), .CK(clk), .Q(\ram[41][7] ) );
  DFFHQX1 \ram_reg[41][6]  ( .D(n1244), .CK(clk), .Q(\ram[41][6] ) );
  DFFHQX1 \ram_reg[41][5]  ( .D(n1243), .CK(clk), .Q(\ram[41][5] ) );
  DFFHQX1 \ram_reg[41][4]  ( .D(n1242), .CK(clk), .Q(\ram[41][4] ) );
  DFFHQX1 \ram_reg[41][3]  ( .D(n1241), .CK(clk), .Q(\ram[41][3] ) );
  DFFHQX1 \ram_reg[41][2]  ( .D(n1240), .CK(clk), .Q(\ram[41][2] ) );
  DFFHQX1 \ram_reg[41][1]  ( .D(n1239), .CK(clk), .Q(\ram[41][1] ) );
  DFFHQX1 \ram_reg[41][0]  ( .D(n1238), .CK(clk), .Q(\ram[41][0] ) );
  DFFHQX1 \ram_reg[37][15]  ( .D(n1189), .CK(clk), .Q(\ram[37][15] ) );
  DFFHQX1 \ram_reg[37][14]  ( .D(n1188), .CK(clk), .Q(\ram[37][14] ) );
  DFFHQX1 \ram_reg[37][13]  ( .D(n1187), .CK(clk), .Q(\ram[37][13] ) );
  DFFHQX1 \ram_reg[37][12]  ( .D(n1186), .CK(clk), .Q(\ram[37][12] ) );
  DFFHQX1 \ram_reg[37][11]  ( .D(n1185), .CK(clk), .Q(\ram[37][11] ) );
  DFFHQX1 \ram_reg[37][10]  ( .D(n1184), .CK(clk), .Q(\ram[37][10] ) );
  DFFHQX1 \ram_reg[37][9]  ( .D(n1183), .CK(clk), .Q(\ram[37][9] ) );
  DFFHQX1 \ram_reg[37][8]  ( .D(n1182), .CK(clk), .Q(\ram[37][8] ) );
  DFFHQX1 \ram_reg[37][7]  ( .D(n1181), .CK(clk), .Q(\ram[37][7] ) );
  DFFHQX1 \ram_reg[37][6]  ( .D(n1180), .CK(clk), .Q(\ram[37][6] ) );
  DFFHQX1 \ram_reg[37][5]  ( .D(n1179), .CK(clk), .Q(\ram[37][5] ) );
  DFFHQX1 \ram_reg[37][4]  ( .D(n1178), .CK(clk), .Q(\ram[37][4] ) );
  DFFHQX1 \ram_reg[37][3]  ( .D(n1177), .CK(clk), .Q(\ram[37][3] ) );
  DFFHQX1 \ram_reg[37][2]  ( .D(n1176), .CK(clk), .Q(\ram[37][2] ) );
  DFFHQX1 \ram_reg[37][1]  ( .D(n1175), .CK(clk), .Q(\ram[37][1] ) );
  DFFHQX1 \ram_reg[37][0]  ( .D(n1174), .CK(clk), .Q(\ram[37][0] ) );
  DFFHQX1 \ram_reg[33][15]  ( .D(n1125), .CK(clk), .Q(\ram[33][15] ) );
  DFFHQX1 \ram_reg[33][14]  ( .D(n1124), .CK(clk), .Q(\ram[33][14] ) );
  DFFHQX1 \ram_reg[33][13]  ( .D(n1123), .CK(clk), .Q(\ram[33][13] ) );
  DFFHQX1 \ram_reg[33][12]  ( .D(n1122), .CK(clk), .Q(\ram[33][12] ) );
  DFFHQX1 \ram_reg[33][11]  ( .D(n1121), .CK(clk), .Q(\ram[33][11] ) );
  DFFHQX1 \ram_reg[33][10]  ( .D(n1120), .CK(clk), .Q(\ram[33][10] ) );
  DFFHQX1 \ram_reg[33][9]  ( .D(n1119), .CK(clk), .Q(\ram[33][9] ) );
  DFFHQX1 \ram_reg[33][8]  ( .D(n1118), .CK(clk), .Q(\ram[33][8] ) );
  DFFHQX1 \ram_reg[33][7]  ( .D(n1117), .CK(clk), .Q(\ram[33][7] ) );
  DFFHQX1 \ram_reg[33][6]  ( .D(n1116), .CK(clk), .Q(\ram[33][6] ) );
  DFFHQX1 \ram_reg[33][5]  ( .D(n1115), .CK(clk), .Q(\ram[33][5] ) );
  DFFHQX1 \ram_reg[33][4]  ( .D(n1114), .CK(clk), .Q(\ram[33][4] ) );
  DFFHQX1 \ram_reg[33][3]  ( .D(n1113), .CK(clk), .Q(\ram[33][3] ) );
  DFFHQX1 \ram_reg[33][2]  ( .D(n1112), .CK(clk), .Q(\ram[33][2] ) );
  DFFHQX1 \ram_reg[33][1]  ( .D(n1111), .CK(clk), .Q(\ram[33][1] ) );
  DFFHQX1 \ram_reg[33][0]  ( .D(n1110), .CK(clk), .Q(\ram[33][0] ) );
  DFFHQX1 \ram_reg[29][15]  ( .D(n1061), .CK(clk), .Q(\ram[29][15] ) );
  DFFHQX1 \ram_reg[29][14]  ( .D(n1060), .CK(clk), .Q(\ram[29][14] ) );
  DFFHQX1 \ram_reg[29][13]  ( .D(n1059), .CK(clk), .Q(\ram[29][13] ) );
  DFFHQX1 \ram_reg[29][12]  ( .D(n1058), .CK(clk), .Q(\ram[29][12] ) );
  DFFHQX1 \ram_reg[29][11]  ( .D(n1057), .CK(clk), .Q(\ram[29][11] ) );
  DFFHQX1 \ram_reg[29][10]  ( .D(n1056), .CK(clk), .Q(\ram[29][10] ) );
  DFFHQX1 \ram_reg[29][9]  ( .D(n1055), .CK(clk), .Q(\ram[29][9] ) );
  DFFHQX1 \ram_reg[29][8]  ( .D(n1054), .CK(clk), .Q(\ram[29][8] ) );
  DFFHQX1 \ram_reg[29][7]  ( .D(n1053), .CK(clk), .Q(\ram[29][7] ) );
  DFFHQX1 \ram_reg[29][6]  ( .D(n1052), .CK(clk), .Q(\ram[29][6] ) );
  DFFHQX1 \ram_reg[29][5]  ( .D(n1051), .CK(clk), .Q(\ram[29][5] ) );
  DFFHQX1 \ram_reg[29][4]  ( .D(n1050), .CK(clk), .Q(\ram[29][4] ) );
  DFFHQX1 \ram_reg[29][3]  ( .D(n1049), .CK(clk), .Q(\ram[29][3] ) );
  DFFHQX1 \ram_reg[29][2]  ( .D(n1048), .CK(clk), .Q(\ram[29][2] ) );
  DFFHQX1 \ram_reg[29][1]  ( .D(n1047), .CK(clk), .Q(\ram[29][1] ) );
  DFFHQX1 \ram_reg[29][0]  ( .D(n1046), .CK(clk), .Q(\ram[29][0] ) );
  DFFHQX1 \ram_reg[25][15]  ( .D(n997), .CK(clk), .Q(\ram[25][15] ) );
  DFFHQX1 \ram_reg[25][14]  ( .D(n996), .CK(clk), .Q(\ram[25][14] ) );
  DFFHQX1 \ram_reg[25][13]  ( .D(n995), .CK(clk), .Q(\ram[25][13] ) );
  DFFHQX1 \ram_reg[25][12]  ( .D(n994), .CK(clk), .Q(\ram[25][12] ) );
  DFFHQX1 \ram_reg[25][11]  ( .D(n993), .CK(clk), .Q(\ram[25][11] ) );
  DFFHQX1 \ram_reg[25][10]  ( .D(n992), .CK(clk), .Q(\ram[25][10] ) );
  DFFHQX1 \ram_reg[25][9]  ( .D(n991), .CK(clk), .Q(\ram[25][9] ) );
  DFFHQX1 \ram_reg[25][8]  ( .D(n990), .CK(clk), .Q(\ram[25][8] ) );
  DFFHQX1 \ram_reg[25][7]  ( .D(n989), .CK(clk), .Q(\ram[25][7] ) );
  DFFHQX1 \ram_reg[25][6]  ( .D(n988), .CK(clk), .Q(\ram[25][6] ) );
  DFFHQX1 \ram_reg[25][5]  ( .D(n987), .CK(clk), .Q(\ram[25][5] ) );
  DFFHQX1 \ram_reg[25][4]  ( .D(n986), .CK(clk), .Q(\ram[25][4] ) );
  DFFHQX1 \ram_reg[25][3]  ( .D(n985), .CK(clk), .Q(\ram[25][3] ) );
  DFFHQX1 \ram_reg[25][2]  ( .D(n984), .CK(clk), .Q(\ram[25][2] ) );
  DFFHQX1 \ram_reg[25][1]  ( .D(n983), .CK(clk), .Q(\ram[25][1] ) );
  DFFHQX1 \ram_reg[25][0]  ( .D(n982), .CK(clk), .Q(\ram[25][0] ) );
  DFFHQX1 \ram_reg[21][15]  ( .D(n933), .CK(clk), .Q(\ram[21][15] ) );
  DFFHQX1 \ram_reg[21][14]  ( .D(n932), .CK(clk), .Q(\ram[21][14] ) );
  DFFHQX1 \ram_reg[21][13]  ( .D(n931), .CK(clk), .Q(\ram[21][13] ) );
  DFFHQX1 \ram_reg[21][12]  ( .D(n930), .CK(clk), .Q(\ram[21][12] ) );
  DFFHQX1 \ram_reg[21][11]  ( .D(n929), .CK(clk), .Q(\ram[21][11] ) );
  DFFHQX1 \ram_reg[21][10]  ( .D(n928), .CK(clk), .Q(\ram[21][10] ) );
  DFFHQX1 \ram_reg[21][9]  ( .D(n927), .CK(clk), .Q(\ram[21][9] ) );
  DFFHQX1 \ram_reg[21][8]  ( .D(n926), .CK(clk), .Q(\ram[21][8] ) );
  DFFHQX1 \ram_reg[21][7]  ( .D(n925), .CK(clk), .Q(\ram[21][7] ) );
  DFFHQX1 \ram_reg[21][6]  ( .D(n924), .CK(clk), .Q(\ram[21][6] ) );
  DFFHQX1 \ram_reg[21][5]  ( .D(n923), .CK(clk), .Q(\ram[21][5] ) );
  DFFHQX1 \ram_reg[21][4]  ( .D(n922), .CK(clk), .Q(\ram[21][4] ) );
  DFFHQX1 \ram_reg[21][3]  ( .D(n921), .CK(clk), .Q(\ram[21][3] ) );
  DFFHQX1 \ram_reg[21][2]  ( .D(n920), .CK(clk), .Q(\ram[21][2] ) );
  DFFHQX1 \ram_reg[21][1]  ( .D(n919), .CK(clk), .Q(\ram[21][1] ) );
  DFFHQX1 \ram_reg[21][0]  ( .D(n918), .CK(clk), .Q(\ram[21][0] ) );
  DFFHQX1 \ram_reg[17][15]  ( .D(n869), .CK(clk), .Q(\ram[17][15] ) );
  DFFHQX1 \ram_reg[17][14]  ( .D(n868), .CK(clk), .Q(\ram[17][14] ) );
  DFFHQX1 \ram_reg[17][13]  ( .D(n867), .CK(clk), .Q(\ram[17][13] ) );
  DFFHQX1 \ram_reg[17][12]  ( .D(n866), .CK(clk), .Q(\ram[17][12] ) );
  DFFHQX1 \ram_reg[17][11]  ( .D(n865), .CK(clk), .Q(\ram[17][11] ) );
  DFFHQX1 \ram_reg[17][10]  ( .D(n864), .CK(clk), .Q(\ram[17][10] ) );
  DFFHQX1 \ram_reg[17][9]  ( .D(n863), .CK(clk), .Q(\ram[17][9] ) );
  DFFHQX1 \ram_reg[17][8]  ( .D(n862), .CK(clk), .Q(\ram[17][8] ) );
  DFFHQX1 \ram_reg[17][7]  ( .D(n861), .CK(clk), .Q(\ram[17][7] ) );
  DFFHQX1 \ram_reg[17][6]  ( .D(n860), .CK(clk), .Q(\ram[17][6] ) );
  DFFHQX1 \ram_reg[17][5]  ( .D(n859), .CK(clk), .Q(\ram[17][5] ) );
  DFFHQX1 \ram_reg[17][4]  ( .D(n858), .CK(clk), .Q(\ram[17][4] ) );
  DFFHQX1 \ram_reg[17][3]  ( .D(n857), .CK(clk), .Q(\ram[17][3] ) );
  DFFHQX1 \ram_reg[17][2]  ( .D(n856), .CK(clk), .Q(\ram[17][2] ) );
  DFFHQX1 \ram_reg[17][1]  ( .D(n855), .CK(clk), .Q(\ram[17][1] ) );
  DFFHQX1 \ram_reg[17][0]  ( .D(n854), .CK(clk), .Q(\ram[17][0] ) );
  DFFHQX1 \ram_reg[13][15]  ( .D(n805), .CK(clk), .Q(\ram[13][15] ) );
  DFFHQX1 \ram_reg[13][14]  ( .D(n804), .CK(clk), .Q(\ram[13][14] ) );
  DFFHQX1 \ram_reg[13][13]  ( .D(n803), .CK(clk), .Q(\ram[13][13] ) );
  DFFHQX1 \ram_reg[13][12]  ( .D(n802), .CK(clk), .Q(\ram[13][12] ) );
  DFFHQX1 \ram_reg[13][11]  ( .D(n801), .CK(clk), .Q(\ram[13][11] ) );
  DFFHQX1 \ram_reg[13][10]  ( .D(n800), .CK(clk), .Q(\ram[13][10] ) );
  DFFHQX1 \ram_reg[13][9]  ( .D(n799), .CK(clk), .Q(\ram[13][9] ) );
  DFFHQX1 \ram_reg[13][8]  ( .D(n798), .CK(clk), .Q(\ram[13][8] ) );
  DFFHQX1 \ram_reg[13][7]  ( .D(n797), .CK(clk), .Q(\ram[13][7] ) );
  DFFHQX1 \ram_reg[13][6]  ( .D(n796), .CK(clk), .Q(\ram[13][6] ) );
  DFFHQX1 \ram_reg[13][5]  ( .D(n795), .CK(clk), .Q(\ram[13][5] ) );
  DFFHQX1 \ram_reg[13][4]  ( .D(n794), .CK(clk), .Q(\ram[13][4] ) );
  DFFHQX1 \ram_reg[13][3]  ( .D(n793), .CK(clk), .Q(\ram[13][3] ) );
  DFFHQX1 \ram_reg[13][2]  ( .D(n792), .CK(clk), .Q(\ram[13][2] ) );
  DFFHQX1 \ram_reg[13][1]  ( .D(n791), .CK(clk), .Q(\ram[13][1] ) );
  DFFHQX1 \ram_reg[13][0]  ( .D(n790), .CK(clk), .Q(\ram[13][0] ) );
  DFFHQX1 \ram_reg[9][15]  ( .D(n741), .CK(clk), .Q(\ram[9][15] ) );
  DFFHQX1 \ram_reg[9][14]  ( .D(n740), .CK(clk), .Q(\ram[9][14] ) );
  DFFHQX1 \ram_reg[9][13]  ( .D(n739), .CK(clk), .Q(\ram[9][13] ) );
  DFFHQX1 \ram_reg[9][12]  ( .D(n738), .CK(clk), .Q(\ram[9][12] ) );
  DFFHQX1 \ram_reg[9][11]  ( .D(n737), .CK(clk), .Q(\ram[9][11] ) );
  DFFHQX1 \ram_reg[9][10]  ( .D(n736), .CK(clk), .Q(\ram[9][10] ) );
  DFFHQX1 \ram_reg[9][9]  ( .D(n735), .CK(clk), .Q(\ram[9][9] ) );
  DFFHQX1 \ram_reg[9][8]  ( .D(n734), .CK(clk), .Q(\ram[9][8] ) );
  DFFHQX1 \ram_reg[9][7]  ( .D(n733), .CK(clk), .Q(\ram[9][7] ) );
  DFFHQX1 \ram_reg[9][6]  ( .D(n732), .CK(clk), .Q(\ram[9][6] ) );
  DFFHQX1 \ram_reg[9][5]  ( .D(n731), .CK(clk), .Q(\ram[9][5] ) );
  DFFHQX1 \ram_reg[9][4]  ( .D(n730), .CK(clk), .Q(\ram[9][4] ) );
  DFFHQX1 \ram_reg[9][3]  ( .D(n729), .CK(clk), .Q(\ram[9][3] ) );
  DFFHQX1 \ram_reg[9][2]  ( .D(n728), .CK(clk), .Q(\ram[9][2] ) );
  DFFHQX1 \ram_reg[9][1]  ( .D(n727), .CK(clk), .Q(\ram[9][1] ) );
  DFFHQX1 \ram_reg[9][0]  ( .D(n726), .CK(clk), .Q(\ram[9][0] ) );
  DFFHQX1 \ram_reg[5][15]  ( .D(n677), .CK(clk), .Q(\ram[5][15] ) );
  DFFHQX1 \ram_reg[5][14]  ( .D(n676), .CK(clk), .Q(\ram[5][14] ) );
  DFFHQX1 \ram_reg[5][13]  ( .D(n675), .CK(clk), .Q(\ram[5][13] ) );
  DFFHQX1 \ram_reg[5][12]  ( .D(n674), .CK(clk), .Q(\ram[5][12] ) );
  DFFHQX1 \ram_reg[5][11]  ( .D(n673), .CK(clk), .Q(\ram[5][11] ) );
  DFFHQX1 \ram_reg[5][10]  ( .D(n672), .CK(clk), .Q(\ram[5][10] ) );
  DFFHQX1 \ram_reg[5][9]  ( .D(n671), .CK(clk), .Q(\ram[5][9] ) );
  DFFHQX1 \ram_reg[5][8]  ( .D(n670), .CK(clk), .Q(\ram[5][8] ) );
  DFFHQX1 \ram_reg[5][7]  ( .D(n669), .CK(clk), .Q(\ram[5][7] ) );
  DFFHQX1 \ram_reg[5][6]  ( .D(n668), .CK(clk), .Q(\ram[5][6] ) );
  DFFHQX1 \ram_reg[5][5]  ( .D(n667), .CK(clk), .Q(\ram[5][5] ) );
  DFFHQX1 \ram_reg[5][4]  ( .D(n666), .CK(clk), .Q(\ram[5][4] ) );
  DFFHQX1 \ram_reg[5][3]  ( .D(n665), .CK(clk), .Q(\ram[5][3] ) );
  DFFHQX1 \ram_reg[5][2]  ( .D(n664), .CK(clk), .Q(\ram[5][2] ) );
  DFFHQX1 \ram_reg[5][1]  ( .D(n663), .CK(clk), .Q(\ram[5][1] ) );
  DFFHQX1 \ram_reg[5][0]  ( .D(n662), .CK(clk), .Q(\ram[5][0] ) );
  DFFHQX1 \ram_reg[1][15]  ( .D(n613), .CK(clk), .Q(\ram[1][15] ) );
  DFFHQX1 \ram_reg[1][14]  ( .D(n612), .CK(clk), .Q(\ram[1][14] ) );
  DFFHQX1 \ram_reg[1][13]  ( .D(n611), .CK(clk), .Q(\ram[1][13] ) );
  DFFHQX1 \ram_reg[1][12]  ( .D(n610), .CK(clk), .Q(\ram[1][12] ) );
  DFFHQX1 \ram_reg[1][11]  ( .D(n609), .CK(clk), .Q(\ram[1][11] ) );
  DFFHQX1 \ram_reg[1][10]  ( .D(n608), .CK(clk), .Q(\ram[1][10] ) );
  DFFHQX1 \ram_reg[1][9]  ( .D(n607), .CK(clk), .Q(\ram[1][9] ) );
  DFFHQX1 \ram_reg[1][8]  ( .D(n606), .CK(clk), .Q(\ram[1][8] ) );
  DFFHQX1 \ram_reg[1][7]  ( .D(n605), .CK(clk), .Q(\ram[1][7] ) );
  DFFHQX1 \ram_reg[1][6]  ( .D(n604), .CK(clk), .Q(\ram[1][6] ) );
  DFFHQX1 \ram_reg[1][5]  ( .D(n603), .CK(clk), .Q(\ram[1][5] ) );
  DFFHQX1 \ram_reg[1][4]  ( .D(n602), .CK(clk), .Q(\ram[1][4] ) );
  DFFHQX1 \ram_reg[1][3]  ( .D(n601), .CK(clk), .Q(\ram[1][3] ) );
  DFFHQX1 \ram_reg[1][2]  ( .D(n600), .CK(clk), .Q(\ram[1][2] ) );
  DFFHQX1 \ram_reg[1][1]  ( .D(n599), .CK(clk), .Q(\ram[1][1] ) );
  DFFHQX1 \ram_reg[1][0]  ( .D(n598), .CK(clk), .Q(\ram[1][0] ) );
  DFFHQX1 \ram_reg[255][15]  ( .D(n4677), .CK(clk), .Q(\ram[255][15] ) );
  DFFHQX1 \ram_reg[255][14]  ( .D(n4676), .CK(clk), .Q(\ram[255][14] ) );
  DFFHQX1 \ram_reg[255][13]  ( .D(n4675), .CK(clk), .Q(\ram[255][13] ) );
  DFFHQX1 \ram_reg[255][12]  ( .D(n4674), .CK(clk), .Q(\ram[255][12] ) );
  DFFHQX1 \ram_reg[255][11]  ( .D(n4673), .CK(clk), .Q(\ram[255][11] ) );
  DFFHQX1 \ram_reg[255][10]  ( .D(n4672), .CK(clk), .Q(\ram[255][10] ) );
  DFFHQX1 \ram_reg[255][9]  ( .D(n4671), .CK(clk), .Q(\ram[255][9] ) );
  DFFHQX1 \ram_reg[255][8]  ( .D(n4670), .CK(clk), .Q(\ram[255][8] ) );
  DFFHQX1 \ram_reg[255][7]  ( .D(n4669), .CK(clk), .Q(\ram[255][7] ) );
  DFFHQX1 \ram_reg[255][6]  ( .D(n4668), .CK(clk), .Q(\ram[255][6] ) );
  DFFHQX1 \ram_reg[255][5]  ( .D(n4667), .CK(clk), .Q(\ram[255][5] ) );
  DFFHQX1 \ram_reg[255][4]  ( .D(n4666), .CK(clk), .Q(\ram[255][4] ) );
  DFFHQX1 \ram_reg[255][3]  ( .D(n4665), .CK(clk), .Q(\ram[255][3] ) );
  DFFHQX1 \ram_reg[255][2]  ( .D(n4664), .CK(clk), .Q(\ram[255][2] ) );
  DFFHQX1 \ram_reg[255][1]  ( .D(n4663), .CK(clk), .Q(\ram[255][1] ) );
  DFFHQX1 \ram_reg[255][0]  ( .D(n4662), .CK(clk), .Q(\ram[255][0] ) );
  DFFHQX1 \ram_reg[251][15]  ( .D(n4613), .CK(clk), .Q(\ram[251][15] ) );
  DFFHQX1 \ram_reg[251][14]  ( .D(n4612), .CK(clk), .Q(\ram[251][14] ) );
  DFFHQX1 \ram_reg[251][13]  ( .D(n4611), .CK(clk), .Q(\ram[251][13] ) );
  DFFHQX1 \ram_reg[251][12]  ( .D(n4610), .CK(clk), .Q(\ram[251][12] ) );
  DFFHQX1 \ram_reg[251][11]  ( .D(n4609), .CK(clk), .Q(\ram[251][11] ) );
  DFFHQX1 \ram_reg[251][10]  ( .D(n4608), .CK(clk), .Q(\ram[251][10] ) );
  DFFHQX1 \ram_reg[251][9]  ( .D(n4607), .CK(clk), .Q(\ram[251][9] ) );
  DFFHQX1 \ram_reg[251][8]  ( .D(n4606), .CK(clk), .Q(\ram[251][8] ) );
  DFFHQX1 \ram_reg[251][7]  ( .D(n4605), .CK(clk), .Q(\ram[251][7] ) );
  DFFHQX1 \ram_reg[251][6]  ( .D(n4604), .CK(clk), .Q(\ram[251][6] ) );
  DFFHQX1 \ram_reg[251][5]  ( .D(n4603), .CK(clk), .Q(\ram[251][5] ) );
  DFFHQX1 \ram_reg[251][4]  ( .D(n4602), .CK(clk), .Q(\ram[251][4] ) );
  DFFHQX1 \ram_reg[251][3]  ( .D(n4601), .CK(clk), .Q(\ram[251][3] ) );
  DFFHQX1 \ram_reg[251][2]  ( .D(n4600), .CK(clk), .Q(\ram[251][2] ) );
  DFFHQX1 \ram_reg[251][1]  ( .D(n4599), .CK(clk), .Q(\ram[251][1] ) );
  DFFHQX1 \ram_reg[251][0]  ( .D(n4598), .CK(clk), .Q(\ram[251][0] ) );
  DFFHQX1 \ram_reg[247][15]  ( .D(n4549), .CK(clk), .Q(\ram[247][15] ) );
  DFFHQX1 \ram_reg[247][14]  ( .D(n4548), .CK(clk), .Q(\ram[247][14] ) );
  DFFHQX1 \ram_reg[247][13]  ( .D(n4547), .CK(clk), .Q(\ram[247][13] ) );
  DFFHQX1 \ram_reg[247][12]  ( .D(n4546), .CK(clk), .Q(\ram[247][12] ) );
  DFFHQX1 \ram_reg[247][11]  ( .D(n4545), .CK(clk), .Q(\ram[247][11] ) );
  DFFHQX1 \ram_reg[247][10]  ( .D(n4544), .CK(clk), .Q(\ram[247][10] ) );
  DFFHQX1 \ram_reg[247][9]  ( .D(n4543), .CK(clk), .Q(\ram[247][9] ) );
  DFFHQX1 \ram_reg[247][8]  ( .D(n4542), .CK(clk), .Q(\ram[247][8] ) );
  DFFHQX1 \ram_reg[247][7]  ( .D(n4541), .CK(clk), .Q(\ram[247][7] ) );
  DFFHQX1 \ram_reg[247][6]  ( .D(n4540), .CK(clk), .Q(\ram[247][6] ) );
  DFFHQX1 \ram_reg[247][5]  ( .D(n4539), .CK(clk), .Q(\ram[247][5] ) );
  DFFHQX1 \ram_reg[247][4]  ( .D(n4538), .CK(clk), .Q(\ram[247][4] ) );
  DFFHQX1 \ram_reg[247][3]  ( .D(n4537), .CK(clk), .Q(\ram[247][3] ) );
  DFFHQX1 \ram_reg[247][2]  ( .D(n4536), .CK(clk), .Q(\ram[247][2] ) );
  DFFHQX1 \ram_reg[247][1]  ( .D(n4535), .CK(clk), .Q(\ram[247][1] ) );
  DFFHQX1 \ram_reg[247][0]  ( .D(n4534), .CK(clk), .Q(\ram[247][0] ) );
  DFFHQX1 \ram_reg[243][15]  ( .D(n4485), .CK(clk), .Q(\ram[243][15] ) );
  DFFHQX1 \ram_reg[243][14]  ( .D(n4484), .CK(clk), .Q(\ram[243][14] ) );
  DFFHQX1 \ram_reg[243][13]  ( .D(n4483), .CK(clk), .Q(\ram[243][13] ) );
  DFFHQX1 \ram_reg[243][12]  ( .D(n4482), .CK(clk), .Q(\ram[243][12] ) );
  DFFHQX1 \ram_reg[243][11]  ( .D(n4481), .CK(clk), .Q(\ram[243][11] ) );
  DFFHQX1 \ram_reg[243][10]  ( .D(n4480), .CK(clk), .Q(\ram[243][10] ) );
  DFFHQX1 \ram_reg[243][9]  ( .D(n4479), .CK(clk), .Q(\ram[243][9] ) );
  DFFHQX1 \ram_reg[243][8]  ( .D(n4478), .CK(clk), .Q(\ram[243][8] ) );
  DFFHQX1 \ram_reg[243][7]  ( .D(n4477), .CK(clk), .Q(\ram[243][7] ) );
  DFFHQX1 \ram_reg[243][6]  ( .D(n4476), .CK(clk), .Q(\ram[243][6] ) );
  DFFHQX1 \ram_reg[243][5]  ( .D(n4475), .CK(clk), .Q(\ram[243][5] ) );
  DFFHQX1 \ram_reg[243][4]  ( .D(n4474), .CK(clk), .Q(\ram[243][4] ) );
  DFFHQX1 \ram_reg[243][3]  ( .D(n4473), .CK(clk), .Q(\ram[243][3] ) );
  DFFHQX1 \ram_reg[243][2]  ( .D(n4472), .CK(clk), .Q(\ram[243][2] ) );
  DFFHQX1 \ram_reg[243][1]  ( .D(n4471), .CK(clk), .Q(\ram[243][1] ) );
  DFFHQX1 \ram_reg[243][0]  ( .D(n4470), .CK(clk), .Q(\ram[243][0] ) );
  DFFHQX1 \ram_reg[239][15]  ( .D(n4421), .CK(clk), .Q(\ram[239][15] ) );
  DFFHQX1 \ram_reg[239][14]  ( .D(n4420), .CK(clk), .Q(\ram[239][14] ) );
  DFFHQX1 \ram_reg[239][13]  ( .D(n4419), .CK(clk), .Q(\ram[239][13] ) );
  DFFHQX1 \ram_reg[239][12]  ( .D(n4418), .CK(clk), .Q(\ram[239][12] ) );
  DFFHQX1 \ram_reg[239][11]  ( .D(n4417), .CK(clk), .Q(\ram[239][11] ) );
  DFFHQX1 \ram_reg[239][10]  ( .D(n4416), .CK(clk), .Q(\ram[239][10] ) );
  DFFHQX1 \ram_reg[239][9]  ( .D(n4415), .CK(clk), .Q(\ram[239][9] ) );
  DFFHQX1 \ram_reg[239][8]  ( .D(n4414), .CK(clk), .Q(\ram[239][8] ) );
  DFFHQX1 \ram_reg[239][7]  ( .D(n4413), .CK(clk), .Q(\ram[239][7] ) );
  DFFHQX1 \ram_reg[239][6]  ( .D(n4412), .CK(clk), .Q(\ram[239][6] ) );
  DFFHQX1 \ram_reg[239][5]  ( .D(n4411), .CK(clk), .Q(\ram[239][5] ) );
  DFFHQX1 \ram_reg[239][4]  ( .D(n4410), .CK(clk), .Q(\ram[239][4] ) );
  DFFHQX1 \ram_reg[239][3]  ( .D(n4409), .CK(clk), .Q(\ram[239][3] ) );
  DFFHQX1 \ram_reg[239][2]  ( .D(n4408), .CK(clk), .Q(\ram[239][2] ) );
  DFFHQX1 \ram_reg[239][1]  ( .D(n4407), .CK(clk), .Q(\ram[239][1] ) );
  DFFHQX1 \ram_reg[239][0]  ( .D(n4406), .CK(clk), .Q(\ram[239][0] ) );
  DFFHQX1 \ram_reg[235][15]  ( .D(n4357), .CK(clk), .Q(\ram[235][15] ) );
  DFFHQX1 \ram_reg[235][14]  ( .D(n4356), .CK(clk), .Q(\ram[235][14] ) );
  DFFHQX1 \ram_reg[235][13]  ( .D(n4355), .CK(clk), .Q(\ram[235][13] ) );
  DFFHQX1 \ram_reg[235][12]  ( .D(n4354), .CK(clk), .Q(\ram[235][12] ) );
  DFFHQX1 \ram_reg[235][11]  ( .D(n4353), .CK(clk), .Q(\ram[235][11] ) );
  DFFHQX1 \ram_reg[235][10]  ( .D(n4352), .CK(clk), .Q(\ram[235][10] ) );
  DFFHQX1 \ram_reg[235][9]  ( .D(n4351), .CK(clk), .Q(\ram[235][9] ) );
  DFFHQX1 \ram_reg[235][8]  ( .D(n4350), .CK(clk), .Q(\ram[235][8] ) );
  DFFHQX1 \ram_reg[235][7]  ( .D(n4349), .CK(clk), .Q(\ram[235][7] ) );
  DFFHQX1 \ram_reg[235][6]  ( .D(n4348), .CK(clk), .Q(\ram[235][6] ) );
  DFFHQX1 \ram_reg[235][5]  ( .D(n4347), .CK(clk), .Q(\ram[235][5] ) );
  DFFHQX1 \ram_reg[235][4]  ( .D(n4346), .CK(clk), .Q(\ram[235][4] ) );
  DFFHQX1 \ram_reg[235][3]  ( .D(n4345), .CK(clk), .Q(\ram[235][3] ) );
  DFFHQX1 \ram_reg[235][2]  ( .D(n4344), .CK(clk), .Q(\ram[235][2] ) );
  DFFHQX1 \ram_reg[235][1]  ( .D(n4343), .CK(clk), .Q(\ram[235][1] ) );
  DFFHQX1 \ram_reg[235][0]  ( .D(n4342), .CK(clk), .Q(\ram[235][0] ) );
  DFFHQX1 \ram_reg[231][15]  ( .D(n4293), .CK(clk), .Q(\ram[231][15] ) );
  DFFHQX1 \ram_reg[231][14]  ( .D(n4292), .CK(clk), .Q(\ram[231][14] ) );
  DFFHQX1 \ram_reg[231][13]  ( .D(n4291), .CK(clk), .Q(\ram[231][13] ) );
  DFFHQX1 \ram_reg[231][12]  ( .D(n4290), .CK(clk), .Q(\ram[231][12] ) );
  DFFHQX1 \ram_reg[231][11]  ( .D(n4289), .CK(clk), .Q(\ram[231][11] ) );
  DFFHQX1 \ram_reg[231][10]  ( .D(n4288), .CK(clk), .Q(\ram[231][10] ) );
  DFFHQX1 \ram_reg[231][9]  ( .D(n4287), .CK(clk), .Q(\ram[231][9] ) );
  DFFHQX1 \ram_reg[231][8]  ( .D(n4286), .CK(clk), .Q(\ram[231][8] ) );
  DFFHQX1 \ram_reg[231][7]  ( .D(n4285), .CK(clk), .Q(\ram[231][7] ) );
  DFFHQX1 \ram_reg[231][6]  ( .D(n4284), .CK(clk), .Q(\ram[231][6] ) );
  DFFHQX1 \ram_reg[231][5]  ( .D(n4283), .CK(clk), .Q(\ram[231][5] ) );
  DFFHQX1 \ram_reg[231][4]  ( .D(n4282), .CK(clk), .Q(\ram[231][4] ) );
  DFFHQX1 \ram_reg[231][3]  ( .D(n4281), .CK(clk), .Q(\ram[231][3] ) );
  DFFHQX1 \ram_reg[231][2]  ( .D(n4280), .CK(clk), .Q(\ram[231][2] ) );
  DFFHQX1 \ram_reg[231][1]  ( .D(n4279), .CK(clk), .Q(\ram[231][1] ) );
  DFFHQX1 \ram_reg[231][0]  ( .D(n4278), .CK(clk), .Q(\ram[231][0] ) );
  DFFHQX1 \ram_reg[227][15]  ( .D(n4229), .CK(clk), .Q(\ram[227][15] ) );
  DFFHQX1 \ram_reg[227][14]  ( .D(n4228), .CK(clk), .Q(\ram[227][14] ) );
  DFFHQX1 \ram_reg[227][13]  ( .D(n4227), .CK(clk), .Q(\ram[227][13] ) );
  DFFHQX1 \ram_reg[227][12]  ( .D(n4226), .CK(clk), .Q(\ram[227][12] ) );
  DFFHQX1 \ram_reg[227][11]  ( .D(n4225), .CK(clk), .Q(\ram[227][11] ) );
  DFFHQX1 \ram_reg[227][10]  ( .D(n4224), .CK(clk), .Q(\ram[227][10] ) );
  DFFHQX1 \ram_reg[227][9]  ( .D(n4223), .CK(clk), .Q(\ram[227][9] ) );
  DFFHQX1 \ram_reg[227][8]  ( .D(n4222), .CK(clk), .Q(\ram[227][8] ) );
  DFFHQX1 \ram_reg[227][7]  ( .D(n4221), .CK(clk), .Q(\ram[227][7] ) );
  DFFHQX1 \ram_reg[227][6]  ( .D(n4220), .CK(clk), .Q(\ram[227][6] ) );
  DFFHQX1 \ram_reg[227][5]  ( .D(n4219), .CK(clk), .Q(\ram[227][5] ) );
  DFFHQX1 \ram_reg[227][4]  ( .D(n4218), .CK(clk), .Q(\ram[227][4] ) );
  DFFHQX1 \ram_reg[227][3]  ( .D(n4217), .CK(clk), .Q(\ram[227][3] ) );
  DFFHQX1 \ram_reg[227][2]  ( .D(n4216), .CK(clk), .Q(\ram[227][2] ) );
  DFFHQX1 \ram_reg[227][1]  ( .D(n4215), .CK(clk), .Q(\ram[227][1] ) );
  DFFHQX1 \ram_reg[227][0]  ( .D(n4214), .CK(clk), .Q(\ram[227][0] ) );
  DFFHQX1 \ram_reg[223][15]  ( .D(n4165), .CK(clk), .Q(\ram[223][15] ) );
  DFFHQX1 \ram_reg[223][14]  ( .D(n4164), .CK(clk), .Q(\ram[223][14] ) );
  DFFHQX1 \ram_reg[223][13]  ( .D(n4163), .CK(clk), .Q(\ram[223][13] ) );
  DFFHQX1 \ram_reg[223][12]  ( .D(n4162), .CK(clk), .Q(\ram[223][12] ) );
  DFFHQX1 \ram_reg[223][11]  ( .D(n4161), .CK(clk), .Q(\ram[223][11] ) );
  DFFHQX1 \ram_reg[223][10]  ( .D(n4160), .CK(clk), .Q(\ram[223][10] ) );
  DFFHQX1 \ram_reg[223][9]  ( .D(n4159), .CK(clk), .Q(\ram[223][9] ) );
  DFFHQX1 \ram_reg[223][8]  ( .D(n4158), .CK(clk), .Q(\ram[223][8] ) );
  DFFHQX1 \ram_reg[223][7]  ( .D(n4157), .CK(clk), .Q(\ram[223][7] ) );
  DFFHQX1 \ram_reg[223][6]  ( .D(n4156), .CK(clk), .Q(\ram[223][6] ) );
  DFFHQX1 \ram_reg[223][5]  ( .D(n4155), .CK(clk), .Q(\ram[223][5] ) );
  DFFHQX1 \ram_reg[223][4]  ( .D(n4154), .CK(clk), .Q(\ram[223][4] ) );
  DFFHQX1 \ram_reg[223][3]  ( .D(n4153), .CK(clk), .Q(\ram[223][3] ) );
  DFFHQX1 \ram_reg[223][2]  ( .D(n4152), .CK(clk), .Q(\ram[223][2] ) );
  DFFHQX1 \ram_reg[223][1]  ( .D(n4151), .CK(clk), .Q(\ram[223][1] ) );
  DFFHQX1 \ram_reg[223][0]  ( .D(n4150), .CK(clk), .Q(\ram[223][0] ) );
  DFFHQX1 \ram_reg[219][15]  ( .D(n4101), .CK(clk), .Q(\ram[219][15] ) );
  DFFHQX1 \ram_reg[219][14]  ( .D(n4100), .CK(clk), .Q(\ram[219][14] ) );
  DFFHQX1 \ram_reg[219][13]  ( .D(n4099), .CK(clk), .Q(\ram[219][13] ) );
  DFFHQX1 \ram_reg[219][12]  ( .D(n4098), .CK(clk), .Q(\ram[219][12] ) );
  DFFHQX1 \ram_reg[219][11]  ( .D(n4097), .CK(clk), .Q(\ram[219][11] ) );
  DFFHQX1 \ram_reg[219][10]  ( .D(n4096), .CK(clk), .Q(\ram[219][10] ) );
  DFFHQX1 \ram_reg[219][9]  ( .D(n4095), .CK(clk), .Q(\ram[219][9] ) );
  DFFHQX1 \ram_reg[219][8]  ( .D(n4094), .CK(clk), .Q(\ram[219][8] ) );
  DFFHQX1 \ram_reg[219][7]  ( .D(n4093), .CK(clk), .Q(\ram[219][7] ) );
  DFFHQX1 \ram_reg[219][6]  ( .D(n4092), .CK(clk), .Q(\ram[219][6] ) );
  DFFHQX1 \ram_reg[219][5]  ( .D(n4091), .CK(clk), .Q(\ram[219][5] ) );
  DFFHQX1 \ram_reg[219][4]  ( .D(n4090), .CK(clk), .Q(\ram[219][4] ) );
  DFFHQX1 \ram_reg[219][3]  ( .D(n4089), .CK(clk), .Q(\ram[219][3] ) );
  DFFHQX1 \ram_reg[219][2]  ( .D(n4088), .CK(clk), .Q(\ram[219][2] ) );
  DFFHQX1 \ram_reg[219][1]  ( .D(n4087), .CK(clk), .Q(\ram[219][1] ) );
  DFFHQX1 \ram_reg[219][0]  ( .D(n4086), .CK(clk), .Q(\ram[219][0] ) );
  DFFHQX1 \ram_reg[215][15]  ( .D(n4037), .CK(clk), .Q(\ram[215][15] ) );
  DFFHQX1 \ram_reg[215][14]  ( .D(n4036), .CK(clk), .Q(\ram[215][14] ) );
  DFFHQX1 \ram_reg[215][13]  ( .D(n4035), .CK(clk), .Q(\ram[215][13] ) );
  DFFHQX1 \ram_reg[215][12]  ( .D(n4034), .CK(clk), .Q(\ram[215][12] ) );
  DFFHQX1 \ram_reg[215][11]  ( .D(n4033), .CK(clk), .Q(\ram[215][11] ) );
  DFFHQX1 \ram_reg[215][10]  ( .D(n4032), .CK(clk), .Q(\ram[215][10] ) );
  DFFHQX1 \ram_reg[215][9]  ( .D(n4031), .CK(clk), .Q(\ram[215][9] ) );
  DFFHQX1 \ram_reg[215][8]  ( .D(n4030), .CK(clk), .Q(\ram[215][8] ) );
  DFFHQX1 \ram_reg[215][7]  ( .D(n4029), .CK(clk), .Q(\ram[215][7] ) );
  DFFHQX1 \ram_reg[215][6]  ( .D(n4028), .CK(clk), .Q(\ram[215][6] ) );
  DFFHQX1 \ram_reg[215][5]  ( .D(n4027), .CK(clk), .Q(\ram[215][5] ) );
  DFFHQX1 \ram_reg[215][4]  ( .D(n4026), .CK(clk), .Q(\ram[215][4] ) );
  DFFHQX1 \ram_reg[215][3]  ( .D(n4025), .CK(clk), .Q(\ram[215][3] ) );
  DFFHQX1 \ram_reg[215][2]  ( .D(n4024), .CK(clk), .Q(\ram[215][2] ) );
  DFFHQX1 \ram_reg[215][1]  ( .D(n4023), .CK(clk), .Q(\ram[215][1] ) );
  DFFHQX1 \ram_reg[215][0]  ( .D(n4022), .CK(clk), .Q(\ram[215][0] ) );
  DFFHQX1 \ram_reg[211][15]  ( .D(n3973), .CK(clk), .Q(\ram[211][15] ) );
  DFFHQX1 \ram_reg[211][14]  ( .D(n3972), .CK(clk), .Q(\ram[211][14] ) );
  DFFHQX1 \ram_reg[211][13]  ( .D(n3971), .CK(clk), .Q(\ram[211][13] ) );
  DFFHQX1 \ram_reg[211][12]  ( .D(n3970), .CK(clk), .Q(\ram[211][12] ) );
  DFFHQX1 \ram_reg[211][11]  ( .D(n3969), .CK(clk), .Q(\ram[211][11] ) );
  DFFHQX1 \ram_reg[211][10]  ( .D(n3968), .CK(clk), .Q(\ram[211][10] ) );
  DFFHQX1 \ram_reg[211][9]  ( .D(n3967), .CK(clk), .Q(\ram[211][9] ) );
  DFFHQX1 \ram_reg[211][8]  ( .D(n3966), .CK(clk), .Q(\ram[211][8] ) );
  DFFHQX1 \ram_reg[211][7]  ( .D(n3965), .CK(clk), .Q(\ram[211][7] ) );
  DFFHQX1 \ram_reg[211][6]  ( .D(n3964), .CK(clk), .Q(\ram[211][6] ) );
  DFFHQX1 \ram_reg[211][5]  ( .D(n3963), .CK(clk), .Q(\ram[211][5] ) );
  DFFHQX1 \ram_reg[211][4]  ( .D(n3962), .CK(clk), .Q(\ram[211][4] ) );
  DFFHQX1 \ram_reg[211][3]  ( .D(n3961), .CK(clk), .Q(\ram[211][3] ) );
  DFFHQX1 \ram_reg[211][2]  ( .D(n3960), .CK(clk), .Q(\ram[211][2] ) );
  DFFHQX1 \ram_reg[211][1]  ( .D(n3959), .CK(clk), .Q(\ram[211][1] ) );
  DFFHQX1 \ram_reg[211][0]  ( .D(n3958), .CK(clk), .Q(\ram[211][0] ) );
  DFFHQX1 \ram_reg[207][15]  ( .D(n3909), .CK(clk), .Q(\ram[207][15] ) );
  DFFHQX1 \ram_reg[207][14]  ( .D(n3908), .CK(clk), .Q(\ram[207][14] ) );
  DFFHQX1 \ram_reg[207][13]  ( .D(n3907), .CK(clk), .Q(\ram[207][13] ) );
  DFFHQX1 \ram_reg[207][12]  ( .D(n3906), .CK(clk), .Q(\ram[207][12] ) );
  DFFHQX1 \ram_reg[207][11]  ( .D(n3905), .CK(clk), .Q(\ram[207][11] ) );
  DFFHQX1 \ram_reg[207][10]  ( .D(n3904), .CK(clk), .Q(\ram[207][10] ) );
  DFFHQX1 \ram_reg[207][9]  ( .D(n3903), .CK(clk), .Q(\ram[207][9] ) );
  DFFHQX1 \ram_reg[207][8]  ( .D(n3902), .CK(clk), .Q(\ram[207][8] ) );
  DFFHQX1 \ram_reg[207][7]  ( .D(n3901), .CK(clk), .Q(\ram[207][7] ) );
  DFFHQX1 \ram_reg[207][6]  ( .D(n3900), .CK(clk), .Q(\ram[207][6] ) );
  DFFHQX1 \ram_reg[207][5]  ( .D(n3899), .CK(clk), .Q(\ram[207][5] ) );
  DFFHQX1 \ram_reg[207][4]  ( .D(n3898), .CK(clk), .Q(\ram[207][4] ) );
  DFFHQX1 \ram_reg[207][3]  ( .D(n3897), .CK(clk), .Q(\ram[207][3] ) );
  DFFHQX1 \ram_reg[207][2]  ( .D(n3896), .CK(clk), .Q(\ram[207][2] ) );
  DFFHQX1 \ram_reg[207][1]  ( .D(n3895), .CK(clk), .Q(\ram[207][1] ) );
  DFFHQX1 \ram_reg[207][0]  ( .D(n3894), .CK(clk), .Q(\ram[207][0] ) );
  DFFHQX1 \ram_reg[203][15]  ( .D(n3845), .CK(clk), .Q(\ram[203][15] ) );
  DFFHQX1 \ram_reg[203][14]  ( .D(n3844), .CK(clk), .Q(\ram[203][14] ) );
  DFFHQX1 \ram_reg[203][13]  ( .D(n3843), .CK(clk), .Q(\ram[203][13] ) );
  DFFHQX1 \ram_reg[203][12]  ( .D(n3842), .CK(clk), .Q(\ram[203][12] ) );
  DFFHQX1 \ram_reg[203][11]  ( .D(n3841), .CK(clk), .Q(\ram[203][11] ) );
  DFFHQX1 \ram_reg[203][10]  ( .D(n3840), .CK(clk), .Q(\ram[203][10] ) );
  DFFHQX1 \ram_reg[203][9]  ( .D(n3839), .CK(clk), .Q(\ram[203][9] ) );
  DFFHQX1 \ram_reg[203][8]  ( .D(n3838), .CK(clk), .Q(\ram[203][8] ) );
  DFFHQX1 \ram_reg[203][7]  ( .D(n3837), .CK(clk), .Q(\ram[203][7] ) );
  DFFHQX1 \ram_reg[203][6]  ( .D(n3836), .CK(clk), .Q(\ram[203][6] ) );
  DFFHQX1 \ram_reg[203][5]  ( .D(n3835), .CK(clk), .Q(\ram[203][5] ) );
  DFFHQX1 \ram_reg[203][4]  ( .D(n3834), .CK(clk), .Q(\ram[203][4] ) );
  DFFHQX1 \ram_reg[203][3]  ( .D(n3833), .CK(clk), .Q(\ram[203][3] ) );
  DFFHQX1 \ram_reg[203][2]  ( .D(n3832), .CK(clk), .Q(\ram[203][2] ) );
  DFFHQX1 \ram_reg[203][1]  ( .D(n3831), .CK(clk), .Q(\ram[203][1] ) );
  DFFHQX1 \ram_reg[203][0]  ( .D(n3830), .CK(clk), .Q(\ram[203][0] ) );
  DFFHQX1 \ram_reg[199][15]  ( .D(n3781), .CK(clk), .Q(\ram[199][15] ) );
  DFFHQX1 \ram_reg[199][14]  ( .D(n3780), .CK(clk), .Q(\ram[199][14] ) );
  DFFHQX1 \ram_reg[199][13]  ( .D(n3779), .CK(clk), .Q(\ram[199][13] ) );
  DFFHQX1 \ram_reg[199][12]  ( .D(n3778), .CK(clk), .Q(\ram[199][12] ) );
  DFFHQX1 \ram_reg[199][11]  ( .D(n3777), .CK(clk), .Q(\ram[199][11] ) );
  DFFHQX1 \ram_reg[199][10]  ( .D(n3776), .CK(clk), .Q(\ram[199][10] ) );
  DFFHQX1 \ram_reg[199][9]  ( .D(n3775), .CK(clk), .Q(\ram[199][9] ) );
  DFFHQX1 \ram_reg[199][8]  ( .D(n3774), .CK(clk), .Q(\ram[199][8] ) );
  DFFHQX1 \ram_reg[199][7]  ( .D(n3773), .CK(clk), .Q(\ram[199][7] ) );
  DFFHQX1 \ram_reg[199][6]  ( .D(n3772), .CK(clk), .Q(\ram[199][6] ) );
  DFFHQX1 \ram_reg[199][5]  ( .D(n3771), .CK(clk), .Q(\ram[199][5] ) );
  DFFHQX1 \ram_reg[199][4]  ( .D(n3770), .CK(clk), .Q(\ram[199][4] ) );
  DFFHQX1 \ram_reg[199][3]  ( .D(n3769), .CK(clk), .Q(\ram[199][3] ) );
  DFFHQX1 \ram_reg[199][2]  ( .D(n3768), .CK(clk), .Q(\ram[199][2] ) );
  DFFHQX1 \ram_reg[199][1]  ( .D(n3767), .CK(clk), .Q(\ram[199][1] ) );
  DFFHQX1 \ram_reg[199][0]  ( .D(n3766), .CK(clk), .Q(\ram[199][0] ) );
  DFFHQX1 \ram_reg[195][15]  ( .D(n3717), .CK(clk), .Q(\ram[195][15] ) );
  DFFHQX1 \ram_reg[195][14]  ( .D(n3716), .CK(clk), .Q(\ram[195][14] ) );
  DFFHQX1 \ram_reg[195][13]  ( .D(n3715), .CK(clk), .Q(\ram[195][13] ) );
  DFFHQX1 \ram_reg[195][12]  ( .D(n3714), .CK(clk), .Q(\ram[195][12] ) );
  DFFHQX1 \ram_reg[195][11]  ( .D(n3713), .CK(clk), .Q(\ram[195][11] ) );
  DFFHQX1 \ram_reg[195][10]  ( .D(n3712), .CK(clk), .Q(\ram[195][10] ) );
  DFFHQX1 \ram_reg[195][9]  ( .D(n3711), .CK(clk), .Q(\ram[195][9] ) );
  DFFHQX1 \ram_reg[195][8]  ( .D(n3710), .CK(clk), .Q(\ram[195][8] ) );
  DFFHQX1 \ram_reg[195][7]  ( .D(n3709), .CK(clk), .Q(\ram[195][7] ) );
  DFFHQX1 \ram_reg[195][6]  ( .D(n3708), .CK(clk), .Q(\ram[195][6] ) );
  DFFHQX1 \ram_reg[195][5]  ( .D(n3707), .CK(clk), .Q(\ram[195][5] ) );
  DFFHQX1 \ram_reg[195][4]  ( .D(n3706), .CK(clk), .Q(\ram[195][4] ) );
  DFFHQX1 \ram_reg[195][3]  ( .D(n3705), .CK(clk), .Q(\ram[195][3] ) );
  DFFHQX1 \ram_reg[195][2]  ( .D(n3704), .CK(clk), .Q(\ram[195][2] ) );
  DFFHQX1 \ram_reg[195][1]  ( .D(n3703), .CK(clk), .Q(\ram[195][1] ) );
  DFFHQX1 \ram_reg[195][0]  ( .D(n3702), .CK(clk), .Q(\ram[195][0] ) );
  DFFHQX1 \ram_reg[191][15]  ( .D(n3653), .CK(clk), .Q(\ram[191][15] ) );
  DFFHQX1 \ram_reg[191][14]  ( .D(n3652), .CK(clk), .Q(\ram[191][14] ) );
  DFFHQX1 \ram_reg[191][13]  ( .D(n3651), .CK(clk), .Q(\ram[191][13] ) );
  DFFHQX1 \ram_reg[191][12]  ( .D(n3650), .CK(clk), .Q(\ram[191][12] ) );
  DFFHQX1 \ram_reg[191][11]  ( .D(n3649), .CK(clk), .Q(\ram[191][11] ) );
  DFFHQX1 \ram_reg[191][10]  ( .D(n3648), .CK(clk), .Q(\ram[191][10] ) );
  DFFHQX1 \ram_reg[191][9]  ( .D(n3647), .CK(clk), .Q(\ram[191][9] ) );
  DFFHQX1 \ram_reg[191][8]  ( .D(n3646), .CK(clk), .Q(\ram[191][8] ) );
  DFFHQX1 \ram_reg[191][7]  ( .D(n3645), .CK(clk), .Q(\ram[191][7] ) );
  DFFHQX1 \ram_reg[191][6]  ( .D(n3644), .CK(clk), .Q(\ram[191][6] ) );
  DFFHQX1 \ram_reg[191][5]  ( .D(n3643), .CK(clk), .Q(\ram[191][5] ) );
  DFFHQX1 \ram_reg[191][4]  ( .D(n3642), .CK(clk), .Q(\ram[191][4] ) );
  DFFHQX1 \ram_reg[191][3]  ( .D(n3641), .CK(clk), .Q(\ram[191][3] ) );
  DFFHQX1 \ram_reg[191][2]  ( .D(n3640), .CK(clk), .Q(\ram[191][2] ) );
  DFFHQX1 \ram_reg[191][1]  ( .D(n3639), .CK(clk), .Q(\ram[191][1] ) );
  DFFHQX1 \ram_reg[191][0]  ( .D(n3638), .CK(clk), .Q(\ram[191][0] ) );
  DFFHQX1 \ram_reg[187][15]  ( .D(n3589), .CK(clk), .Q(\ram[187][15] ) );
  DFFHQX1 \ram_reg[187][14]  ( .D(n3588), .CK(clk), .Q(\ram[187][14] ) );
  DFFHQX1 \ram_reg[187][13]  ( .D(n3587), .CK(clk), .Q(\ram[187][13] ) );
  DFFHQX1 \ram_reg[187][12]  ( .D(n3586), .CK(clk), .Q(\ram[187][12] ) );
  DFFHQX1 \ram_reg[187][11]  ( .D(n3585), .CK(clk), .Q(\ram[187][11] ) );
  DFFHQX1 \ram_reg[187][10]  ( .D(n3584), .CK(clk), .Q(\ram[187][10] ) );
  DFFHQX1 \ram_reg[187][9]  ( .D(n3583), .CK(clk), .Q(\ram[187][9] ) );
  DFFHQX1 \ram_reg[187][8]  ( .D(n3582), .CK(clk), .Q(\ram[187][8] ) );
  DFFHQX1 \ram_reg[187][7]  ( .D(n3581), .CK(clk), .Q(\ram[187][7] ) );
  DFFHQX1 \ram_reg[187][6]  ( .D(n3580), .CK(clk), .Q(\ram[187][6] ) );
  DFFHQX1 \ram_reg[187][5]  ( .D(n3579), .CK(clk), .Q(\ram[187][5] ) );
  DFFHQX1 \ram_reg[187][4]  ( .D(n3578), .CK(clk), .Q(\ram[187][4] ) );
  DFFHQX1 \ram_reg[187][3]  ( .D(n3577), .CK(clk), .Q(\ram[187][3] ) );
  DFFHQX1 \ram_reg[187][2]  ( .D(n3576), .CK(clk), .Q(\ram[187][2] ) );
  DFFHQX1 \ram_reg[187][1]  ( .D(n3575), .CK(clk), .Q(\ram[187][1] ) );
  DFFHQX1 \ram_reg[187][0]  ( .D(n3574), .CK(clk), .Q(\ram[187][0] ) );
  DFFHQX1 \ram_reg[183][15]  ( .D(n3525), .CK(clk), .Q(\ram[183][15] ) );
  DFFHQX1 \ram_reg[183][14]  ( .D(n3524), .CK(clk), .Q(\ram[183][14] ) );
  DFFHQX1 \ram_reg[183][13]  ( .D(n3523), .CK(clk), .Q(\ram[183][13] ) );
  DFFHQX1 \ram_reg[183][12]  ( .D(n3522), .CK(clk), .Q(\ram[183][12] ) );
  DFFHQX1 \ram_reg[183][11]  ( .D(n3521), .CK(clk), .Q(\ram[183][11] ) );
  DFFHQX1 \ram_reg[183][10]  ( .D(n3520), .CK(clk), .Q(\ram[183][10] ) );
  DFFHQX1 \ram_reg[183][9]  ( .D(n3519), .CK(clk), .Q(\ram[183][9] ) );
  DFFHQX1 \ram_reg[183][8]  ( .D(n3518), .CK(clk), .Q(\ram[183][8] ) );
  DFFHQX1 \ram_reg[183][7]  ( .D(n3517), .CK(clk), .Q(\ram[183][7] ) );
  DFFHQX1 \ram_reg[183][6]  ( .D(n3516), .CK(clk), .Q(\ram[183][6] ) );
  DFFHQX1 \ram_reg[183][5]  ( .D(n3515), .CK(clk), .Q(\ram[183][5] ) );
  DFFHQX1 \ram_reg[183][4]  ( .D(n3514), .CK(clk), .Q(\ram[183][4] ) );
  DFFHQX1 \ram_reg[183][3]  ( .D(n3513), .CK(clk), .Q(\ram[183][3] ) );
  DFFHQX1 \ram_reg[183][2]  ( .D(n3512), .CK(clk), .Q(\ram[183][2] ) );
  DFFHQX1 \ram_reg[183][1]  ( .D(n3511), .CK(clk), .Q(\ram[183][1] ) );
  DFFHQX1 \ram_reg[183][0]  ( .D(n3510), .CK(clk), .Q(\ram[183][0] ) );
  DFFHQX1 \ram_reg[179][15]  ( .D(n3461), .CK(clk), .Q(\ram[179][15] ) );
  DFFHQX1 \ram_reg[179][14]  ( .D(n3460), .CK(clk), .Q(\ram[179][14] ) );
  DFFHQX1 \ram_reg[179][13]  ( .D(n3459), .CK(clk), .Q(\ram[179][13] ) );
  DFFHQX1 \ram_reg[179][12]  ( .D(n3458), .CK(clk), .Q(\ram[179][12] ) );
  DFFHQX1 \ram_reg[179][11]  ( .D(n3457), .CK(clk), .Q(\ram[179][11] ) );
  DFFHQX1 \ram_reg[179][10]  ( .D(n3456), .CK(clk), .Q(\ram[179][10] ) );
  DFFHQX1 \ram_reg[179][9]  ( .D(n3455), .CK(clk), .Q(\ram[179][9] ) );
  DFFHQX1 \ram_reg[179][8]  ( .D(n3454), .CK(clk), .Q(\ram[179][8] ) );
  DFFHQX1 \ram_reg[179][7]  ( .D(n3453), .CK(clk), .Q(\ram[179][7] ) );
  DFFHQX1 \ram_reg[179][6]  ( .D(n3452), .CK(clk), .Q(\ram[179][6] ) );
  DFFHQX1 \ram_reg[179][5]  ( .D(n3451), .CK(clk), .Q(\ram[179][5] ) );
  DFFHQX1 \ram_reg[179][4]  ( .D(n3450), .CK(clk), .Q(\ram[179][4] ) );
  DFFHQX1 \ram_reg[179][3]  ( .D(n3449), .CK(clk), .Q(\ram[179][3] ) );
  DFFHQX1 \ram_reg[179][2]  ( .D(n3448), .CK(clk), .Q(\ram[179][2] ) );
  DFFHQX1 \ram_reg[179][1]  ( .D(n3447), .CK(clk), .Q(\ram[179][1] ) );
  DFFHQX1 \ram_reg[179][0]  ( .D(n3446), .CK(clk), .Q(\ram[179][0] ) );
  DFFHQX1 \ram_reg[175][15]  ( .D(n3397), .CK(clk), .Q(\ram[175][15] ) );
  DFFHQX1 \ram_reg[175][14]  ( .D(n3396), .CK(clk), .Q(\ram[175][14] ) );
  DFFHQX1 \ram_reg[175][13]  ( .D(n3395), .CK(clk), .Q(\ram[175][13] ) );
  DFFHQX1 \ram_reg[175][12]  ( .D(n3394), .CK(clk), .Q(\ram[175][12] ) );
  DFFHQX1 \ram_reg[175][11]  ( .D(n3393), .CK(clk), .Q(\ram[175][11] ) );
  DFFHQX1 \ram_reg[175][10]  ( .D(n3392), .CK(clk), .Q(\ram[175][10] ) );
  DFFHQX1 \ram_reg[175][9]  ( .D(n3391), .CK(clk), .Q(\ram[175][9] ) );
  DFFHQX1 \ram_reg[175][8]  ( .D(n3390), .CK(clk), .Q(\ram[175][8] ) );
  DFFHQX1 \ram_reg[175][7]  ( .D(n3389), .CK(clk), .Q(\ram[175][7] ) );
  DFFHQX1 \ram_reg[175][6]  ( .D(n3388), .CK(clk), .Q(\ram[175][6] ) );
  DFFHQX1 \ram_reg[175][5]  ( .D(n3387), .CK(clk), .Q(\ram[175][5] ) );
  DFFHQX1 \ram_reg[175][4]  ( .D(n3386), .CK(clk), .Q(\ram[175][4] ) );
  DFFHQX1 \ram_reg[175][3]  ( .D(n3385), .CK(clk), .Q(\ram[175][3] ) );
  DFFHQX1 \ram_reg[175][2]  ( .D(n3384), .CK(clk), .Q(\ram[175][2] ) );
  DFFHQX1 \ram_reg[175][1]  ( .D(n3383), .CK(clk), .Q(\ram[175][1] ) );
  DFFHQX1 \ram_reg[175][0]  ( .D(n3382), .CK(clk), .Q(\ram[175][0] ) );
  DFFHQX1 \ram_reg[171][15]  ( .D(n3333), .CK(clk), .Q(\ram[171][15] ) );
  DFFHQX1 \ram_reg[171][14]  ( .D(n3332), .CK(clk), .Q(\ram[171][14] ) );
  DFFHQX1 \ram_reg[171][13]  ( .D(n3331), .CK(clk), .Q(\ram[171][13] ) );
  DFFHQX1 \ram_reg[171][12]  ( .D(n3330), .CK(clk), .Q(\ram[171][12] ) );
  DFFHQX1 \ram_reg[171][11]  ( .D(n3329), .CK(clk), .Q(\ram[171][11] ) );
  DFFHQX1 \ram_reg[171][10]  ( .D(n3328), .CK(clk), .Q(\ram[171][10] ) );
  DFFHQX1 \ram_reg[171][9]  ( .D(n3327), .CK(clk), .Q(\ram[171][9] ) );
  DFFHQX1 \ram_reg[171][8]  ( .D(n3326), .CK(clk), .Q(\ram[171][8] ) );
  DFFHQX1 \ram_reg[171][7]  ( .D(n3325), .CK(clk), .Q(\ram[171][7] ) );
  DFFHQX1 \ram_reg[171][6]  ( .D(n3324), .CK(clk), .Q(\ram[171][6] ) );
  DFFHQX1 \ram_reg[171][5]  ( .D(n3323), .CK(clk), .Q(\ram[171][5] ) );
  DFFHQX1 \ram_reg[171][4]  ( .D(n3322), .CK(clk), .Q(\ram[171][4] ) );
  DFFHQX1 \ram_reg[171][3]  ( .D(n3321), .CK(clk), .Q(\ram[171][3] ) );
  DFFHQX1 \ram_reg[171][2]  ( .D(n3320), .CK(clk), .Q(\ram[171][2] ) );
  DFFHQX1 \ram_reg[171][1]  ( .D(n3319), .CK(clk), .Q(\ram[171][1] ) );
  DFFHQX1 \ram_reg[171][0]  ( .D(n3318), .CK(clk), .Q(\ram[171][0] ) );
  DFFHQX1 \ram_reg[167][15]  ( .D(n3269), .CK(clk), .Q(\ram[167][15] ) );
  DFFHQX1 \ram_reg[167][14]  ( .D(n3268), .CK(clk), .Q(\ram[167][14] ) );
  DFFHQX1 \ram_reg[167][13]  ( .D(n3267), .CK(clk), .Q(\ram[167][13] ) );
  DFFHQX1 \ram_reg[167][12]  ( .D(n3266), .CK(clk), .Q(\ram[167][12] ) );
  DFFHQX1 \ram_reg[167][11]  ( .D(n3265), .CK(clk), .Q(\ram[167][11] ) );
  DFFHQX1 \ram_reg[167][10]  ( .D(n3264), .CK(clk), .Q(\ram[167][10] ) );
  DFFHQX1 \ram_reg[167][9]  ( .D(n3263), .CK(clk), .Q(\ram[167][9] ) );
  DFFHQX1 \ram_reg[167][8]  ( .D(n3262), .CK(clk), .Q(\ram[167][8] ) );
  DFFHQX1 \ram_reg[167][7]  ( .D(n3261), .CK(clk), .Q(\ram[167][7] ) );
  DFFHQX1 \ram_reg[167][6]  ( .D(n3260), .CK(clk), .Q(\ram[167][6] ) );
  DFFHQX1 \ram_reg[167][5]  ( .D(n3259), .CK(clk), .Q(\ram[167][5] ) );
  DFFHQX1 \ram_reg[167][4]  ( .D(n3258), .CK(clk), .Q(\ram[167][4] ) );
  DFFHQX1 \ram_reg[167][3]  ( .D(n3257), .CK(clk), .Q(\ram[167][3] ) );
  DFFHQX1 \ram_reg[167][2]  ( .D(n3256), .CK(clk), .Q(\ram[167][2] ) );
  DFFHQX1 \ram_reg[167][1]  ( .D(n3255), .CK(clk), .Q(\ram[167][1] ) );
  DFFHQX1 \ram_reg[167][0]  ( .D(n3254), .CK(clk), .Q(\ram[167][0] ) );
  DFFHQX1 \ram_reg[163][15]  ( .D(n3205), .CK(clk), .Q(\ram[163][15] ) );
  DFFHQX1 \ram_reg[163][14]  ( .D(n3204), .CK(clk), .Q(\ram[163][14] ) );
  DFFHQX1 \ram_reg[163][13]  ( .D(n3203), .CK(clk), .Q(\ram[163][13] ) );
  DFFHQX1 \ram_reg[163][12]  ( .D(n3202), .CK(clk), .Q(\ram[163][12] ) );
  DFFHQX1 \ram_reg[163][11]  ( .D(n3201), .CK(clk), .Q(\ram[163][11] ) );
  DFFHQX1 \ram_reg[163][10]  ( .D(n3200), .CK(clk), .Q(\ram[163][10] ) );
  DFFHQX1 \ram_reg[163][9]  ( .D(n3199), .CK(clk), .Q(\ram[163][9] ) );
  DFFHQX1 \ram_reg[163][8]  ( .D(n3198), .CK(clk), .Q(\ram[163][8] ) );
  DFFHQX1 \ram_reg[163][7]  ( .D(n3197), .CK(clk), .Q(\ram[163][7] ) );
  DFFHQX1 \ram_reg[163][6]  ( .D(n3196), .CK(clk), .Q(\ram[163][6] ) );
  DFFHQX1 \ram_reg[163][5]  ( .D(n3195), .CK(clk), .Q(\ram[163][5] ) );
  DFFHQX1 \ram_reg[163][4]  ( .D(n3194), .CK(clk), .Q(\ram[163][4] ) );
  DFFHQX1 \ram_reg[163][3]  ( .D(n3193), .CK(clk), .Q(\ram[163][3] ) );
  DFFHQX1 \ram_reg[163][2]  ( .D(n3192), .CK(clk), .Q(\ram[163][2] ) );
  DFFHQX1 \ram_reg[163][1]  ( .D(n3191), .CK(clk), .Q(\ram[163][1] ) );
  DFFHQX1 \ram_reg[163][0]  ( .D(n3190), .CK(clk), .Q(\ram[163][0] ) );
  DFFHQX1 \ram_reg[159][15]  ( .D(n3141), .CK(clk), .Q(\ram[159][15] ) );
  DFFHQX1 \ram_reg[159][14]  ( .D(n3140), .CK(clk), .Q(\ram[159][14] ) );
  DFFHQX1 \ram_reg[159][13]  ( .D(n3139), .CK(clk), .Q(\ram[159][13] ) );
  DFFHQX1 \ram_reg[159][12]  ( .D(n3138), .CK(clk), .Q(\ram[159][12] ) );
  DFFHQX1 \ram_reg[159][11]  ( .D(n3137), .CK(clk), .Q(\ram[159][11] ) );
  DFFHQX1 \ram_reg[159][10]  ( .D(n3136), .CK(clk), .Q(\ram[159][10] ) );
  DFFHQX1 \ram_reg[159][9]  ( .D(n3135), .CK(clk), .Q(\ram[159][9] ) );
  DFFHQX1 \ram_reg[159][8]  ( .D(n3134), .CK(clk), .Q(\ram[159][8] ) );
  DFFHQX1 \ram_reg[159][7]  ( .D(n3133), .CK(clk), .Q(\ram[159][7] ) );
  DFFHQX1 \ram_reg[159][6]  ( .D(n3132), .CK(clk), .Q(\ram[159][6] ) );
  DFFHQX1 \ram_reg[159][5]  ( .D(n3131), .CK(clk), .Q(\ram[159][5] ) );
  DFFHQX1 \ram_reg[159][4]  ( .D(n3130), .CK(clk), .Q(\ram[159][4] ) );
  DFFHQX1 \ram_reg[159][3]  ( .D(n3129), .CK(clk), .Q(\ram[159][3] ) );
  DFFHQX1 \ram_reg[159][2]  ( .D(n3128), .CK(clk), .Q(\ram[159][2] ) );
  DFFHQX1 \ram_reg[159][1]  ( .D(n3127), .CK(clk), .Q(\ram[159][1] ) );
  DFFHQX1 \ram_reg[159][0]  ( .D(n3126), .CK(clk), .Q(\ram[159][0] ) );
  DFFHQX1 \ram_reg[155][15]  ( .D(n3077), .CK(clk), .Q(\ram[155][15] ) );
  DFFHQX1 \ram_reg[155][14]  ( .D(n3076), .CK(clk), .Q(\ram[155][14] ) );
  DFFHQX1 \ram_reg[155][13]  ( .D(n3075), .CK(clk), .Q(\ram[155][13] ) );
  DFFHQX1 \ram_reg[155][12]  ( .D(n3074), .CK(clk), .Q(\ram[155][12] ) );
  DFFHQX1 \ram_reg[155][11]  ( .D(n3073), .CK(clk), .Q(\ram[155][11] ) );
  DFFHQX1 \ram_reg[155][10]  ( .D(n3072), .CK(clk), .Q(\ram[155][10] ) );
  DFFHQX1 \ram_reg[155][9]  ( .D(n3071), .CK(clk), .Q(\ram[155][9] ) );
  DFFHQX1 \ram_reg[155][8]  ( .D(n3070), .CK(clk), .Q(\ram[155][8] ) );
  DFFHQX1 \ram_reg[155][7]  ( .D(n3069), .CK(clk), .Q(\ram[155][7] ) );
  DFFHQX1 \ram_reg[155][6]  ( .D(n3068), .CK(clk), .Q(\ram[155][6] ) );
  DFFHQX1 \ram_reg[155][5]  ( .D(n3067), .CK(clk), .Q(\ram[155][5] ) );
  DFFHQX1 \ram_reg[155][4]  ( .D(n3066), .CK(clk), .Q(\ram[155][4] ) );
  DFFHQX1 \ram_reg[155][3]  ( .D(n3065), .CK(clk), .Q(\ram[155][3] ) );
  DFFHQX1 \ram_reg[155][2]  ( .D(n3064), .CK(clk), .Q(\ram[155][2] ) );
  DFFHQX1 \ram_reg[155][1]  ( .D(n3063), .CK(clk), .Q(\ram[155][1] ) );
  DFFHQX1 \ram_reg[155][0]  ( .D(n3062), .CK(clk), .Q(\ram[155][0] ) );
  DFFHQX1 \ram_reg[151][15]  ( .D(n3013), .CK(clk), .Q(\ram[151][15] ) );
  DFFHQX1 \ram_reg[151][14]  ( .D(n3012), .CK(clk), .Q(\ram[151][14] ) );
  DFFHQX1 \ram_reg[151][13]  ( .D(n3011), .CK(clk), .Q(\ram[151][13] ) );
  DFFHQX1 \ram_reg[151][12]  ( .D(n3010), .CK(clk), .Q(\ram[151][12] ) );
  DFFHQX1 \ram_reg[151][11]  ( .D(n3009), .CK(clk), .Q(\ram[151][11] ) );
  DFFHQX1 \ram_reg[151][10]  ( .D(n3008), .CK(clk), .Q(\ram[151][10] ) );
  DFFHQX1 \ram_reg[151][9]  ( .D(n3007), .CK(clk), .Q(\ram[151][9] ) );
  DFFHQX1 \ram_reg[151][8]  ( .D(n3006), .CK(clk), .Q(\ram[151][8] ) );
  DFFHQX1 \ram_reg[151][7]  ( .D(n3005), .CK(clk), .Q(\ram[151][7] ) );
  DFFHQX1 \ram_reg[151][6]  ( .D(n3004), .CK(clk), .Q(\ram[151][6] ) );
  DFFHQX1 \ram_reg[151][5]  ( .D(n3003), .CK(clk), .Q(\ram[151][5] ) );
  DFFHQX1 \ram_reg[151][4]  ( .D(n3002), .CK(clk), .Q(\ram[151][4] ) );
  DFFHQX1 \ram_reg[151][3]  ( .D(n3001), .CK(clk), .Q(\ram[151][3] ) );
  DFFHQX1 \ram_reg[151][2]  ( .D(n3000), .CK(clk), .Q(\ram[151][2] ) );
  DFFHQX1 \ram_reg[151][1]  ( .D(n2999), .CK(clk), .Q(\ram[151][1] ) );
  DFFHQX1 \ram_reg[151][0]  ( .D(n2998), .CK(clk), .Q(\ram[151][0] ) );
  DFFHQX1 \ram_reg[147][15]  ( .D(n2949), .CK(clk), .Q(\ram[147][15] ) );
  DFFHQX1 \ram_reg[147][14]  ( .D(n2948), .CK(clk), .Q(\ram[147][14] ) );
  DFFHQX1 \ram_reg[147][13]  ( .D(n2947), .CK(clk), .Q(\ram[147][13] ) );
  DFFHQX1 \ram_reg[147][12]  ( .D(n2946), .CK(clk), .Q(\ram[147][12] ) );
  DFFHQX1 \ram_reg[147][11]  ( .D(n2945), .CK(clk), .Q(\ram[147][11] ) );
  DFFHQX1 \ram_reg[147][10]  ( .D(n2944), .CK(clk), .Q(\ram[147][10] ) );
  DFFHQX1 \ram_reg[147][9]  ( .D(n2943), .CK(clk), .Q(\ram[147][9] ) );
  DFFHQX1 \ram_reg[147][8]  ( .D(n2942), .CK(clk), .Q(\ram[147][8] ) );
  DFFHQX1 \ram_reg[147][7]  ( .D(n2941), .CK(clk), .Q(\ram[147][7] ) );
  DFFHQX1 \ram_reg[147][6]  ( .D(n2940), .CK(clk), .Q(\ram[147][6] ) );
  DFFHQX1 \ram_reg[147][5]  ( .D(n2939), .CK(clk), .Q(\ram[147][5] ) );
  DFFHQX1 \ram_reg[147][4]  ( .D(n2938), .CK(clk), .Q(\ram[147][4] ) );
  DFFHQX1 \ram_reg[147][3]  ( .D(n2937), .CK(clk), .Q(\ram[147][3] ) );
  DFFHQX1 \ram_reg[147][2]  ( .D(n2936), .CK(clk), .Q(\ram[147][2] ) );
  DFFHQX1 \ram_reg[147][1]  ( .D(n2935), .CK(clk), .Q(\ram[147][1] ) );
  DFFHQX1 \ram_reg[147][0]  ( .D(n2934), .CK(clk), .Q(\ram[147][0] ) );
  DFFHQX1 \ram_reg[143][15]  ( .D(n2885), .CK(clk), .Q(\ram[143][15] ) );
  DFFHQX1 \ram_reg[143][14]  ( .D(n2884), .CK(clk), .Q(\ram[143][14] ) );
  DFFHQX1 \ram_reg[143][13]  ( .D(n2883), .CK(clk), .Q(\ram[143][13] ) );
  DFFHQX1 \ram_reg[143][12]  ( .D(n2882), .CK(clk), .Q(\ram[143][12] ) );
  DFFHQX1 \ram_reg[143][11]  ( .D(n2881), .CK(clk), .Q(\ram[143][11] ) );
  DFFHQX1 \ram_reg[143][10]  ( .D(n2880), .CK(clk), .Q(\ram[143][10] ) );
  DFFHQX1 \ram_reg[143][9]  ( .D(n2879), .CK(clk), .Q(\ram[143][9] ) );
  DFFHQX1 \ram_reg[143][8]  ( .D(n2878), .CK(clk), .Q(\ram[143][8] ) );
  DFFHQX1 \ram_reg[143][7]  ( .D(n2877), .CK(clk), .Q(\ram[143][7] ) );
  DFFHQX1 \ram_reg[143][6]  ( .D(n2876), .CK(clk), .Q(\ram[143][6] ) );
  DFFHQX1 \ram_reg[143][5]  ( .D(n2875), .CK(clk), .Q(\ram[143][5] ) );
  DFFHQX1 \ram_reg[143][4]  ( .D(n2874), .CK(clk), .Q(\ram[143][4] ) );
  DFFHQX1 \ram_reg[143][3]  ( .D(n2873), .CK(clk), .Q(\ram[143][3] ) );
  DFFHQX1 \ram_reg[143][2]  ( .D(n2872), .CK(clk), .Q(\ram[143][2] ) );
  DFFHQX1 \ram_reg[143][1]  ( .D(n2871), .CK(clk), .Q(\ram[143][1] ) );
  DFFHQX1 \ram_reg[143][0]  ( .D(n2870), .CK(clk), .Q(\ram[143][0] ) );
  DFFHQX1 \ram_reg[139][15]  ( .D(n2821), .CK(clk), .Q(\ram[139][15] ) );
  DFFHQX1 \ram_reg[139][14]  ( .D(n2820), .CK(clk), .Q(\ram[139][14] ) );
  DFFHQX1 \ram_reg[139][13]  ( .D(n2819), .CK(clk), .Q(\ram[139][13] ) );
  DFFHQX1 \ram_reg[139][12]  ( .D(n2818), .CK(clk), .Q(\ram[139][12] ) );
  DFFHQX1 \ram_reg[139][11]  ( .D(n2817), .CK(clk), .Q(\ram[139][11] ) );
  DFFHQX1 \ram_reg[139][10]  ( .D(n2816), .CK(clk), .Q(\ram[139][10] ) );
  DFFHQX1 \ram_reg[139][9]  ( .D(n2815), .CK(clk), .Q(\ram[139][9] ) );
  DFFHQX1 \ram_reg[139][8]  ( .D(n2814), .CK(clk), .Q(\ram[139][8] ) );
  DFFHQX1 \ram_reg[139][7]  ( .D(n2813), .CK(clk), .Q(\ram[139][7] ) );
  DFFHQX1 \ram_reg[139][6]  ( .D(n2812), .CK(clk), .Q(\ram[139][6] ) );
  DFFHQX1 \ram_reg[139][5]  ( .D(n2811), .CK(clk), .Q(\ram[139][5] ) );
  DFFHQX1 \ram_reg[139][4]  ( .D(n2810), .CK(clk), .Q(\ram[139][4] ) );
  DFFHQX1 \ram_reg[139][3]  ( .D(n2809), .CK(clk), .Q(\ram[139][3] ) );
  DFFHQX1 \ram_reg[139][2]  ( .D(n2808), .CK(clk), .Q(\ram[139][2] ) );
  DFFHQX1 \ram_reg[139][1]  ( .D(n2807), .CK(clk), .Q(\ram[139][1] ) );
  DFFHQX1 \ram_reg[139][0]  ( .D(n2806), .CK(clk), .Q(\ram[139][0] ) );
  DFFHQX1 \ram_reg[135][15]  ( .D(n2757), .CK(clk), .Q(\ram[135][15] ) );
  DFFHQX1 \ram_reg[135][14]  ( .D(n2756), .CK(clk), .Q(\ram[135][14] ) );
  DFFHQX1 \ram_reg[135][13]  ( .D(n2755), .CK(clk), .Q(\ram[135][13] ) );
  DFFHQX1 \ram_reg[135][12]  ( .D(n2754), .CK(clk), .Q(\ram[135][12] ) );
  DFFHQX1 \ram_reg[135][11]  ( .D(n2753), .CK(clk), .Q(\ram[135][11] ) );
  DFFHQX1 \ram_reg[135][10]  ( .D(n2752), .CK(clk), .Q(\ram[135][10] ) );
  DFFHQX1 \ram_reg[135][9]  ( .D(n2751), .CK(clk), .Q(\ram[135][9] ) );
  DFFHQX1 \ram_reg[135][8]  ( .D(n2750), .CK(clk), .Q(\ram[135][8] ) );
  DFFHQX1 \ram_reg[135][7]  ( .D(n2749), .CK(clk), .Q(\ram[135][7] ) );
  DFFHQX1 \ram_reg[135][6]  ( .D(n2748), .CK(clk), .Q(\ram[135][6] ) );
  DFFHQX1 \ram_reg[135][5]  ( .D(n2747), .CK(clk), .Q(\ram[135][5] ) );
  DFFHQX1 \ram_reg[135][4]  ( .D(n2746), .CK(clk), .Q(\ram[135][4] ) );
  DFFHQX1 \ram_reg[135][3]  ( .D(n2745), .CK(clk), .Q(\ram[135][3] ) );
  DFFHQX1 \ram_reg[135][2]  ( .D(n2744), .CK(clk), .Q(\ram[135][2] ) );
  DFFHQX1 \ram_reg[135][1]  ( .D(n2743), .CK(clk), .Q(\ram[135][1] ) );
  DFFHQX1 \ram_reg[135][0]  ( .D(n2742), .CK(clk), .Q(\ram[135][0] ) );
  DFFHQX1 \ram_reg[131][15]  ( .D(n2693), .CK(clk), .Q(\ram[131][15] ) );
  DFFHQX1 \ram_reg[131][14]  ( .D(n2692), .CK(clk), .Q(\ram[131][14] ) );
  DFFHQX1 \ram_reg[131][13]  ( .D(n2691), .CK(clk), .Q(\ram[131][13] ) );
  DFFHQX1 \ram_reg[131][12]  ( .D(n2690), .CK(clk), .Q(\ram[131][12] ) );
  DFFHQX1 \ram_reg[131][11]  ( .D(n2689), .CK(clk), .Q(\ram[131][11] ) );
  DFFHQX1 \ram_reg[131][10]  ( .D(n2688), .CK(clk), .Q(\ram[131][10] ) );
  DFFHQX1 \ram_reg[131][9]  ( .D(n2687), .CK(clk), .Q(\ram[131][9] ) );
  DFFHQX1 \ram_reg[131][8]  ( .D(n2686), .CK(clk), .Q(\ram[131][8] ) );
  DFFHQX1 \ram_reg[131][7]  ( .D(n2685), .CK(clk), .Q(\ram[131][7] ) );
  DFFHQX1 \ram_reg[131][6]  ( .D(n2684), .CK(clk), .Q(\ram[131][6] ) );
  DFFHQX1 \ram_reg[131][5]  ( .D(n2683), .CK(clk), .Q(\ram[131][5] ) );
  DFFHQX1 \ram_reg[131][4]  ( .D(n2682), .CK(clk), .Q(\ram[131][4] ) );
  DFFHQX1 \ram_reg[131][3]  ( .D(n2681), .CK(clk), .Q(\ram[131][3] ) );
  DFFHQX1 \ram_reg[131][2]  ( .D(n2680), .CK(clk), .Q(\ram[131][2] ) );
  DFFHQX1 \ram_reg[131][1]  ( .D(n2679), .CK(clk), .Q(\ram[131][1] ) );
  DFFHQX1 \ram_reg[131][0]  ( .D(n2678), .CK(clk), .Q(\ram[131][0] ) );
  DFFHQX1 \ram_reg[127][15]  ( .D(n2629), .CK(clk), .Q(\ram[127][15] ) );
  DFFHQX1 \ram_reg[127][14]  ( .D(n2628), .CK(clk), .Q(\ram[127][14] ) );
  DFFHQX1 \ram_reg[127][13]  ( .D(n2627), .CK(clk), .Q(\ram[127][13] ) );
  DFFHQX1 \ram_reg[127][12]  ( .D(n2626), .CK(clk), .Q(\ram[127][12] ) );
  DFFHQX1 \ram_reg[127][11]  ( .D(n2625), .CK(clk), .Q(\ram[127][11] ) );
  DFFHQX1 \ram_reg[127][10]  ( .D(n2624), .CK(clk), .Q(\ram[127][10] ) );
  DFFHQX1 \ram_reg[127][9]  ( .D(n2623), .CK(clk), .Q(\ram[127][9] ) );
  DFFHQX1 \ram_reg[127][8]  ( .D(n2622), .CK(clk), .Q(\ram[127][8] ) );
  DFFHQX1 \ram_reg[127][7]  ( .D(n2621), .CK(clk), .Q(\ram[127][7] ) );
  DFFHQX1 \ram_reg[127][6]  ( .D(n2620), .CK(clk), .Q(\ram[127][6] ) );
  DFFHQX1 \ram_reg[127][5]  ( .D(n2619), .CK(clk), .Q(\ram[127][5] ) );
  DFFHQX1 \ram_reg[127][4]  ( .D(n2618), .CK(clk), .Q(\ram[127][4] ) );
  DFFHQX1 \ram_reg[127][3]  ( .D(n2617), .CK(clk), .Q(\ram[127][3] ) );
  DFFHQX1 \ram_reg[127][2]  ( .D(n2616), .CK(clk), .Q(\ram[127][2] ) );
  DFFHQX1 \ram_reg[127][1]  ( .D(n2615), .CK(clk), .Q(\ram[127][1] ) );
  DFFHQX1 \ram_reg[127][0]  ( .D(n2614), .CK(clk), .Q(\ram[127][0] ) );
  DFFHQX1 \ram_reg[123][15]  ( .D(n2565), .CK(clk), .Q(\ram[123][15] ) );
  DFFHQX1 \ram_reg[123][14]  ( .D(n2564), .CK(clk), .Q(\ram[123][14] ) );
  DFFHQX1 \ram_reg[123][13]  ( .D(n2563), .CK(clk), .Q(\ram[123][13] ) );
  DFFHQX1 \ram_reg[123][12]  ( .D(n2562), .CK(clk), .Q(\ram[123][12] ) );
  DFFHQX1 \ram_reg[123][11]  ( .D(n2561), .CK(clk), .Q(\ram[123][11] ) );
  DFFHQX1 \ram_reg[123][10]  ( .D(n2560), .CK(clk), .Q(\ram[123][10] ) );
  DFFHQX1 \ram_reg[123][9]  ( .D(n2559), .CK(clk), .Q(\ram[123][9] ) );
  DFFHQX1 \ram_reg[123][8]  ( .D(n2558), .CK(clk), .Q(\ram[123][8] ) );
  DFFHQX1 \ram_reg[123][7]  ( .D(n2557), .CK(clk), .Q(\ram[123][7] ) );
  DFFHQX1 \ram_reg[123][6]  ( .D(n2556), .CK(clk), .Q(\ram[123][6] ) );
  DFFHQX1 \ram_reg[123][5]  ( .D(n2555), .CK(clk), .Q(\ram[123][5] ) );
  DFFHQX1 \ram_reg[123][4]  ( .D(n2554), .CK(clk), .Q(\ram[123][4] ) );
  DFFHQX1 \ram_reg[123][3]  ( .D(n2553), .CK(clk), .Q(\ram[123][3] ) );
  DFFHQX1 \ram_reg[123][2]  ( .D(n2552), .CK(clk), .Q(\ram[123][2] ) );
  DFFHQX1 \ram_reg[123][1]  ( .D(n2551), .CK(clk), .Q(\ram[123][1] ) );
  DFFHQX1 \ram_reg[123][0]  ( .D(n2550), .CK(clk), .Q(\ram[123][0] ) );
  DFFHQX1 \ram_reg[119][15]  ( .D(n2501), .CK(clk), .Q(\ram[119][15] ) );
  DFFHQX1 \ram_reg[119][14]  ( .D(n2500), .CK(clk), .Q(\ram[119][14] ) );
  DFFHQX1 \ram_reg[119][13]  ( .D(n2499), .CK(clk), .Q(\ram[119][13] ) );
  DFFHQX1 \ram_reg[119][12]  ( .D(n2498), .CK(clk), .Q(\ram[119][12] ) );
  DFFHQX1 \ram_reg[119][11]  ( .D(n2497), .CK(clk), .Q(\ram[119][11] ) );
  DFFHQX1 \ram_reg[119][10]  ( .D(n2496), .CK(clk), .Q(\ram[119][10] ) );
  DFFHQX1 \ram_reg[119][9]  ( .D(n2495), .CK(clk), .Q(\ram[119][9] ) );
  DFFHQX1 \ram_reg[119][8]  ( .D(n2494), .CK(clk), .Q(\ram[119][8] ) );
  DFFHQX1 \ram_reg[119][7]  ( .D(n2493), .CK(clk), .Q(\ram[119][7] ) );
  DFFHQX1 \ram_reg[119][6]  ( .D(n2492), .CK(clk), .Q(\ram[119][6] ) );
  DFFHQX1 \ram_reg[119][5]  ( .D(n2491), .CK(clk), .Q(\ram[119][5] ) );
  DFFHQX1 \ram_reg[119][4]  ( .D(n2490), .CK(clk), .Q(\ram[119][4] ) );
  DFFHQX1 \ram_reg[119][3]  ( .D(n2489), .CK(clk), .Q(\ram[119][3] ) );
  DFFHQX1 \ram_reg[119][2]  ( .D(n2488), .CK(clk), .Q(\ram[119][2] ) );
  DFFHQX1 \ram_reg[119][1]  ( .D(n2487), .CK(clk), .Q(\ram[119][1] ) );
  DFFHQX1 \ram_reg[119][0]  ( .D(n2486), .CK(clk), .Q(\ram[119][0] ) );
  DFFHQX1 \ram_reg[115][15]  ( .D(n2437), .CK(clk), .Q(\ram[115][15] ) );
  DFFHQX1 \ram_reg[115][14]  ( .D(n2436), .CK(clk), .Q(\ram[115][14] ) );
  DFFHQX1 \ram_reg[115][13]  ( .D(n2435), .CK(clk), .Q(\ram[115][13] ) );
  DFFHQX1 \ram_reg[115][12]  ( .D(n2434), .CK(clk), .Q(\ram[115][12] ) );
  DFFHQX1 \ram_reg[115][11]  ( .D(n2433), .CK(clk), .Q(\ram[115][11] ) );
  DFFHQX1 \ram_reg[115][10]  ( .D(n2432), .CK(clk), .Q(\ram[115][10] ) );
  DFFHQX1 \ram_reg[115][9]  ( .D(n2431), .CK(clk), .Q(\ram[115][9] ) );
  DFFHQX1 \ram_reg[115][8]  ( .D(n2430), .CK(clk), .Q(\ram[115][8] ) );
  DFFHQX1 \ram_reg[115][7]  ( .D(n2429), .CK(clk), .Q(\ram[115][7] ) );
  DFFHQX1 \ram_reg[115][6]  ( .D(n2428), .CK(clk), .Q(\ram[115][6] ) );
  DFFHQX1 \ram_reg[115][5]  ( .D(n2427), .CK(clk), .Q(\ram[115][5] ) );
  DFFHQX1 \ram_reg[115][4]  ( .D(n2426), .CK(clk), .Q(\ram[115][4] ) );
  DFFHQX1 \ram_reg[115][3]  ( .D(n2425), .CK(clk), .Q(\ram[115][3] ) );
  DFFHQX1 \ram_reg[115][2]  ( .D(n2424), .CK(clk), .Q(\ram[115][2] ) );
  DFFHQX1 \ram_reg[115][1]  ( .D(n2423), .CK(clk), .Q(\ram[115][1] ) );
  DFFHQX1 \ram_reg[115][0]  ( .D(n2422), .CK(clk), .Q(\ram[115][0] ) );
  DFFHQX1 \ram_reg[111][15]  ( .D(n2373), .CK(clk), .Q(\ram[111][15] ) );
  DFFHQX1 \ram_reg[111][14]  ( .D(n2372), .CK(clk), .Q(\ram[111][14] ) );
  DFFHQX1 \ram_reg[111][13]  ( .D(n2371), .CK(clk), .Q(\ram[111][13] ) );
  DFFHQX1 \ram_reg[111][12]  ( .D(n2370), .CK(clk), .Q(\ram[111][12] ) );
  DFFHQX1 \ram_reg[111][11]  ( .D(n2369), .CK(clk), .Q(\ram[111][11] ) );
  DFFHQX1 \ram_reg[111][10]  ( .D(n2368), .CK(clk), .Q(\ram[111][10] ) );
  DFFHQX1 \ram_reg[111][9]  ( .D(n2367), .CK(clk), .Q(\ram[111][9] ) );
  DFFHQX1 \ram_reg[111][8]  ( .D(n2366), .CK(clk), .Q(\ram[111][8] ) );
  DFFHQX1 \ram_reg[111][7]  ( .D(n2365), .CK(clk), .Q(\ram[111][7] ) );
  DFFHQX1 \ram_reg[111][6]  ( .D(n2364), .CK(clk), .Q(\ram[111][6] ) );
  DFFHQX1 \ram_reg[111][5]  ( .D(n2363), .CK(clk), .Q(\ram[111][5] ) );
  DFFHQX1 \ram_reg[111][4]  ( .D(n2362), .CK(clk), .Q(\ram[111][4] ) );
  DFFHQX1 \ram_reg[111][3]  ( .D(n2361), .CK(clk), .Q(\ram[111][3] ) );
  DFFHQX1 \ram_reg[111][2]  ( .D(n2360), .CK(clk), .Q(\ram[111][2] ) );
  DFFHQX1 \ram_reg[111][1]  ( .D(n2359), .CK(clk), .Q(\ram[111][1] ) );
  DFFHQX1 \ram_reg[111][0]  ( .D(n2358), .CK(clk), .Q(\ram[111][0] ) );
  DFFHQX1 \ram_reg[107][15]  ( .D(n2309), .CK(clk), .Q(\ram[107][15] ) );
  DFFHQX1 \ram_reg[107][14]  ( .D(n2308), .CK(clk), .Q(\ram[107][14] ) );
  DFFHQX1 \ram_reg[107][13]  ( .D(n2307), .CK(clk), .Q(\ram[107][13] ) );
  DFFHQX1 \ram_reg[107][12]  ( .D(n2306), .CK(clk), .Q(\ram[107][12] ) );
  DFFHQX1 \ram_reg[107][11]  ( .D(n2305), .CK(clk), .Q(\ram[107][11] ) );
  DFFHQX1 \ram_reg[107][10]  ( .D(n2304), .CK(clk), .Q(\ram[107][10] ) );
  DFFHQX1 \ram_reg[107][9]  ( .D(n2303), .CK(clk), .Q(\ram[107][9] ) );
  DFFHQX1 \ram_reg[107][8]  ( .D(n2302), .CK(clk), .Q(\ram[107][8] ) );
  DFFHQX1 \ram_reg[107][7]  ( .D(n2301), .CK(clk), .Q(\ram[107][7] ) );
  DFFHQX1 \ram_reg[107][6]  ( .D(n2300), .CK(clk), .Q(\ram[107][6] ) );
  DFFHQX1 \ram_reg[107][5]  ( .D(n2299), .CK(clk), .Q(\ram[107][5] ) );
  DFFHQX1 \ram_reg[107][4]  ( .D(n2298), .CK(clk), .Q(\ram[107][4] ) );
  DFFHQX1 \ram_reg[107][3]  ( .D(n2297), .CK(clk), .Q(\ram[107][3] ) );
  DFFHQX1 \ram_reg[107][2]  ( .D(n2296), .CK(clk), .Q(\ram[107][2] ) );
  DFFHQX1 \ram_reg[107][1]  ( .D(n2295), .CK(clk), .Q(\ram[107][1] ) );
  DFFHQX1 \ram_reg[107][0]  ( .D(n2294), .CK(clk), .Q(\ram[107][0] ) );
  DFFHQX1 \ram_reg[103][15]  ( .D(n2245), .CK(clk), .Q(\ram[103][15] ) );
  DFFHQX1 \ram_reg[103][14]  ( .D(n2244), .CK(clk), .Q(\ram[103][14] ) );
  DFFHQX1 \ram_reg[103][13]  ( .D(n2243), .CK(clk), .Q(\ram[103][13] ) );
  DFFHQX1 \ram_reg[103][12]  ( .D(n2242), .CK(clk), .Q(\ram[103][12] ) );
  DFFHQX1 \ram_reg[103][11]  ( .D(n2241), .CK(clk), .Q(\ram[103][11] ) );
  DFFHQX1 \ram_reg[103][10]  ( .D(n2240), .CK(clk), .Q(\ram[103][10] ) );
  DFFHQX1 \ram_reg[103][9]  ( .D(n2239), .CK(clk), .Q(\ram[103][9] ) );
  DFFHQX1 \ram_reg[103][8]  ( .D(n2238), .CK(clk), .Q(\ram[103][8] ) );
  DFFHQX1 \ram_reg[103][7]  ( .D(n2237), .CK(clk), .Q(\ram[103][7] ) );
  DFFHQX1 \ram_reg[103][6]  ( .D(n2236), .CK(clk), .Q(\ram[103][6] ) );
  DFFHQX1 \ram_reg[103][5]  ( .D(n2235), .CK(clk), .Q(\ram[103][5] ) );
  DFFHQX1 \ram_reg[103][4]  ( .D(n2234), .CK(clk), .Q(\ram[103][4] ) );
  DFFHQX1 \ram_reg[103][3]  ( .D(n2233), .CK(clk), .Q(\ram[103][3] ) );
  DFFHQX1 \ram_reg[103][2]  ( .D(n2232), .CK(clk), .Q(\ram[103][2] ) );
  DFFHQX1 \ram_reg[103][1]  ( .D(n2231), .CK(clk), .Q(\ram[103][1] ) );
  DFFHQX1 \ram_reg[103][0]  ( .D(n2230), .CK(clk), .Q(\ram[103][0] ) );
  DFFHQX1 \ram_reg[99][15]  ( .D(n2181), .CK(clk), .Q(\ram[99][15] ) );
  DFFHQX1 \ram_reg[99][14]  ( .D(n2180), .CK(clk), .Q(\ram[99][14] ) );
  DFFHQX1 \ram_reg[99][13]  ( .D(n2179), .CK(clk), .Q(\ram[99][13] ) );
  DFFHQX1 \ram_reg[99][12]  ( .D(n2178), .CK(clk), .Q(\ram[99][12] ) );
  DFFHQX1 \ram_reg[99][11]  ( .D(n2177), .CK(clk), .Q(\ram[99][11] ) );
  DFFHQX1 \ram_reg[99][10]  ( .D(n2176), .CK(clk), .Q(\ram[99][10] ) );
  DFFHQX1 \ram_reg[99][9]  ( .D(n2175), .CK(clk), .Q(\ram[99][9] ) );
  DFFHQX1 \ram_reg[99][8]  ( .D(n2174), .CK(clk), .Q(\ram[99][8] ) );
  DFFHQX1 \ram_reg[99][7]  ( .D(n2173), .CK(clk), .Q(\ram[99][7] ) );
  DFFHQX1 \ram_reg[99][6]  ( .D(n2172), .CK(clk), .Q(\ram[99][6] ) );
  DFFHQX1 \ram_reg[99][5]  ( .D(n2171), .CK(clk), .Q(\ram[99][5] ) );
  DFFHQX1 \ram_reg[99][4]  ( .D(n2170), .CK(clk), .Q(\ram[99][4] ) );
  DFFHQX1 \ram_reg[99][3]  ( .D(n2169), .CK(clk), .Q(\ram[99][3] ) );
  DFFHQX1 \ram_reg[99][2]  ( .D(n2168), .CK(clk), .Q(\ram[99][2] ) );
  DFFHQX1 \ram_reg[99][1]  ( .D(n2167), .CK(clk), .Q(\ram[99][1] ) );
  DFFHQX1 \ram_reg[99][0]  ( .D(n2166), .CK(clk), .Q(\ram[99][0] ) );
  DFFHQX1 \ram_reg[95][15]  ( .D(n2117), .CK(clk), .Q(\ram[95][15] ) );
  DFFHQX1 \ram_reg[95][14]  ( .D(n2116), .CK(clk), .Q(\ram[95][14] ) );
  DFFHQX1 \ram_reg[95][13]  ( .D(n2115), .CK(clk), .Q(\ram[95][13] ) );
  DFFHQX1 \ram_reg[95][12]  ( .D(n2114), .CK(clk), .Q(\ram[95][12] ) );
  DFFHQX1 \ram_reg[95][11]  ( .D(n2113), .CK(clk), .Q(\ram[95][11] ) );
  DFFHQX1 \ram_reg[95][10]  ( .D(n2112), .CK(clk), .Q(\ram[95][10] ) );
  DFFHQX1 \ram_reg[95][9]  ( .D(n2111), .CK(clk), .Q(\ram[95][9] ) );
  DFFHQX1 \ram_reg[95][8]  ( .D(n2110), .CK(clk), .Q(\ram[95][8] ) );
  DFFHQX1 \ram_reg[95][7]  ( .D(n2109), .CK(clk), .Q(\ram[95][7] ) );
  DFFHQX1 \ram_reg[95][6]  ( .D(n2108), .CK(clk), .Q(\ram[95][6] ) );
  DFFHQX1 \ram_reg[95][5]  ( .D(n2107), .CK(clk), .Q(\ram[95][5] ) );
  DFFHQX1 \ram_reg[95][4]  ( .D(n2106), .CK(clk), .Q(\ram[95][4] ) );
  DFFHQX1 \ram_reg[95][3]  ( .D(n2105), .CK(clk), .Q(\ram[95][3] ) );
  DFFHQX1 \ram_reg[95][2]  ( .D(n2104), .CK(clk), .Q(\ram[95][2] ) );
  DFFHQX1 \ram_reg[95][1]  ( .D(n2103), .CK(clk), .Q(\ram[95][1] ) );
  DFFHQX1 \ram_reg[95][0]  ( .D(n2102), .CK(clk), .Q(\ram[95][0] ) );
  DFFHQX1 \ram_reg[91][15]  ( .D(n2053), .CK(clk), .Q(\ram[91][15] ) );
  DFFHQX1 \ram_reg[91][14]  ( .D(n2052), .CK(clk), .Q(\ram[91][14] ) );
  DFFHQX1 \ram_reg[91][13]  ( .D(n2051), .CK(clk), .Q(\ram[91][13] ) );
  DFFHQX1 \ram_reg[91][12]  ( .D(n2050), .CK(clk), .Q(\ram[91][12] ) );
  DFFHQX1 \ram_reg[91][11]  ( .D(n2049), .CK(clk), .Q(\ram[91][11] ) );
  DFFHQX1 \ram_reg[91][10]  ( .D(n2048), .CK(clk), .Q(\ram[91][10] ) );
  DFFHQX1 \ram_reg[91][9]  ( .D(n2047), .CK(clk), .Q(\ram[91][9] ) );
  DFFHQX1 \ram_reg[91][8]  ( .D(n2046), .CK(clk), .Q(\ram[91][8] ) );
  DFFHQX1 \ram_reg[91][7]  ( .D(n2045), .CK(clk), .Q(\ram[91][7] ) );
  DFFHQX1 \ram_reg[91][6]  ( .D(n2044), .CK(clk), .Q(\ram[91][6] ) );
  DFFHQX1 \ram_reg[91][5]  ( .D(n2043), .CK(clk), .Q(\ram[91][5] ) );
  DFFHQX1 \ram_reg[91][4]  ( .D(n2042), .CK(clk), .Q(\ram[91][4] ) );
  DFFHQX1 \ram_reg[91][3]  ( .D(n2041), .CK(clk), .Q(\ram[91][3] ) );
  DFFHQX1 \ram_reg[91][2]  ( .D(n2040), .CK(clk), .Q(\ram[91][2] ) );
  DFFHQX1 \ram_reg[91][1]  ( .D(n2039), .CK(clk), .Q(\ram[91][1] ) );
  DFFHQX1 \ram_reg[91][0]  ( .D(n2038), .CK(clk), .Q(\ram[91][0] ) );
  DFFHQX1 \ram_reg[87][15]  ( .D(n1989), .CK(clk), .Q(\ram[87][15] ) );
  DFFHQX1 \ram_reg[87][14]  ( .D(n1988), .CK(clk), .Q(\ram[87][14] ) );
  DFFHQX1 \ram_reg[87][13]  ( .D(n1987), .CK(clk), .Q(\ram[87][13] ) );
  DFFHQX1 \ram_reg[87][12]  ( .D(n1986), .CK(clk), .Q(\ram[87][12] ) );
  DFFHQX1 \ram_reg[87][11]  ( .D(n1985), .CK(clk), .Q(\ram[87][11] ) );
  DFFHQX1 \ram_reg[87][10]  ( .D(n1984), .CK(clk), .Q(\ram[87][10] ) );
  DFFHQX1 \ram_reg[87][9]  ( .D(n1983), .CK(clk), .Q(\ram[87][9] ) );
  DFFHQX1 \ram_reg[87][8]  ( .D(n1982), .CK(clk), .Q(\ram[87][8] ) );
  DFFHQX1 \ram_reg[87][7]  ( .D(n1981), .CK(clk), .Q(\ram[87][7] ) );
  DFFHQX1 \ram_reg[87][6]  ( .D(n1980), .CK(clk), .Q(\ram[87][6] ) );
  DFFHQX1 \ram_reg[87][5]  ( .D(n1979), .CK(clk), .Q(\ram[87][5] ) );
  DFFHQX1 \ram_reg[87][4]  ( .D(n1978), .CK(clk), .Q(\ram[87][4] ) );
  DFFHQX1 \ram_reg[87][3]  ( .D(n1977), .CK(clk), .Q(\ram[87][3] ) );
  DFFHQX1 \ram_reg[87][2]  ( .D(n1976), .CK(clk), .Q(\ram[87][2] ) );
  DFFHQX1 \ram_reg[87][1]  ( .D(n1975), .CK(clk), .Q(\ram[87][1] ) );
  DFFHQX1 \ram_reg[87][0]  ( .D(n1974), .CK(clk), .Q(\ram[87][0] ) );
  DFFHQX1 \ram_reg[83][15]  ( .D(n1925), .CK(clk), .Q(\ram[83][15] ) );
  DFFHQX1 \ram_reg[83][14]  ( .D(n1924), .CK(clk), .Q(\ram[83][14] ) );
  DFFHQX1 \ram_reg[83][13]  ( .D(n1923), .CK(clk), .Q(\ram[83][13] ) );
  DFFHQX1 \ram_reg[83][12]  ( .D(n1922), .CK(clk), .Q(\ram[83][12] ) );
  DFFHQX1 \ram_reg[83][11]  ( .D(n1921), .CK(clk), .Q(\ram[83][11] ) );
  DFFHQX1 \ram_reg[83][10]  ( .D(n1920), .CK(clk), .Q(\ram[83][10] ) );
  DFFHQX1 \ram_reg[83][9]  ( .D(n1919), .CK(clk), .Q(\ram[83][9] ) );
  DFFHQX1 \ram_reg[83][8]  ( .D(n1918), .CK(clk), .Q(\ram[83][8] ) );
  DFFHQX1 \ram_reg[83][7]  ( .D(n1917), .CK(clk), .Q(\ram[83][7] ) );
  DFFHQX1 \ram_reg[83][6]  ( .D(n1916), .CK(clk), .Q(\ram[83][6] ) );
  DFFHQX1 \ram_reg[83][5]  ( .D(n1915), .CK(clk), .Q(\ram[83][5] ) );
  DFFHQX1 \ram_reg[83][4]  ( .D(n1914), .CK(clk), .Q(\ram[83][4] ) );
  DFFHQX1 \ram_reg[83][3]  ( .D(n1913), .CK(clk), .Q(\ram[83][3] ) );
  DFFHQX1 \ram_reg[83][2]  ( .D(n1912), .CK(clk), .Q(\ram[83][2] ) );
  DFFHQX1 \ram_reg[83][1]  ( .D(n1911), .CK(clk), .Q(\ram[83][1] ) );
  DFFHQX1 \ram_reg[83][0]  ( .D(n1910), .CK(clk), .Q(\ram[83][0] ) );
  DFFHQX1 \ram_reg[79][15]  ( .D(n1861), .CK(clk), .Q(\ram[79][15] ) );
  DFFHQX1 \ram_reg[79][14]  ( .D(n1860), .CK(clk), .Q(\ram[79][14] ) );
  DFFHQX1 \ram_reg[79][13]  ( .D(n1859), .CK(clk), .Q(\ram[79][13] ) );
  DFFHQX1 \ram_reg[79][12]  ( .D(n1858), .CK(clk), .Q(\ram[79][12] ) );
  DFFHQX1 \ram_reg[79][11]  ( .D(n1857), .CK(clk), .Q(\ram[79][11] ) );
  DFFHQX1 \ram_reg[79][10]  ( .D(n1856), .CK(clk), .Q(\ram[79][10] ) );
  DFFHQX1 \ram_reg[79][9]  ( .D(n1855), .CK(clk), .Q(\ram[79][9] ) );
  DFFHQX1 \ram_reg[79][8]  ( .D(n1854), .CK(clk), .Q(\ram[79][8] ) );
  DFFHQX1 \ram_reg[79][7]  ( .D(n1853), .CK(clk), .Q(\ram[79][7] ) );
  DFFHQX1 \ram_reg[79][6]  ( .D(n1852), .CK(clk), .Q(\ram[79][6] ) );
  DFFHQX1 \ram_reg[79][5]  ( .D(n1851), .CK(clk), .Q(\ram[79][5] ) );
  DFFHQX1 \ram_reg[79][4]  ( .D(n1850), .CK(clk), .Q(\ram[79][4] ) );
  DFFHQX1 \ram_reg[79][3]  ( .D(n1849), .CK(clk), .Q(\ram[79][3] ) );
  DFFHQX1 \ram_reg[79][2]  ( .D(n1848), .CK(clk), .Q(\ram[79][2] ) );
  DFFHQX1 \ram_reg[79][1]  ( .D(n1847), .CK(clk), .Q(\ram[79][1] ) );
  DFFHQX1 \ram_reg[79][0]  ( .D(n1846), .CK(clk), .Q(\ram[79][0] ) );
  DFFHQX1 \ram_reg[75][15]  ( .D(n1797), .CK(clk), .Q(\ram[75][15] ) );
  DFFHQX1 \ram_reg[75][14]  ( .D(n1796), .CK(clk), .Q(\ram[75][14] ) );
  DFFHQX1 \ram_reg[75][13]  ( .D(n1795), .CK(clk), .Q(\ram[75][13] ) );
  DFFHQX1 \ram_reg[75][12]  ( .D(n1794), .CK(clk), .Q(\ram[75][12] ) );
  DFFHQX1 \ram_reg[75][11]  ( .D(n1793), .CK(clk), .Q(\ram[75][11] ) );
  DFFHQX1 \ram_reg[75][10]  ( .D(n1792), .CK(clk), .Q(\ram[75][10] ) );
  DFFHQX1 \ram_reg[75][9]  ( .D(n1791), .CK(clk), .Q(\ram[75][9] ) );
  DFFHQX1 \ram_reg[75][8]  ( .D(n1790), .CK(clk), .Q(\ram[75][8] ) );
  DFFHQX1 \ram_reg[75][7]  ( .D(n1789), .CK(clk), .Q(\ram[75][7] ) );
  DFFHQX1 \ram_reg[75][6]  ( .D(n1788), .CK(clk), .Q(\ram[75][6] ) );
  DFFHQX1 \ram_reg[75][5]  ( .D(n1787), .CK(clk), .Q(\ram[75][5] ) );
  DFFHQX1 \ram_reg[75][4]  ( .D(n1786), .CK(clk), .Q(\ram[75][4] ) );
  DFFHQX1 \ram_reg[75][3]  ( .D(n1785), .CK(clk), .Q(\ram[75][3] ) );
  DFFHQX1 \ram_reg[75][2]  ( .D(n1784), .CK(clk), .Q(\ram[75][2] ) );
  DFFHQX1 \ram_reg[75][1]  ( .D(n1783), .CK(clk), .Q(\ram[75][1] ) );
  DFFHQX1 \ram_reg[75][0]  ( .D(n1782), .CK(clk), .Q(\ram[75][0] ) );
  DFFHQX1 \ram_reg[71][15]  ( .D(n1733), .CK(clk), .Q(\ram[71][15] ) );
  DFFHQX1 \ram_reg[71][14]  ( .D(n1732), .CK(clk), .Q(\ram[71][14] ) );
  DFFHQX1 \ram_reg[71][13]  ( .D(n1731), .CK(clk), .Q(\ram[71][13] ) );
  DFFHQX1 \ram_reg[71][12]  ( .D(n1730), .CK(clk), .Q(\ram[71][12] ) );
  DFFHQX1 \ram_reg[71][11]  ( .D(n1729), .CK(clk), .Q(\ram[71][11] ) );
  DFFHQX1 \ram_reg[71][10]  ( .D(n1728), .CK(clk), .Q(\ram[71][10] ) );
  DFFHQX1 \ram_reg[71][9]  ( .D(n1727), .CK(clk), .Q(\ram[71][9] ) );
  DFFHQX1 \ram_reg[71][8]  ( .D(n1726), .CK(clk), .Q(\ram[71][8] ) );
  DFFHQX1 \ram_reg[71][7]  ( .D(n1725), .CK(clk), .Q(\ram[71][7] ) );
  DFFHQX1 \ram_reg[71][6]  ( .D(n1724), .CK(clk), .Q(\ram[71][6] ) );
  DFFHQX1 \ram_reg[71][5]  ( .D(n1723), .CK(clk), .Q(\ram[71][5] ) );
  DFFHQX1 \ram_reg[71][4]  ( .D(n1722), .CK(clk), .Q(\ram[71][4] ) );
  DFFHQX1 \ram_reg[71][3]  ( .D(n1721), .CK(clk), .Q(\ram[71][3] ) );
  DFFHQX1 \ram_reg[71][2]  ( .D(n1720), .CK(clk), .Q(\ram[71][2] ) );
  DFFHQX1 \ram_reg[71][1]  ( .D(n1719), .CK(clk), .Q(\ram[71][1] ) );
  DFFHQX1 \ram_reg[71][0]  ( .D(n1718), .CK(clk), .Q(\ram[71][0] ) );
  DFFHQX1 \ram_reg[67][15]  ( .D(n1669), .CK(clk), .Q(\ram[67][15] ) );
  DFFHQX1 \ram_reg[67][14]  ( .D(n1668), .CK(clk), .Q(\ram[67][14] ) );
  DFFHQX1 \ram_reg[67][13]  ( .D(n1667), .CK(clk), .Q(\ram[67][13] ) );
  DFFHQX1 \ram_reg[67][12]  ( .D(n1666), .CK(clk), .Q(\ram[67][12] ) );
  DFFHQX1 \ram_reg[67][11]  ( .D(n1665), .CK(clk), .Q(\ram[67][11] ) );
  DFFHQX1 \ram_reg[67][10]  ( .D(n1664), .CK(clk), .Q(\ram[67][10] ) );
  DFFHQX1 \ram_reg[67][9]  ( .D(n1663), .CK(clk), .Q(\ram[67][9] ) );
  DFFHQX1 \ram_reg[67][8]  ( .D(n1662), .CK(clk), .Q(\ram[67][8] ) );
  DFFHQX1 \ram_reg[67][7]  ( .D(n1661), .CK(clk), .Q(\ram[67][7] ) );
  DFFHQX1 \ram_reg[67][6]  ( .D(n1660), .CK(clk), .Q(\ram[67][6] ) );
  DFFHQX1 \ram_reg[67][5]  ( .D(n1659), .CK(clk), .Q(\ram[67][5] ) );
  DFFHQX1 \ram_reg[67][4]  ( .D(n1658), .CK(clk), .Q(\ram[67][4] ) );
  DFFHQX1 \ram_reg[67][3]  ( .D(n1657), .CK(clk), .Q(\ram[67][3] ) );
  DFFHQX1 \ram_reg[67][2]  ( .D(n1656), .CK(clk), .Q(\ram[67][2] ) );
  DFFHQX1 \ram_reg[67][1]  ( .D(n1655), .CK(clk), .Q(\ram[67][1] ) );
  DFFHQX1 \ram_reg[67][0]  ( .D(n1654), .CK(clk), .Q(\ram[67][0] ) );
  DFFHQX1 \ram_reg[63][15]  ( .D(n1605), .CK(clk), .Q(\ram[63][15] ) );
  DFFHQX1 \ram_reg[63][14]  ( .D(n1604), .CK(clk), .Q(\ram[63][14] ) );
  DFFHQX1 \ram_reg[63][13]  ( .D(n1603), .CK(clk), .Q(\ram[63][13] ) );
  DFFHQX1 \ram_reg[63][12]  ( .D(n1602), .CK(clk), .Q(\ram[63][12] ) );
  DFFHQX1 \ram_reg[63][11]  ( .D(n1601), .CK(clk), .Q(\ram[63][11] ) );
  DFFHQX1 \ram_reg[63][10]  ( .D(n1600), .CK(clk), .Q(\ram[63][10] ) );
  DFFHQX1 \ram_reg[63][9]  ( .D(n1599), .CK(clk), .Q(\ram[63][9] ) );
  DFFHQX1 \ram_reg[63][8]  ( .D(n1598), .CK(clk), .Q(\ram[63][8] ) );
  DFFHQX1 \ram_reg[63][7]  ( .D(n1597), .CK(clk), .Q(\ram[63][7] ) );
  DFFHQX1 \ram_reg[63][6]  ( .D(n1596), .CK(clk), .Q(\ram[63][6] ) );
  DFFHQX1 \ram_reg[63][5]  ( .D(n1595), .CK(clk), .Q(\ram[63][5] ) );
  DFFHQX1 \ram_reg[63][4]  ( .D(n1594), .CK(clk), .Q(\ram[63][4] ) );
  DFFHQX1 \ram_reg[63][3]  ( .D(n1593), .CK(clk), .Q(\ram[63][3] ) );
  DFFHQX1 \ram_reg[63][2]  ( .D(n1592), .CK(clk), .Q(\ram[63][2] ) );
  DFFHQX1 \ram_reg[63][1]  ( .D(n1591), .CK(clk), .Q(\ram[63][1] ) );
  DFFHQX1 \ram_reg[63][0]  ( .D(n1590), .CK(clk), .Q(\ram[63][0] ) );
  DFFHQX1 \ram_reg[59][15]  ( .D(n1541), .CK(clk), .Q(\ram[59][15] ) );
  DFFHQX1 \ram_reg[59][14]  ( .D(n1540), .CK(clk), .Q(\ram[59][14] ) );
  DFFHQX1 \ram_reg[59][13]  ( .D(n1539), .CK(clk), .Q(\ram[59][13] ) );
  DFFHQX1 \ram_reg[59][12]  ( .D(n1538), .CK(clk), .Q(\ram[59][12] ) );
  DFFHQX1 \ram_reg[59][11]  ( .D(n1537), .CK(clk), .Q(\ram[59][11] ) );
  DFFHQX1 \ram_reg[59][10]  ( .D(n1536), .CK(clk), .Q(\ram[59][10] ) );
  DFFHQX1 \ram_reg[59][9]  ( .D(n1535), .CK(clk), .Q(\ram[59][9] ) );
  DFFHQX1 \ram_reg[59][8]  ( .D(n1534), .CK(clk), .Q(\ram[59][8] ) );
  DFFHQX1 \ram_reg[59][7]  ( .D(n1533), .CK(clk), .Q(\ram[59][7] ) );
  DFFHQX1 \ram_reg[59][6]  ( .D(n1532), .CK(clk), .Q(\ram[59][6] ) );
  DFFHQX1 \ram_reg[59][5]  ( .D(n1531), .CK(clk), .Q(\ram[59][5] ) );
  DFFHQX1 \ram_reg[59][4]  ( .D(n1530), .CK(clk), .Q(\ram[59][4] ) );
  DFFHQX1 \ram_reg[59][3]  ( .D(n1529), .CK(clk), .Q(\ram[59][3] ) );
  DFFHQX1 \ram_reg[59][2]  ( .D(n1528), .CK(clk), .Q(\ram[59][2] ) );
  DFFHQX1 \ram_reg[59][1]  ( .D(n1527), .CK(clk), .Q(\ram[59][1] ) );
  DFFHQX1 \ram_reg[59][0]  ( .D(n1526), .CK(clk), .Q(\ram[59][0] ) );
  DFFHQX1 \ram_reg[55][15]  ( .D(n1477), .CK(clk), .Q(\ram[55][15] ) );
  DFFHQX1 \ram_reg[55][14]  ( .D(n1476), .CK(clk), .Q(\ram[55][14] ) );
  DFFHQX1 \ram_reg[55][13]  ( .D(n1475), .CK(clk), .Q(\ram[55][13] ) );
  DFFHQX1 \ram_reg[55][12]  ( .D(n1474), .CK(clk), .Q(\ram[55][12] ) );
  DFFHQX1 \ram_reg[55][11]  ( .D(n1473), .CK(clk), .Q(\ram[55][11] ) );
  DFFHQX1 \ram_reg[55][10]  ( .D(n1472), .CK(clk), .Q(\ram[55][10] ) );
  DFFHQX1 \ram_reg[55][9]  ( .D(n1471), .CK(clk), .Q(\ram[55][9] ) );
  DFFHQX1 \ram_reg[55][8]  ( .D(n1470), .CK(clk), .Q(\ram[55][8] ) );
  DFFHQX1 \ram_reg[55][7]  ( .D(n1469), .CK(clk), .Q(\ram[55][7] ) );
  DFFHQX1 \ram_reg[55][6]  ( .D(n1468), .CK(clk), .Q(\ram[55][6] ) );
  DFFHQX1 \ram_reg[55][5]  ( .D(n1467), .CK(clk), .Q(\ram[55][5] ) );
  DFFHQX1 \ram_reg[55][4]  ( .D(n1466), .CK(clk), .Q(\ram[55][4] ) );
  DFFHQX1 \ram_reg[55][3]  ( .D(n1465), .CK(clk), .Q(\ram[55][3] ) );
  DFFHQX1 \ram_reg[55][2]  ( .D(n1464), .CK(clk), .Q(\ram[55][2] ) );
  DFFHQX1 \ram_reg[55][1]  ( .D(n1463), .CK(clk), .Q(\ram[55][1] ) );
  DFFHQX1 \ram_reg[55][0]  ( .D(n1462), .CK(clk), .Q(\ram[55][0] ) );
  DFFHQX1 \ram_reg[51][15]  ( .D(n1413), .CK(clk), .Q(\ram[51][15] ) );
  DFFHQX1 \ram_reg[51][14]  ( .D(n1412), .CK(clk), .Q(\ram[51][14] ) );
  DFFHQX1 \ram_reg[51][13]  ( .D(n1411), .CK(clk), .Q(\ram[51][13] ) );
  DFFHQX1 \ram_reg[51][12]  ( .D(n1410), .CK(clk), .Q(\ram[51][12] ) );
  DFFHQX1 \ram_reg[51][11]  ( .D(n1409), .CK(clk), .Q(\ram[51][11] ) );
  DFFHQX1 \ram_reg[51][10]  ( .D(n1408), .CK(clk), .Q(\ram[51][10] ) );
  DFFHQX1 \ram_reg[51][9]  ( .D(n1407), .CK(clk), .Q(\ram[51][9] ) );
  DFFHQX1 \ram_reg[51][8]  ( .D(n1406), .CK(clk), .Q(\ram[51][8] ) );
  DFFHQX1 \ram_reg[51][7]  ( .D(n1405), .CK(clk), .Q(\ram[51][7] ) );
  DFFHQX1 \ram_reg[51][6]  ( .D(n1404), .CK(clk), .Q(\ram[51][6] ) );
  DFFHQX1 \ram_reg[51][5]  ( .D(n1403), .CK(clk), .Q(\ram[51][5] ) );
  DFFHQX1 \ram_reg[51][4]  ( .D(n1402), .CK(clk), .Q(\ram[51][4] ) );
  DFFHQX1 \ram_reg[51][3]  ( .D(n1401), .CK(clk), .Q(\ram[51][3] ) );
  DFFHQX1 \ram_reg[51][2]  ( .D(n1400), .CK(clk), .Q(\ram[51][2] ) );
  DFFHQX1 \ram_reg[51][1]  ( .D(n1399), .CK(clk), .Q(\ram[51][1] ) );
  DFFHQX1 \ram_reg[51][0]  ( .D(n1398), .CK(clk), .Q(\ram[51][0] ) );
  DFFHQX1 \ram_reg[47][15]  ( .D(n1349), .CK(clk), .Q(\ram[47][15] ) );
  DFFHQX1 \ram_reg[47][14]  ( .D(n1348), .CK(clk), .Q(\ram[47][14] ) );
  DFFHQX1 \ram_reg[47][13]  ( .D(n1347), .CK(clk), .Q(\ram[47][13] ) );
  DFFHQX1 \ram_reg[47][12]  ( .D(n1346), .CK(clk), .Q(\ram[47][12] ) );
  DFFHQX1 \ram_reg[47][11]  ( .D(n1345), .CK(clk), .Q(\ram[47][11] ) );
  DFFHQX1 \ram_reg[47][10]  ( .D(n1344), .CK(clk), .Q(\ram[47][10] ) );
  DFFHQX1 \ram_reg[47][9]  ( .D(n1343), .CK(clk), .Q(\ram[47][9] ) );
  DFFHQX1 \ram_reg[47][8]  ( .D(n1342), .CK(clk), .Q(\ram[47][8] ) );
  DFFHQX1 \ram_reg[47][7]  ( .D(n1341), .CK(clk), .Q(\ram[47][7] ) );
  DFFHQX1 \ram_reg[47][6]  ( .D(n1340), .CK(clk), .Q(\ram[47][6] ) );
  DFFHQX1 \ram_reg[47][5]  ( .D(n1339), .CK(clk), .Q(\ram[47][5] ) );
  DFFHQX1 \ram_reg[47][4]  ( .D(n1338), .CK(clk), .Q(\ram[47][4] ) );
  DFFHQX1 \ram_reg[47][3]  ( .D(n1337), .CK(clk), .Q(\ram[47][3] ) );
  DFFHQX1 \ram_reg[47][2]  ( .D(n1336), .CK(clk), .Q(\ram[47][2] ) );
  DFFHQX1 \ram_reg[47][1]  ( .D(n1335), .CK(clk), .Q(\ram[47][1] ) );
  DFFHQX1 \ram_reg[47][0]  ( .D(n1334), .CK(clk), .Q(\ram[47][0] ) );
  DFFHQX1 \ram_reg[43][15]  ( .D(n1285), .CK(clk), .Q(\ram[43][15] ) );
  DFFHQX1 \ram_reg[43][14]  ( .D(n1284), .CK(clk), .Q(\ram[43][14] ) );
  DFFHQX1 \ram_reg[43][13]  ( .D(n1283), .CK(clk), .Q(\ram[43][13] ) );
  DFFHQX1 \ram_reg[43][12]  ( .D(n1282), .CK(clk), .Q(\ram[43][12] ) );
  DFFHQX1 \ram_reg[43][11]  ( .D(n1281), .CK(clk), .Q(\ram[43][11] ) );
  DFFHQX1 \ram_reg[43][10]  ( .D(n1280), .CK(clk), .Q(\ram[43][10] ) );
  DFFHQX1 \ram_reg[43][9]  ( .D(n1279), .CK(clk), .Q(\ram[43][9] ) );
  DFFHQX1 \ram_reg[43][8]  ( .D(n1278), .CK(clk), .Q(\ram[43][8] ) );
  DFFHQX1 \ram_reg[43][7]  ( .D(n1277), .CK(clk), .Q(\ram[43][7] ) );
  DFFHQX1 \ram_reg[43][6]  ( .D(n1276), .CK(clk), .Q(\ram[43][6] ) );
  DFFHQX1 \ram_reg[43][5]  ( .D(n1275), .CK(clk), .Q(\ram[43][5] ) );
  DFFHQX1 \ram_reg[43][4]  ( .D(n1274), .CK(clk), .Q(\ram[43][4] ) );
  DFFHQX1 \ram_reg[43][3]  ( .D(n1273), .CK(clk), .Q(\ram[43][3] ) );
  DFFHQX1 \ram_reg[43][2]  ( .D(n1272), .CK(clk), .Q(\ram[43][2] ) );
  DFFHQX1 \ram_reg[43][1]  ( .D(n1271), .CK(clk), .Q(\ram[43][1] ) );
  DFFHQX1 \ram_reg[43][0]  ( .D(n1270), .CK(clk), .Q(\ram[43][0] ) );
  DFFHQX1 \ram_reg[39][15]  ( .D(n1221), .CK(clk), .Q(\ram[39][15] ) );
  DFFHQX1 \ram_reg[39][14]  ( .D(n1220), .CK(clk), .Q(\ram[39][14] ) );
  DFFHQX1 \ram_reg[39][13]  ( .D(n1219), .CK(clk), .Q(\ram[39][13] ) );
  DFFHQX1 \ram_reg[39][12]  ( .D(n1218), .CK(clk), .Q(\ram[39][12] ) );
  DFFHQX1 \ram_reg[39][11]  ( .D(n1217), .CK(clk), .Q(\ram[39][11] ) );
  DFFHQX1 \ram_reg[39][10]  ( .D(n1216), .CK(clk), .Q(\ram[39][10] ) );
  DFFHQX1 \ram_reg[39][9]  ( .D(n1215), .CK(clk), .Q(\ram[39][9] ) );
  DFFHQX1 \ram_reg[39][8]  ( .D(n1214), .CK(clk), .Q(\ram[39][8] ) );
  DFFHQX1 \ram_reg[39][7]  ( .D(n1213), .CK(clk), .Q(\ram[39][7] ) );
  DFFHQX1 \ram_reg[39][6]  ( .D(n1212), .CK(clk), .Q(\ram[39][6] ) );
  DFFHQX1 \ram_reg[39][5]  ( .D(n1211), .CK(clk), .Q(\ram[39][5] ) );
  DFFHQX1 \ram_reg[39][4]  ( .D(n1210), .CK(clk), .Q(\ram[39][4] ) );
  DFFHQX1 \ram_reg[39][3]  ( .D(n1209), .CK(clk), .Q(\ram[39][3] ) );
  DFFHQX1 \ram_reg[39][2]  ( .D(n1208), .CK(clk), .Q(\ram[39][2] ) );
  DFFHQX1 \ram_reg[39][1]  ( .D(n1207), .CK(clk), .Q(\ram[39][1] ) );
  DFFHQX1 \ram_reg[39][0]  ( .D(n1206), .CK(clk), .Q(\ram[39][0] ) );
  DFFHQX1 \ram_reg[35][15]  ( .D(n1157), .CK(clk), .Q(\ram[35][15] ) );
  DFFHQX1 \ram_reg[35][14]  ( .D(n1156), .CK(clk), .Q(\ram[35][14] ) );
  DFFHQX1 \ram_reg[35][13]  ( .D(n1155), .CK(clk), .Q(\ram[35][13] ) );
  DFFHQX1 \ram_reg[35][12]  ( .D(n1154), .CK(clk), .Q(\ram[35][12] ) );
  DFFHQX1 \ram_reg[35][11]  ( .D(n1153), .CK(clk), .Q(\ram[35][11] ) );
  DFFHQX1 \ram_reg[35][10]  ( .D(n1152), .CK(clk), .Q(\ram[35][10] ) );
  DFFHQX1 \ram_reg[35][9]  ( .D(n1151), .CK(clk), .Q(\ram[35][9] ) );
  DFFHQX1 \ram_reg[35][8]  ( .D(n1150), .CK(clk), .Q(\ram[35][8] ) );
  DFFHQX1 \ram_reg[35][7]  ( .D(n1149), .CK(clk), .Q(\ram[35][7] ) );
  DFFHQX1 \ram_reg[35][6]  ( .D(n1148), .CK(clk), .Q(\ram[35][6] ) );
  DFFHQX1 \ram_reg[35][5]  ( .D(n1147), .CK(clk), .Q(\ram[35][5] ) );
  DFFHQX1 \ram_reg[35][4]  ( .D(n1146), .CK(clk), .Q(\ram[35][4] ) );
  DFFHQX1 \ram_reg[35][3]  ( .D(n1145), .CK(clk), .Q(\ram[35][3] ) );
  DFFHQX1 \ram_reg[35][2]  ( .D(n1144), .CK(clk), .Q(\ram[35][2] ) );
  DFFHQX1 \ram_reg[35][1]  ( .D(n1143), .CK(clk), .Q(\ram[35][1] ) );
  DFFHQX1 \ram_reg[35][0]  ( .D(n1142), .CK(clk), .Q(\ram[35][0] ) );
  DFFHQX1 \ram_reg[31][15]  ( .D(n1093), .CK(clk), .Q(\ram[31][15] ) );
  DFFHQX1 \ram_reg[31][14]  ( .D(n1092), .CK(clk), .Q(\ram[31][14] ) );
  DFFHQX1 \ram_reg[31][13]  ( .D(n1091), .CK(clk), .Q(\ram[31][13] ) );
  DFFHQX1 \ram_reg[31][12]  ( .D(n1090), .CK(clk), .Q(\ram[31][12] ) );
  DFFHQX1 \ram_reg[31][11]  ( .D(n1089), .CK(clk), .Q(\ram[31][11] ) );
  DFFHQX1 \ram_reg[31][10]  ( .D(n1088), .CK(clk), .Q(\ram[31][10] ) );
  DFFHQX1 \ram_reg[31][9]  ( .D(n1087), .CK(clk), .Q(\ram[31][9] ) );
  DFFHQX1 \ram_reg[31][8]  ( .D(n1086), .CK(clk), .Q(\ram[31][8] ) );
  DFFHQX1 \ram_reg[31][7]  ( .D(n1085), .CK(clk), .Q(\ram[31][7] ) );
  DFFHQX1 \ram_reg[31][6]  ( .D(n1084), .CK(clk), .Q(\ram[31][6] ) );
  DFFHQX1 \ram_reg[31][5]  ( .D(n1083), .CK(clk), .Q(\ram[31][5] ) );
  DFFHQX1 \ram_reg[31][4]  ( .D(n1082), .CK(clk), .Q(\ram[31][4] ) );
  DFFHQX1 \ram_reg[31][3]  ( .D(n1081), .CK(clk), .Q(\ram[31][3] ) );
  DFFHQX1 \ram_reg[31][2]  ( .D(n1080), .CK(clk), .Q(\ram[31][2] ) );
  DFFHQX1 \ram_reg[31][1]  ( .D(n1079), .CK(clk), .Q(\ram[31][1] ) );
  DFFHQX1 \ram_reg[31][0]  ( .D(n1078), .CK(clk), .Q(\ram[31][0] ) );
  DFFHQX1 \ram_reg[27][15]  ( .D(n1029), .CK(clk), .Q(\ram[27][15] ) );
  DFFHQX1 \ram_reg[27][14]  ( .D(n1028), .CK(clk), .Q(\ram[27][14] ) );
  DFFHQX1 \ram_reg[27][13]  ( .D(n1027), .CK(clk), .Q(\ram[27][13] ) );
  DFFHQX1 \ram_reg[27][12]  ( .D(n1026), .CK(clk), .Q(\ram[27][12] ) );
  DFFHQX1 \ram_reg[27][11]  ( .D(n1025), .CK(clk), .Q(\ram[27][11] ) );
  DFFHQX1 \ram_reg[27][10]  ( .D(n1024), .CK(clk), .Q(\ram[27][10] ) );
  DFFHQX1 \ram_reg[27][9]  ( .D(n1023), .CK(clk), .Q(\ram[27][9] ) );
  DFFHQX1 \ram_reg[27][8]  ( .D(n1022), .CK(clk), .Q(\ram[27][8] ) );
  DFFHQX1 \ram_reg[27][7]  ( .D(n1021), .CK(clk), .Q(\ram[27][7] ) );
  DFFHQX1 \ram_reg[27][6]  ( .D(n1020), .CK(clk), .Q(\ram[27][6] ) );
  DFFHQX1 \ram_reg[27][5]  ( .D(n1019), .CK(clk), .Q(\ram[27][5] ) );
  DFFHQX1 \ram_reg[27][4]  ( .D(n1018), .CK(clk), .Q(\ram[27][4] ) );
  DFFHQX1 \ram_reg[27][3]  ( .D(n1017), .CK(clk), .Q(\ram[27][3] ) );
  DFFHQX1 \ram_reg[27][2]  ( .D(n1016), .CK(clk), .Q(\ram[27][2] ) );
  DFFHQX1 \ram_reg[27][1]  ( .D(n1015), .CK(clk), .Q(\ram[27][1] ) );
  DFFHQX1 \ram_reg[27][0]  ( .D(n1014), .CK(clk), .Q(\ram[27][0] ) );
  DFFHQX1 \ram_reg[23][15]  ( .D(n965), .CK(clk), .Q(\ram[23][15] ) );
  DFFHQX1 \ram_reg[23][14]  ( .D(n964), .CK(clk), .Q(\ram[23][14] ) );
  DFFHQX1 \ram_reg[23][13]  ( .D(n963), .CK(clk), .Q(\ram[23][13] ) );
  DFFHQX1 \ram_reg[23][12]  ( .D(n962), .CK(clk), .Q(\ram[23][12] ) );
  DFFHQX1 \ram_reg[23][11]  ( .D(n961), .CK(clk), .Q(\ram[23][11] ) );
  DFFHQX1 \ram_reg[23][10]  ( .D(n960), .CK(clk), .Q(\ram[23][10] ) );
  DFFHQX1 \ram_reg[23][9]  ( .D(n959), .CK(clk), .Q(\ram[23][9] ) );
  DFFHQX1 \ram_reg[23][8]  ( .D(n958), .CK(clk), .Q(\ram[23][8] ) );
  DFFHQX1 \ram_reg[23][7]  ( .D(n957), .CK(clk), .Q(\ram[23][7] ) );
  DFFHQX1 \ram_reg[23][6]  ( .D(n956), .CK(clk), .Q(\ram[23][6] ) );
  DFFHQX1 \ram_reg[23][5]  ( .D(n955), .CK(clk), .Q(\ram[23][5] ) );
  DFFHQX1 \ram_reg[23][4]  ( .D(n954), .CK(clk), .Q(\ram[23][4] ) );
  DFFHQX1 \ram_reg[23][3]  ( .D(n953), .CK(clk), .Q(\ram[23][3] ) );
  DFFHQX1 \ram_reg[23][2]  ( .D(n952), .CK(clk), .Q(\ram[23][2] ) );
  DFFHQX1 \ram_reg[23][1]  ( .D(n951), .CK(clk), .Q(\ram[23][1] ) );
  DFFHQX1 \ram_reg[23][0]  ( .D(n950), .CK(clk), .Q(\ram[23][0] ) );
  DFFHQX1 \ram_reg[19][15]  ( .D(n901), .CK(clk), .Q(\ram[19][15] ) );
  DFFHQX1 \ram_reg[19][14]  ( .D(n900), .CK(clk), .Q(\ram[19][14] ) );
  DFFHQX1 \ram_reg[19][13]  ( .D(n899), .CK(clk), .Q(\ram[19][13] ) );
  DFFHQX1 \ram_reg[19][12]  ( .D(n898), .CK(clk), .Q(\ram[19][12] ) );
  DFFHQX1 \ram_reg[19][11]  ( .D(n897), .CK(clk), .Q(\ram[19][11] ) );
  DFFHQX1 \ram_reg[19][10]  ( .D(n896), .CK(clk), .Q(\ram[19][10] ) );
  DFFHQX1 \ram_reg[19][9]  ( .D(n895), .CK(clk), .Q(\ram[19][9] ) );
  DFFHQX1 \ram_reg[19][8]  ( .D(n894), .CK(clk), .Q(\ram[19][8] ) );
  DFFHQX1 \ram_reg[19][7]  ( .D(n893), .CK(clk), .Q(\ram[19][7] ) );
  DFFHQX1 \ram_reg[19][6]  ( .D(n892), .CK(clk), .Q(\ram[19][6] ) );
  DFFHQX1 \ram_reg[19][5]  ( .D(n891), .CK(clk), .Q(\ram[19][5] ) );
  DFFHQX1 \ram_reg[19][4]  ( .D(n890), .CK(clk), .Q(\ram[19][4] ) );
  DFFHQX1 \ram_reg[19][3]  ( .D(n889), .CK(clk), .Q(\ram[19][3] ) );
  DFFHQX1 \ram_reg[19][2]  ( .D(n888), .CK(clk), .Q(\ram[19][2] ) );
  DFFHQX1 \ram_reg[19][1]  ( .D(n887), .CK(clk), .Q(\ram[19][1] ) );
  DFFHQX1 \ram_reg[19][0]  ( .D(n886), .CK(clk), .Q(\ram[19][0] ) );
  DFFHQX1 \ram_reg[15][15]  ( .D(n837), .CK(clk), .Q(\ram[15][15] ) );
  DFFHQX1 \ram_reg[15][14]  ( .D(n836), .CK(clk), .Q(\ram[15][14] ) );
  DFFHQX1 \ram_reg[15][13]  ( .D(n835), .CK(clk), .Q(\ram[15][13] ) );
  DFFHQX1 \ram_reg[15][12]  ( .D(n834), .CK(clk), .Q(\ram[15][12] ) );
  DFFHQX1 \ram_reg[15][11]  ( .D(n833), .CK(clk), .Q(\ram[15][11] ) );
  DFFHQX1 \ram_reg[15][10]  ( .D(n832), .CK(clk), .Q(\ram[15][10] ) );
  DFFHQX1 \ram_reg[15][9]  ( .D(n831), .CK(clk), .Q(\ram[15][9] ) );
  DFFHQX1 \ram_reg[15][8]  ( .D(n830), .CK(clk), .Q(\ram[15][8] ) );
  DFFHQX1 \ram_reg[15][7]  ( .D(n829), .CK(clk), .Q(\ram[15][7] ) );
  DFFHQX1 \ram_reg[15][6]  ( .D(n828), .CK(clk), .Q(\ram[15][6] ) );
  DFFHQX1 \ram_reg[15][5]  ( .D(n827), .CK(clk), .Q(\ram[15][5] ) );
  DFFHQX1 \ram_reg[15][4]  ( .D(n826), .CK(clk), .Q(\ram[15][4] ) );
  DFFHQX1 \ram_reg[15][3]  ( .D(n825), .CK(clk), .Q(\ram[15][3] ) );
  DFFHQX1 \ram_reg[15][2]  ( .D(n824), .CK(clk), .Q(\ram[15][2] ) );
  DFFHQX1 \ram_reg[15][1]  ( .D(n823), .CK(clk), .Q(\ram[15][1] ) );
  DFFHQX1 \ram_reg[15][0]  ( .D(n822), .CK(clk), .Q(\ram[15][0] ) );
  DFFHQX1 \ram_reg[11][15]  ( .D(n773), .CK(clk), .Q(\ram[11][15] ) );
  DFFHQX1 \ram_reg[11][14]  ( .D(n772), .CK(clk), .Q(\ram[11][14] ) );
  DFFHQX1 \ram_reg[11][13]  ( .D(n771), .CK(clk), .Q(\ram[11][13] ) );
  DFFHQX1 \ram_reg[11][12]  ( .D(n770), .CK(clk), .Q(\ram[11][12] ) );
  DFFHQX1 \ram_reg[11][11]  ( .D(n769), .CK(clk), .Q(\ram[11][11] ) );
  DFFHQX1 \ram_reg[11][10]  ( .D(n768), .CK(clk), .Q(\ram[11][10] ) );
  DFFHQX1 \ram_reg[11][9]  ( .D(n767), .CK(clk), .Q(\ram[11][9] ) );
  DFFHQX1 \ram_reg[11][8]  ( .D(n766), .CK(clk), .Q(\ram[11][8] ) );
  DFFHQX1 \ram_reg[11][7]  ( .D(n765), .CK(clk), .Q(\ram[11][7] ) );
  DFFHQX1 \ram_reg[11][6]  ( .D(n764), .CK(clk), .Q(\ram[11][6] ) );
  DFFHQX1 \ram_reg[11][5]  ( .D(n763), .CK(clk), .Q(\ram[11][5] ) );
  DFFHQX1 \ram_reg[11][4]  ( .D(n762), .CK(clk), .Q(\ram[11][4] ) );
  DFFHQX1 \ram_reg[11][3]  ( .D(n761), .CK(clk), .Q(\ram[11][3] ) );
  DFFHQX1 \ram_reg[11][2]  ( .D(n760), .CK(clk), .Q(\ram[11][2] ) );
  DFFHQX1 \ram_reg[11][1]  ( .D(n759), .CK(clk), .Q(\ram[11][1] ) );
  DFFHQX1 \ram_reg[11][0]  ( .D(n758), .CK(clk), .Q(\ram[11][0] ) );
  DFFHQX1 \ram_reg[7][15]  ( .D(n709), .CK(clk), .Q(\ram[7][15] ) );
  DFFHQX1 \ram_reg[7][14]  ( .D(n708), .CK(clk), .Q(\ram[7][14] ) );
  DFFHQX1 \ram_reg[7][13]  ( .D(n707), .CK(clk), .Q(\ram[7][13] ) );
  DFFHQX1 \ram_reg[7][12]  ( .D(n706), .CK(clk), .Q(\ram[7][12] ) );
  DFFHQX1 \ram_reg[7][11]  ( .D(n705), .CK(clk), .Q(\ram[7][11] ) );
  DFFHQX1 \ram_reg[7][10]  ( .D(n704), .CK(clk), .Q(\ram[7][10] ) );
  DFFHQX1 \ram_reg[7][9]  ( .D(n703), .CK(clk), .Q(\ram[7][9] ) );
  DFFHQX1 \ram_reg[7][8]  ( .D(n702), .CK(clk), .Q(\ram[7][8] ) );
  DFFHQX1 \ram_reg[7][7]  ( .D(n701), .CK(clk), .Q(\ram[7][7] ) );
  DFFHQX1 \ram_reg[7][6]  ( .D(n700), .CK(clk), .Q(\ram[7][6] ) );
  DFFHQX1 \ram_reg[7][5]  ( .D(n699), .CK(clk), .Q(\ram[7][5] ) );
  DFFHQX1 \ram_reg[7][4]  ( .D(n698), .CK(clk), .Q(\ram[7][4] ) );
  DFFHQX1 \ram_reg[7][3]  ( .D(n697), .CK(clk), .Q(\ram[7][3] ) );
  DFFHQX1 \ram_reg[7][2]  ( .D(n696), .CK(clk), .Q(\ram[7][2] ) );
  DFFHQX1 \ram_reg[7][1]  ( .D(n695), .CK(clk), .Q(\ram[7][1] ) );
  DFFHQX1 \ram_reg[7][0]  ( .D(n694), .CK(clk), .Q(\ram[7][0] ) );
  DFFHQX1 \ram_reg[3][15]  ( .D(n645), .CK(clk), .Q(\ram[3][15] ) );
  DFFHQX1 \ram_reg[3][14]  ( .D(n644), .CK(clk), .Q(\ram[3][14] ) );
  DFFHQX1 \ram_reg[3][13]  ( .D(n643), .CK(clk), .Q(\ram[3][13] ) );
  DFFHQX1 \ram_reg[3][12]  ( .D(n642), .CK(clk), .Q(\ram[3][12] ) );
  DFFHQX1 \ram_reg[3][11]  ( .D(n641), .CK(clk), .Q(\ram[3][11] ) );
  DFFHQX1 \ram_reg[3][10]  ( .D(n640), .CK(clk), .Q(\ram[3][10] ) );
  DFFHQX1 \ram_reg[3][9]  ( .D(n639), .CK(clk), .Q(\ram[3][9] ) );
  DFFHQX1 \ram_reg[3][8]  ( .D(n638), .CK(clk), .Q(\ram[3][8] ) );
  DFFHQX1 \ram_reg[3][7]  ( .D(n637), .CK(clk), .Q(\ram[3][7] ) );
  DFFHQX1 \ram_reg[3][6]  ( .D(n636), .CK(clk), .Q(\ram[3][6] ) );
  DFFHQX1 \ram_reg[3][5]  ( .D(n635), .CK(clk), .Q(\ram[3][5] ) );
  DFFHQX1 \ram_reg[3][4]  ( .D(n634), .CK(clk), .Q(\ram[3][4] ) );
  DFFHQX1 \ram_reg[3][3]  ( .D(n633), .CK(clk), .Q(\ram[3][3] ) );
  DFFHQX1 \ram_reg[3][2]  ( .D(n632), .CK(clk), .Q(\ram[3][2] ) );
  DFFHQX1 \ram_reg[3][1]  ( .D(n631), .CK(clk), .Q(\ram[3][1] ) );
  DFFHQX1 \ram_reg[3][0]  ( .D(n630), .CK(clk), .Q(\ram[3][0] ) );
  DFFHQX1 \ram_reg[252][15]  ( .D(n4629), .CK(clk), .Q(\ram[252][15] ) );
  DFFHQX1 \ram_reg[252][14]  ( .D(n4628), .CK(clk), .Q(\ram[252][14] ) );
  DFFHQX1 \ram_reg[252][13]  ( .D(n4627), .CK(clk), .Q(\ram[252][13] ) );
  DFFHQX1 \ram_reg[252][12]  ( .D(n4626), .CK(clk), .Q(\ram[252][12] ) );
  DFFHQX1 \ram_reg[252][11]  ( .D(n4625), .CK(clk), .Q(\ram[252][11] ) );
  DFFHQX1 \ram_reg[252][10]  ( .D(n4624), .CK(clk), .Q(\ram[252][10] ) );
  DFFHQX1 \ram_reg[252][9]  ( .D(n4623), .CK(clk), .Q(\ram[252][9] ) );
  DFFHQX1 \ram_reg[252][8]  ( .D(n4622), .CK(clk), .Q(\ram[252][8] ) );
  DFFHQX1 \ram_reg[252][7]  ( .D(n4621), .CK(clk), .Q(\ram[252][7] ) );
  DFFHQX1 \ram_reg[252][6]  ( .D(n4620), .CK(clk), .Q(\ram[252][6] ) );
  DFFHQX1 \ram_reg[252][5]  ( .D(n4619), .CK(clk), .Q(\ram[252][5] ) );
  DFFHQX1 \ram_reg[252][4]  ( .D(n4618), .CK(clk), .Q(\ram[252][4] ) );
  DFFHQX1 \ram_reg[252][3]  ( .D(n4617), .CK(clk), .Q(\ram[252][3] ) );
  DFFHQX1 \ram_reg[252][2]  ( .D(n4616), .CK(clk), .Q(\ram[252][2] ) );
  DFFHQX1 \ram_reg[252][1]  ( .D(n4615), .CK(clk), .Q(\ram[252][1] ) );
  DFFHQX1 \ram_reg[252][0]  ( .D(n4614), .CK(clk), .Q(\ram[252][0] ) );
  DFFHQX1 \ram_reg[248][15]  ( .D(n4565), .CK(clk), .Q(\ram[248][15] ) );
  DFFHQX1 \ram_reg[248][14]  ( .D(n4564), .CK(clk), .Q(\ram[248][14] ) );
  DFFHQX1 \ram_reg[248][13]  ( .D(n4563), .CK(clk), .Q(\ram[248][13] ) );
  DFFHQX1 \ram_reg[248][12]  ( .D(n4562), .CK(clk), .Q(\ram[248][12] ) );
  DFFHQX1 \ram_reg[248][11]  ( .D(n4561), .CK(clk), .Q(\ram[248][11] ) );
  DFFHQX1 \ram_reg[248][10]  ( .D(n4560), .CK(clk), .Q(\ram[248][10] ) );
  DFFHQX1 \ram_reg[248][9]  ( .D(n4559), .CK(clk), .Q(\ram[248][9] ) );
  DFFHQX1 \ram_reg[248][8]  ( .D(n4558), .CK(clk), .Q(\ram[248][8] ) );
  DFFHQX1 \ram_reg[248][7]  ( .D(n4557), .CK(clk), .Q(\ram[248][7] ) );
  DFFHQX1 \ram_reg[248][6]  ( .D(n4556), .CK(clk), .Q(\ram[248][6] ) );
  DFFHQX1 \ram_reg[248][5]  ( .D(n4555), .CK(clk), .Q(\ram[248][5] ) );
  DFFHQX1 \ram_reg[248][4]  ( .D(n4554), .CK(clk), .Q(\ram[248][4] ) );
  DFFHQX1 \ram_reg[248][3]  ( .D(n4553), .CK(clk), .Q(\ram[248][3] ) );
  DFFHQX1 \ram_reg[248][2]  ( .D(n4552), .CK(clk), .Q(\ram[248][2] ) );
  DFFHQX1 \ram_reg[248][1]  ( .D(n4551), .CK(clk), .Q(\ram[248][1] ) );
  DFFHQX1 \ram_reg[248][0]  ( .D(n4550), .CK(clk), .Q(\ram[248][0] ) );
  DFFHQX1 \ram_reg[244][15]  ( .D(n4501), .CK(clk), .Q(\ram[244][15] ) );
  DFFHQX1 \ram_reg[244][14]  ( .D(n4500), .CK(clk), .Q(\ram[244][14] ) );
  DFFHQX1 \ram_reg[244][13]  ( .D(n4499), .CK(clk), .Q(\ram[244][13] ) );
  DFFHQX1 \ram_reg[244][12]  ( .D(n4498), .CK(clk), .Q(\ram[244][12] ) );
  DFFHQX1 \ram_reg[244][11]  ( .D(n4497), .CK(clk), .Q(\ram[244][11] ) );
  DFFHQX1 \ram_reg[244][10]  ( .D(n4496), .CK(clk), .Q(\ram[244][10] ) );
  DFFHQX1 \ram_reg[244][9]  ( .D(n4495), .CK(clk), .Q(\ram[244][9] ) );
  DFFHQX1 \ram_reg[244][8]  ( .D(n4494), .CK(clk), .Q(\ram[244][8] ) );
  DFFHQX1 \ram_reg[244][7]  ( .D(n4493), .CK(clk), .Q(\ram[244][7] ) );
  DFFHQX1 \ram_reg[244][6]  ( .D(n4492), .CK(clk), .Q(\ram[244][6] ) );
  DFFHQX1 \ram_reg[244][5]  ( .D(n4491), .CK(clk), .Q(\ram[244][5] ) );
  DFFHQX1 \ram_reg[244][4]  ( .D(n4490), .CK(clk), .Q(\ram[244][4] ) );
  DFFHQX1 \ram_reg[244][3]  ( .D(n4489), .CK(clk), .Q(\ram[244][3] ) );
  DFFHQX1 \ram_reg[244][2]  ( .D(n4488), .CK(clk), .Q(\ram[244][2] ) );
  DFFHQX1 \ram_reg[244][1]  ( .D(n4487), .CK(clk), .Q(\ram[244][1] ) );
  DFFHQX1 \ram_reg[244][0]  ( .D(n4486), .CK(clk), .Q(\ram[244][0] ) );
  DFFHQX1 \ram_reg[240][15]  ( .D(n4437), .CK(clk), .Q(\ram[240][15] ) );
  DFFHQX1 \ram_reg[240][14]  ( .D(n4436), .CK(clk), .Q(\ram[240][14] ) );
  DFFHQX1 \ram_reg[240][13]  ( .D(n4435), .CK(clk), .Q(\ram[240][13] ) );
  DFFHQX1 \ram_reg[240][12]  ( .D(n4434), .CK(clk), .Q(\ram[240][12] ) );
  DFFHQX1 \ram_reg[240][11]  ( .D(n4433), .CK(clk), .Q(\ram[240][11] ) );
  DFFHQX1 \ram_reg[240][10]  ( .D(n4432), .CK(clk), .Q(\ram[240][10] ) );
  DFFHQX1 \ram_reg[240][9]  ( .D(n4431), .CK(clk), .Q(\ram[240][9] ) );
  DFFHQX1 \ram_reg[240][8]  ( .D(n4430), .CK(clk), .Q(\ram[240][8] ) );
  DFFHQX1 \ram_reg[240][7]  ( .D(n4429), .CK(clk), .Q(\ram[240][7] ) );
  DFFHQX1 \ram_reg[240][6]  ( .D(n4428), .CK(clk), .Q(\ram[240][6] ) );
  DFFHQX1 \ram_reg[240][5]  ( .D(n4427), .CK(clk), .Q(\ram[240][5] ) );
  DFFHQX1 \ram_reg[240][4]  ( .D(n4426), .CK(clk), .Q(\ram[240][4] ) );
  DFFHQX1 \ram_reg[240][3]  ( .D(n4425), .CK(clk), .Q(\ram[240][3] ) );
  DFFHQX1 \ram_reg[240][2]  ( .D(n4424), .CK(clk), .Q(\ram[240][2] ) );
  DFFHQX1 \ram_reg[240][1]  ( .D(n4423), .CK(clk), .Q(\ram[240][1] ) );
  DFFHQX1 \ram_reg[240][0]  ( .D(n4422), .CK(clk), .Q(\ram[240][0] ) );
  DFFHQX1 \ram_reg[236][15]  ( .D(n4373), .CK(clk), .Q(\ram[236][15] ) );
  DFFHQX1 \ram_reg[236][14]  ( .D(n4372), .CK(clk), .Q(\ram[236][14] ) );
  DFFHQX1 \ram_reg[236][13]  ( .D(n4371), .CK(clk), .Q(\ram[236][13] ) );
  DFFHQX1 \ram_reg[236][12]  ( .D(n4370), .CK(clk), .Q(\ram[236][12] ) );
  DFFHQX1 \ram_reg[236][11]  ( .D(n4369), .CK(clk), .Q(\ram[236][11] ) );
  DFFHQX1 \ram_reg[236][10]  ( .D(n4368), .CK(clk), .Q(\ram[236][10] ) );
  DFFHQX1 \ram_reg[236][9]  ( .D(n4367), .CK(clk), .Q(\ram[236][9] ) );
  DFFHQX1 \ram_reg[236][8]  ( .D(n4366), .CK(clk), .Q(\ram[236][8] ) );
  DFFHQX1 \ram_reg[236][7]  ( .D(n4365), .CK(clk), .Q(\ram[236][7] ) );
  DFFHQX1 \ram_reg[236][6]  ( .D(n4364), .CK(clk), .Q(\ram[236][6] ) );
  DFFHQX1 \ram_reg[236][5]  ( .D(n4363), .CK(clk), .Q(\ram[236][5] ) );
  DFFHQX1 \ram_reg[236][4]  ( .D(n4362), .CK(clk), .Q(\ram[236][4] ) );
  DFFHQX1 \ram_reg[236][3]  ( .D(n4361), .CK(clk), .Q(\ram[236][3] ) );
  DFFHQX1 \ram_reg[236][2]  ( .D(n4360), .CK(clk), .Q(\ram[236][2] ) );
  DFFHQX1 \ram_reg[236][1]  ( .D(n4359), .CK(clk), .Q(\ram[236][1] ) );
  DFFHQX1 \ram_reg[236][0]  ( .D(n4358), .CK(clk), .Q(\ram[236][0] ) );
  DFFHQX1 \ram_reg[232][15]  ( .D(n4309), .CK(clk), .Q(\ram[232][15] ) );
  DFFHQX1 \ram_reg[232][14]  ( .D(n4308), .CK(clk), .Q(\ram[232][14] ) );
  DFFHQX1 \ram_reg[232][13]  ( .D(n4307), .CK(clk), .Q(\ram[232][13] ) );
  DFFHQX1 \ram_reg[232][12]  ( .D(n4306), .CK(clk), .Q(\ram[232][12] ) );
  DFFHQX1 \ram_reg[232][11]  ( .D(n4305), .CK(clk), .Q(\ram[232][11] ) );
  DFFHQX1 \ram_reg[232][10]  ( .D(n4304), .CK(clk), .Q(\ram[232][10] ) );
  DFFHQX1 \ram_reg[232][9]  ( .D(n4303), .CK(clk), .Q(\ram[232][9] ) );
  DFFHQX1 \ram_reg[232][8]  ( .D(n4302), .CK(clk), .Q(\ram[232][8] ) );
  DFFHQX1 \ram_reg[232][7]  ( .D(n4301), .CK(clk), .Q(\ram[232][7] ) );
  DFFHQX1 \ram_reg[232][6]  ( .D(n4300), .CK(clk), .Q(\ram[232][6] ) );
  DFFHQX1 \ram_reg[232][5]  ( .D(n4299), .CK(clk), .Q(\ram[232][5] ) );
  DFFHQX1 \ram_reg[232][4]  ( .D(n4298), .CK(clk), .Q(\ram[232][4] ) );
  DFFHQX1 \ram_reg[232][3]  ( .D(n4297), .CK(clk), .Q(\ram[232][3] ) );
  DFFHQX1 \ram_reg[232][2]  ( .D(n4296), .CK(clk), .Q(\ram[232][2] ) );
  DFFHQX1 \ram_reg[232][1]  ( .D(n4295), .CK(clk), .Q(\ram[232][1] ) );
  DFFHQX1 \ram_reg[232][0]  ( .D(n4294), .CK(clk), .Q(\ram[232][0] ) );
  DFFHQX1 \ram_reg[228][15]  ( .D(n4245), .CK(clk), .Q(\ram[228][15] ) );
  DFFHQX1 \ram_reg[228][14]  ( .D(n4244), .CK(clk), .Q(\ram[228][14] ) );
  DFFHQX1 \ram_reg[228][13]  ( .D(n4243), .CK(clk), .Q(\ram[228][13] ) );
  DFFHQX1 \ram_reg[228][12]  ( .D(n4242), .CK(clk), .Q(\ram[228][12] ) );
  DFFHQX1 \ram_reg[228][11]  ( .D(n4241), .CK(clk), .Q(\ram[228][11] ) );
  DFFHQX1 \ram_reg[228][10]  ( .D(n4240), .CK(clk), .Q(\ram[228][10] ) );
  DFFHQX1 \ram_reg[228][9]  ( .D(n4239), .CK(clk), .Q(\ram[228][9] ) );
  DFFHQX1 \ram_reg[228][8]  ( .D(n4238), .CK(clk), .Q(\ram[228][8] ) );
  DFFHQX1 \ram_reg[228][7]  ( .D(n4237), .CK(clk), .Q(\ram[228][7] ) );
  DFFHQX1 \ram_reg[228][6]  ( .D(n4236), .CK(clk), .Q(\ram[228][6] ) );
  DFFHQX1 \ram_reg[228][5]  ( .D(n4235), .CK(clk), .Q(\ram[228][5] ) );
  DFFHQX1 \ram_reg[228][4]  ( .D(n4234), .CK(clk), .Q(\ram[228][4] ) );
  DFFHQX1 \ram_reg[228][3]  ( .D(n4233), .CK(clk), .Q(\ram[228][3] ) );
  DFFHQX1 \ram_reg[228][2]  ( .D(n4232), .CK(clk), .Q(\ram[228][2] ) );
  DFFHQX1 \ram_reg[228][1]  ( .D(n4231), .CK(clk), .Q(\ram[228][1] ) );
  DFFHQX1 \ram_reg[228][0]  ( .D(n4230), .CK(clk), .Q(\ram[228][0] ) );
  DFFHQX1 \ram_reg[224][15]  ( .D(n4181), .CK(clk), .Q(\ram[224][15] ) );
  DFFHQX1 \ram_reg[224][14]  ( .D(n4180), .CK(clk), .Q(\ram[224][14] ) );
  DFFHQX1 \ram_reg[224][13]  ( .D(n4179), .CK(clk), .Q(\ram[224][13] ) );
  DFFHQX1 \ram_reg[224][12]  ( .D(n4178), .CK(clk), .Q(\ram[224][12] ) );
  DFFHQX1 \ram_reg[224][11]  ( .D(n4177), .CK(clk), .Q(\ram[224][11] ) );
  DFFHQX1 \ram_reg[224][10]  ( .D(n4176), .CK(clk), .Q(\ram[224][10] ) );
  DFFHQX1 \ram_reg[224][9]  ( .D(n4175), .CK(clk), .Q(\ram[224][9] ) );
  DFFHQX1 \ram_reg[224][8]  ( .D(n4174), .CK(clk), .Q(\ram[224][8] ) );
  DFFHQX1 \ram_reg[224][7]  ( .D(n4173), .CK(clk), .Q(\ram[224][7] ) );
  DFFHQX1 \ram_reg[224][6]  ( .D(n4172), .CK(clk), .Q(\ram[224][6] ) );
  DFFHQX1 \ram_reg[224][5]  ( .D(n4171), .CK(clk), .Q(\ram[224][5] ) );
  DFFHQX1 \ram_reg[224][4]  ( .D(n4170), .CK(clk), .Q(\ram[224][4] ) );
  DFFHQX1 \ram_reg[224][3]  ( .D(n4169), .CK(clk), .Q(\ram[224][3] ) );
  DFFHQX1 \ram_reg[224][2]  ( .D(n4168), .CK(clk), .Q(\ram[224][2] ) );
  DFFHQX1 \ram_reg[224][1]  ( .D(n4167), .CK(clk), .Q(\ram[224][1] ) );
  DFFHQX1 \ram_reg[224][0]  ( .D(n4166), .CK(clk), .Q(\ram[224][0] ) );
  DFFHQX1 \ram_reg[220][15]  ( .D(n4117), .CK(clk), .Q(\ram[220][15] ) );
  DFFHQX1 \ram_reg[220][14]  ( .D(n4116), .CK(clk), .Q(\ram[220][14] ) );
  DFFHQX1 \ram_reg[220][13]  ( .D(n4115), .CK(clk), .Q(\ram[220][13] ) );
  DFFHQX1 \ram_reg[220][12]  ( .D(n4114), .CK(clk), .Q(\ram[220][12] ) );
  DFFHQX1 \ram_reg[220][11]  ( .D(n4113), .CK(clk), .Q(\ram[220][11] ) );
  DFFHQX1 \ram_reg[220][10]  ( .D(n4112), .CK(clk), .Q(\ram[220][10] ) );
  DFFHQX1 \ram_reg[220][9]  ( .D(n4111), .CK(clk), .Q(\ram[220][9] ) );
  DFFHQX1 \ram_reg[220][8]  ( .D(n4110), .CK(clk), .Q(\ram[220][8] ) );
  DFFHQX1 \ram_reg[220][7]  ( .D(n4109), .CK(clk), .Q(\ram[220][7] ) );
  DFFHQX1 \ram_reg[220][6]  ( .D(n4108), .CK(clk), .Q(\ram[220][6] ) );
  DFFHQX1 \ram_reg[220][5]  ( .D(n4107), .CK(clk), .Q(\ram[220][5] ) );
  DFFHQX1 \ram_reg[220][4]  ( .D(n4106), .CK(clk), .Q(\ram[220][4] ) );
  DFFHQX1 \ram_reg[220][3]  ( .D(n4105), .CK(clk), .Q(\ram[220][3] ) );
  DFFHQX1 \ram_reg[220][2]  ( .D(n4104), .CK(clk), .Q(\ram[220][2] ) );
  DFFHQX1 \ram_reg[220][1]  ( .D(n4103), .CK(clk), .Q(\ram[220][1] ) );
  DFFHQX1 \ram_reg[220][0]  ( .D(n4102), .CK(clk), .Q(\ram[220][0] ) );
  DFFHQX1 \ram_reg[216][15]  ( .D(n4053), .CK(clk), .Q(\ram[216][15] ) );
  DFFHQX1 \ram_reg[216][14]  ( .D(n4052), .CK(clk), .Q(\ram[216][14] ) );
  DFFHQX1 \ram_reg[216][13]  ( .D(n4051), .CK(clk), .Q(\ram[216][13] ) );
  DFFHQX1 \ram_reg[216][12]  ( .D(n4050), .CK(clk), .Q(\ram[216][12] ) );
  DFFHQX1 \ram_reg[216][11]  ( .D(n4049), .CK(clk), .Q(\ram[216][11] ) );
  DFFHQX1 \ram_reg[216][10]  ( .D(n4048), .CK(clk), .Q(\ram[216][10] ) );
  DFFHQX1 \ram_reg[216][9]  ( .D(n4047), .CK(clk), .Q(\ram[216][9] ) );
  DFFHQX1 \ram_reg[216][8]  ( .D(n4046), .CK(clk), .Q(\ram[216][8] ) );
  DFFHQX1 \ram_reg[216][7]  ( .D(n4045), .CK(clk), .Q(\ram[216][7] ) );
  DFFHQX1 \ram_reg[216][6]  ( .D(n4044), .CK(clk), .Q(\ram[216][6] ) );
  DFFHQX1 \ram_reg[216][5]  ( .D(n4043), .CK(clk), .Q(\ram[216][5] ) );
  DFFHQX1 \ram_reg[216][4]  ( .D(n4042), .CK(clk), .Q(\ram[216][4] ) );
  DFFHQX1 \ram_reg[216][3]  ( .D(n4041), .CK(clk), .Q(\ram[216][3] ) );
  DFFHQX1 \ram_reg[216][2]  ( .D(n4040), .CK(clk), .Q(\ram[216][2] ) );
  DFFHQX1 \ram_reg[216][1]  ( .D(n4039), .CK(clk), .Q(\ram[216][1] ) );
  DFFHQX1 \ram_reg[216][0]  ( .D(n4038), .CK(clk), .Q(\ram[216][0] ) );
  DFFHQX1 \ram_reg[212][15]  ( .D(n3989), .CK(clk), .Q(\ram[212][15] ) );
  DFFHQX1 \ram_reg[212][14]  ( .D(n3988), .CK(clk), .Q(\ram[212][14] ) );
  DFFHQX1 \ram_reg[212][13]  ( .D(n3987), .CK(clk), .Q(\ram[212][13] ) );
  DFFHQX1 \ram_reg[212][12]  ( .D(n3986), .CK(clk), .Q(\ram[212][12] ) );
  DFFHQX1 \ram_reg[212][11]  ( .D(n3985), .CK(clk), .Q(\ram[212][11] ) );
  DFFHQX1 \ram_reg[212][10]  ( .D(n3984), .CK(clk), .Q(\ram[212][10] ) );
  DFFHQX1 \ram_reg[212][9]  ( .D(n3983), .CK(clk), .Q(\ram[212][9] ) );
  DFFHQX1 \ram_reg[212][8]  ( .D(n3982), .CK(clk), .Q(\ram[212][8] ) );
  DFFHQX1 \ram_reg[212][7]  ( .D(n3981), .CK(clk), .Q(\ram[212][7] ) );
  DFFHQX1 \ram_reg[212][6]  ( .D(n3980), .CK(clk), .Q(\ram[212][6] ) );
  DFFHQX1 \ram_reg[212][5]  ( .D(n3979), .CK(clk), .Q(\ram[212][5] ) );
  DFFHQX1 \ram_reg[212][4]  ( .D(n3978), .CK(clk), .Q(\ram[212][4] ) );
  DFFHQX1 \ram_reg[212][3]  ( .D(n3977), .CK(clk), .Q(\ram[212][3] ) );
  DFFHQX1 \ram_reg[212][2]  ( .D(n3976), .CK(clk), .Q(\ram[212][2] ) );
  DFFHQX1 \ram_reg[212][1]  ( .D(n3975), .CK(clk), .Q(\ram[212][1] ) );
  DFFHQX1 \ram_reg[212][0]  ( .D(n3974), .CK(clk), .Q(\ram[212][0] ) );
  DFFHQX1 \ram_reg[208][15]  ( .D(n3925), .CK(clk), .Q(\ram[208][15] ) );
  DFFHQX1 \ram_reg[208][14]  ( .D(n3924), .CK(clk), .Q(\ram[208][14] ) );
  DFFHQX1 \ram_reg[208][13]  ( .D(n3923), .CK(clk), .Q(\ram[208][13] ) );
  DFFHQX1 \ram_reg[208][12]  ( .D(n3922), .CK(clk), .Q(\ram[208][12] ) );
  DFFHQX1 \ram_reg[208][11]  ( .D(n3921), .CK(clk), .Q(\ram[208][11] ) );
  DFFHQX1 \ram_reg[208][10]  ( .D(n3920), .CK(clk), .Q(\ram[208][10] ) );
  DFFHQX1 \ram_reg[208][9]  ( .D(n3919), .CK(clk), .Q(\ram[208][9] ) );
  DFFHQX1 \ram_reg[208][8]  ( .D(n3918), .CK(clk), .Q(\ram[208][8] ) );
  DFFHQX1 \ram_reg[208][7]  ( .D(n3917), .CK(clk), .Q(\ram[208][7] ) );
  DFFHQX1 \ram_reg[208][6]  ( .D(n3916), .CK(clk), .Q(\ram[208][6] ) );
  DFFHQX1 \ram_reg[208][5]  ( .D(n3915), .CK(clk), .Q(\ram[208][5] ) );
  DFFHQX1 \ram_reg[208][4]  ( .D(n3914), .CK(clk), .Q(\ram[208][4] ) );
  DFFHQX1 \ram_reg[208][3]  ( .D(n3913), .CK(clk), .Q(\ram[208][3] ) );
  DFFHQX1 \ram_reg[208][2]  ( .D(n3912), .CK(clk), .Q(\ram[208][2] ) );
  DFFHQX1 \ram_reg[208][1]  ( .D(n3911), .CK(clk), .Q(\ram[208][1] ) );
  DFFHQX1 \ram_reg[208][0]  ( .D(n3910), .CK(clk), .Q(\ram[208][0] ) );
  DFFHQX1 \ram_reg[204][15]  ( .D(n3861), .CK(clk), .Q(\ram[204][15] ) );
  DFFHQX1 \ram_reg[204][14]  ( .D(n3860), .CK(clk), .Q(\ram[204][14] ) );
  DFFHQX1 \ram_reg[204][13]  ( .D(n3859), .CK(clk), .Q(\ram[204][13] ) );
  DFFHQX1 \ram_reg[204][12]  ( .D(n3858), .CK(clk), .Q(\ram[204][12] ) );
  DFFHQX1 \ram_reg[204][11]  ( .D(n3857), .CK(clk), .Q(\ram[204][11] ) );
  DFFHQX1 \ram_reg[204][10]  ( .D(n3856), .CK(clk), .Q(\ram[204][10] ) );
  DFFHQX1 \ram_reg[204][9]  ( .D(n3855), .CK(clk), .Q(\ram[204][9] ) );
  DFFHQX1 \ram_reg[204][8]  ( .D(n3854), .CK(clk), .Q(\ram[204][8] ) );
  DFFHQX1 \ram_reg[204][7]  ( .D(n3853), .CK(clk), .Q(\ram[204][7] ) );
  DFFHQX1 \ram_reg[204][6]  ( .D(n3852), .CK(clk), .Q(\ram[204][6] ) );
  DFFHQX1 \ram_reg[204][5]  ( .D(n3851), .CK(clk), .Q(\ram[204][5] ) );
  DFFHQX1 \ram_reg[204][4]  ( .D(n3850), .CK(clk), .Q(\ram[204][4] ) );
  DFFHQX1 \ram_reg[204][3]  ( .D(n3849), .CK(clk), .Q(\ram[204][3] ) );
  DFFHQX1 \ram_reg[204][2]  ( .D(n3848), .CK(clk), .Q(\ram[204][2] ) );
  DFFHQX1 \ram_reg[204][1]  ( .D(n3847), .CK(clk), .Q(\ram[204][1] ) );
  DFFHQX1 \ram_reg[204][0]  ( .D(n3846), .CK(clk), .Q(\ram[204][0] ) );
  DFFHQX1 \ram_reg[200][15]  ( .D(n3797), .CK(clk), .Q(\ram[200][15] ) );
  DFFHQX1 \ram_reg[200][14]  ( .D(n3796), .CK(clk), .Q(\ram[200][14] ) );
  DFFHQX1 \ram_reg[200][13]  ( .D(n3795), .CK(clk), .Q(\ram[200][13] ) );
  DFFHQX1 \ram_reg[200][12]  ( .D(n3794), .CK(clk), .Q(\ram[200][12] ) );
  DFFHQX1 \ram_reg[200][11]  ( .D(n3793), .CK(clk), .Q(\ram[200][11] ) );
  DFFHQX1 \ram_reg[200][10]  ( .D(n3792), .CK(clk), .Q(\ram[200][10] ) );
  DFFHQX1 \ram_reg[200][9]  ( .D(n3791), .CK(clk), .Q(\ram[200][9] ) );
  DFFHQX1 \ram_reg[200][8]  ( .D(n3790), .CK(clk), .Q(\ram[200][8] ) );
  DFFHQX1 \ram_reg[200][7]  ( .D(n3789), .CK(clk), .Q(\ram[200][7] ) );
  DFFHQX1 \ram_reg[200][6]  ( .D(n3788), .CK(clk), .Q(\ram[200][6] ) );
  DFFHQX1 \ram_reg[200][5]  ( .D(n3787), .CK(clk), .Q(\ram[200][5] ) );
  DFFHQX1 \ram_reg[200][4]  ( .D(n3786), .CK(clk), .Q(\ram[200][4] ) );
  DFFHQX1 \ram_reg[200][3]  ( .D(n3785), .CK(clk), .Q(\ram[200][3] ) );
  DFFHQX1 \ram_reg[200][2]  ( .D(n3784), .CK(clk), .Q(\ram[200][2] ) );
  DFFHQX1 \ram_reg[200][1]  ( .D(n3783), .CK(clk), .Q(\ram[200][1] ) );
  DFFHQX1 \ram_reg[200][0]  ( .D(n3782), .CK(clk), .Q(\ram[200][0] ) );
  DFFHQX1 \ram_reg[196][15]  ( .D(n3733), .CK(clk), .Q(\ram[196][15] ) );
  DFFHQX1 \ram_reg[196][14]  ( .D(n3732), .CK(clk), .Q(\ram[196][14] ) );
  DFFHQX1 \ram_reg[196][13]  ( .D(n3731), .CK(clk), .Q(\ram[196][13] ) );
  DFFHQX1 \ram_reg[196][12]  ( .D(n3730), .CK(clk), .Q(\ram[196][12] ) );
  DFFHQX1 \ram_reg[196][11]  ( .D(n3729), .CK(clk), .Q(\ram[196][11] ) );
  DFFHQX1 \ram_reg[196][10]  ( .D(n3728), .CK(clk), .Q(\ram[196][10] ) );
  DFFHQX1 \ram_reg[196][9]  ( .D(n3727), .CK(clk), .Q(\ram[196][9] ) );
  DFFHQX1 \ram_reg[196][8]  ( .D(n3726), .CK(clk), .Q(\ram[196][8] ) );
  DFFHQX1 \ram_reg[196][7]  ( .D(n3725), .CK(clk), .Q(\ram[196][7] ) );
  DFFHQX1 \ram_reg[196][6]  ( .D(n3724), .CK(clk), .Q(\ram[196][6] ) );
  DFFHQX1 \ram_reg[196][5]  ( .D(n3723), .CK(clk), .Q(\ram[196][5] ) );
  DFFHQX1 \ram_reg[196][4]  ( .D(n3722), .CK(clk), .Q(\ram[196][4] ) );
  DFFHQX1 \ram_reg[196][3]  ( .D(n3721), .CK(clk), .Q(\ram[196][3] ) );
  DFFHQX1 \ram_reg[196][2]  ( .D(n3720), .CK(clk), .Q(\ram[196][2] ) );
  DFFHQX1 \ram_reg[196][1]  ( .D(n3719), .CK(clk), .Q(\ram[196][1] ) );
  DFFHQX1 \ram_reg[196][0]  ( .D(n3718), .CK(clk), .Q(\ram[196][0] ) );
  DFFHQX1 \ram_reg[192][15]  ( .D(n3669), .CK(clk), .Q(\ram[192][15] ) );
  DFFHQX1 \ram_reg[192][14]  ( .D(n3668), .CK(clk), .Q(\ram[192][14] ) );
  DFFHQX1 \ram_reg[192][13]  ( .D(n3667), .CK(clk), .Q(\ram[192][13] ) );
  DFFHQX1 \ram_reg[192][12]  ( .D(n3666), .CK(clk), .Q(\ram[192][12] ) );
  DFFHQX1 \ram_reg[192][11]  ( .D(n3665), .CK(clk), .Q(\ram[192][11] ) );
  DFFHQX1 \ram_reg[192][10]  ( .D(n3664), .CK(clk), .Q(\ram[192][10] ) );
  DFFHQX1 \ram_reg[192][9]  ( .D(n3663), .CK(clk), .Q(\ram[192][9] ) );
  DFFHQX1 \ram_reg[192][8]  ( .D(n3662), .CK(clk), .Q(\ram[192][8] ) );
  DFFHQX1 \ram_reg[192][7]  ( .D(n3661), .CK(clk), .Q(\ram[192][7] ) );
  DFFHQX1 \ram_reg[192][6]  ( .D(n3660), .CK(clk), .Q(\ram[192][6] ) );
  DFFHQX1 \ram_reg[192][5]  ( .D(n3659), .CK(clk), .Q(\ram[192][5] ) );
  DFFHQX1 \ram_reg[192][4]  ( .D(n3658), .CK(clk), .Q(\ram[192][4] ) );
  DFFHQX1 \ram_reg[192][3]  ( .D(n3657), .CK(clk), .Q(\ram[192][3] ) );
  DFFHQX1 \ram_reg[192][2]  ( .D(n3656), .CK(clk), .Q(\ram[192][2] ) );
  DFFHQX1 \ram_reg[192][1]  ( .D(n3655), .CK(clk), .Q(\ram[192][1] ) );
  DFFHQX1 \ram_reg[192][0]  ( .D(n3654), .CK(clk), .Q(\ram[192][0] ) );
  DFFHQX1 \ram_reg[188][15]  ( .D(n3605), .CK(clk), .Q(\ram[188][15] ) );
  DFFHQX1 \ram_reg[188][14]  ( .D(n3604), .CK(clk), .Q(\ram[188][14] ) );
  DFFHQX1 \ram_reg[188][13]  ( .D(n3603), .CK(clk), .Q(\ram[188][13] ) );
  DFFHQX1 \ram_reg[188][12]  ( .D(n3602), .CK(clk), .Q(\ram[188][12] ) );
  DFFHQX1 \ram_reg[188][11]  ( .D(n3601), .CK(clk), .Q(\ram[188][11] ) );
  DFFHQX1 \ram_reg[188][10]  ( .D(n3600), .CK(clk), .Q(\ram[188][10] ) );
  DFFHQX1 \ram_reg[188][9]  ( .D(n3599), .CK(clk), .Q(\ram[188][9] ) );
  DFFHQX1 \ram_reg[188][8]  ( .D(n3598), .CK(clk), .Q(\ram[188][8] ) );
  DFFHQX1 \ram_reg[188][7]  ( .D(n3597), .CK(clk), .Q(\ram[188][7] ) );
  DFFHQX1 \ram_reg[188][6]  ( .D(n3596), .CK(clk), .Q(\ram[188][6] ) );
  DFFHQX1 \ram_reg[188][5]  ( .D(n3595), .CK(clk), .Q(\ram[188][5] ) );
  DFFHQX1 \ram_reg[188][4]  ( .D(n3594), .CK(clk), .Q(\ram[188][4] ) );
  DFFHQX1 \ram_reg[188][3]  ( .D(n3593), .CK(clk), .Q(\ram[188][3] ) );
  DFFHQX1 \ram_reg[188][2]  ( .D(n3592), .CK(clk), .Q(\ram[188][2] ) );
  DFFHQX1 \ram_reg[188][1]  ( .D(n3591), .CK(clk), .Q(\ram[188][1] ) );
  DFFHQX1 \ram_reg[188][0]  ( .D(n3590), .CK(clk), .Q(\ram[188][0] ) );
  DFFHQX1 \ram_reg[184][15]  ( .D(n3541), .CK(clk), .Q(\ram[184][15] ) );
  DFFHQX1 \ram_reg[184][14]  ( .D(n3540), .CK(clk), .Q(\ram[184][14] ) );
  DFFHQX1 \ram_reg[184][13]  ( .D(n3539), .CK(clk), .Q(\ram[184][13] ) );
  DFFHQX1 \ram_reg[184][12]  ( .D(n3538), .CK(clk), .Q(\ram[184][12] ) );
  DFFHQX1 \ram_reg[184][11]  ( .D(n3537), .CK(clk), .Q(\ram[184][11] ) );
  DFFHQX1 \ram_reg[184][10]  ( .D(n3536), .CK(clk), .Q(\ram[184][10] ) );
  DFFHQX1 \ram_reg[184][9]  ( .D(n3535), .CK(clk), .Q(\ram[184][9] ) );
  DFFHQX1 \ram_reg[184][8]  ( .D(n3534), .CK(clk), .Q(\ram[184][8] ) );
  DFFHQX1 \ram_reg[184][7]  ( .D(n3533), .CK(clk), .Q(\ram[184][7] ) );
  DFFHQX1 \ram_reg[184][6]  ( .D(n3532), .CK(clk), .Q(\ram[184][6] ) );
  DFFHQX1 \ram_reg[184][5]  ( .D(n3531), .CK(clk), .Q(\ram[184][5] ) );
  DFFHQX1 \ram_reg[184][4]  ( .D(n3530), .CK(clk), .Q(\ram[184][4] ) );
  DFFHQX1 \ram_reg[184][3]  ( .D(n3529), .CK(clk), .Q(\ram[184][3] ) );
  DFFHQX1 \ram_reg[184][2]  ( .D(n3528), .CK(clk), .Q(\ram[184][2] ) );
  DFFHQX1 \ram_reg[184][1]  ( .D(n3527), .CK(clk), .Q(\ram[184][1] ) );
  DFFHQX1 \ram_reg[184][0]  ( .D(n3526), .CK(clk), .Q(\ram[184][0] ) );
  DFFHQX1 \ram_reg[180][15]  ( .D(n3477), .CK(clk), .Q(\ram[180][15] ) );
  DFFHQX1 \ram_reg[180][14]  ( .D(n3476), .CK(clk), .Q(\ram[180][14] ) );
  DFFHQX1 \ram_reg[180][13]  ( .D(n3475), .CK(clk), .Q(\ram[180][13] ) );
  DFFHQX1 \ram_reg[180][12]  ( .D(n3474), .CK(clk), .Q(\ram[180][12] ) );
  DFFHQX1 \ram_reg[180][11]  ( .D(n3473), .CK(clk), .Q(\ram[180][11] ) );
  DFFHQX1 \ram_reg[180][10]  ( .D(n3472), .CK(clk), .Q(\ram[180][10] ) );
  DFFHQX1 \ram_reg[180][9]  ( .D(n3471), .CK(clk), .Q(\ram[180][9] ) );
  DFFHQX1 \ram_reg[180][8]  ( .D(n3470), .CK(clk), .Q(\ram[180][8] ) );
  DFFHQX1 \ram_reg[180][7]  ( .D(n3469), .CK(clk), .Q(\ram[180][7] ) );
  DFFHQX1 \ram_reg[180][6]  ( .D(n3468), .CK(clk), .Q(\ram[180][6] ) );
  DFFHQX1 \ram_reg[180][5]  ( .D(n3467), .CK(clk), .Q(\ram[180][5] ) );
  DFFHQX1 \ram_reg[180][4]  ( .D(n3466), .CK(clk), .Q(\ram[180][4] ) );
  DFFHQX1 \ram_reg[180][3]  ( .D(n3465), .CK(clk), .Q(\ram[180][3] ) );
  DFFHQX1 \ram_reg[180][2]  ( .D(n3464), .CK(clk), .Q(\ram[180][2] ) );
  DFFHQX1 \ram_reg[180][1]  ( .D(n3463), .CK(clk), .Q(\ram[180][1] ) );
  DFFHQX1 \ram_reg[180][0]  ( .D(n3462), .CK(clk), .Q(\ram[180][0] ) );
  DFFHQX1 \ram_reg[176][15]  ( .D(n3413), .CK(clk), .Q(\ram[176][15] ) );
  DFFHQX1 \ram_reg[176][14]  ( .D(n3412), .CK(clk), .Q(\ram[176][14] ) );
  DFFHQX1 \ram_reg[176][13]  ( .D(n3411), .CK(clk), .Q(\ram[176][13] ) );
  DFFHQX1 \ram_reg[176][12]  ( .D(n3410), .CK(clk), .Q(\ram[176][12] ) );
  DFFHQX1 \ram_reg[176][11]  ( .D(n3409), .CK(clk), .Q(\ram[176][11] ) );
  DFFHQX1 \ram_reg[176][10]  ( .D(n3408), .CK(clk), .Q(\ram[176][10] ) );
  DFFHQX1 \ram_reg[176][9]  ( .D(n3407), .CK(clk), .Q(\ram[176][9] ) );
  DFFHQX1 \ram_reg[176][8]  ( .D(n3406), .CK(clk), .Q(\ram[176][8] ) );
  DFFHQX1 \ram_reg[176][7]  ( .D(n3405), .CK(clk), .Q(\ram[176][7] ) );
  DFFHQX1 \ram_reg[176][6]  ( .D(n3404), .CK(clk), .Q(\ram[176][6] ) );
  DFFHQX1 \ram_reg[176][5]  ( .D(n3403), .CK(clk), .Q(\ram[176][5] ) );
  DFFHQX1 \ram_reg[176][4]  ( .D(n3402), .CK(clk), .Q(\ram[176][4] ) );
  DFFHQX1 \ram_reg[176][3]  ( .D(n3401), .CK(clk), .Q(\ram[176][3] ) );
  DFFHQX1 \ram_reg[176][2]  ( .D(n3400), .CK(clk), .Q(\ram[176][2] ) );
  DFFHQX1 \ram_reg[176][1]  ( .D(n3399), .CK(clk), .Q(\ram[176][1] ) );
  DFFHQX1 \ram_reg[176][0]  ( .D(n3398), .CK(clk), .Q(\ram[176][0] ) );
  DFFHQX1 \ram_reg[172][15]  ( .D(n3349), .CK(clk), .Q(\ram[172][15] ) );
  DFFHQX1 \ram_reg[172][14]  ( .D(n3348), .CK(clk), .Q(\ram[172][14] ) );
  DFFHQX1 \ram_reg[172][13]  ( .D(n3347), .CK(clk), .Q(\ram[172][13] ) );
  DFFHQX1 \ram_reg[172][12]  ( .D(n3346), .CK(clk), .Q(\ram[172][12] ) );
  DFFHQX1 \ram_reg[172][11]  ( .D(n3345), .CK(clk), .Q(\ram[172][11] ) );
  DFFHQX1 \ram_reg[172][10]  ( .D(n3344), .CK(clk), .Q(\ram[172][10] ) );
  DFFHQX1 \ram_reg[172][9]  ( .D(n3343), .CK(clk), .Q(\ram[172][9] ) );
  DFFHQX1 \ram_reg[172][8]  ( .D(n3342), .CK(clk), .Q(\ram[172][8] ) );
  DFFHQX1 \ram_reg[172][7]  ( .D(n3341), .CK(clk), .Q(\ram[172][7] ) );
  DFFHQX1 \ram_reg[172][6]  ( .D(n3340), .CK(clk), .Q(\ram[172][6] ) );
  DFFHQX1 \ram_reg[172][5]  ( .D(n3339), .CK(clk), .Q(\ram[172][5] ) );
  DFFHQX1 \ram_reg[172][4]  ( .D(n3338), .CK(clk), .Q(\ram[172][4] ) );
  DFFHQX1 \ram_reg[172][3]  ( .D(n3337), .CK(clk), .Q(\ram[172][3] ) );
  DFFHQX1 \ram_reg[172][2]  ( .D(n3336), .CK(clk), .Q(\ram[172][2] ) );
  DFFHQX1 \ram_reg[172][1]  ( .D(n3335), .CK(clk), .Q(\ram[172][1] ) );
  DFFHQX1 \ram_reg[172][0]  ( .D(n3334), .CK(clk), .Q(\ram[172][0] ) );
  DFFHQX1 \ram_reg[168][15]  ( .D(n3285), .CK(clk), .Q(\ram[168][15] ) );
  DFFHQX1 \ram_reg[168][14]  ( .D(n3284), .CK(clk), .Q(\ram[168][14] ) );
  DFFHQX1 \ram_reg[168][13]  ( .D(n3283), .CK(clk), .Q(\ram[168][13] ) );
  DFFHQX1 \ram_reg[168][12]  ( .D(n3282), .CK(clk), .Q(\ram[168][12] ) );
  DFFHQX1 \ram_reg[168][11]  ( .D(n3281), .CK(clk), .Q(\ram[168][11] ) );
  DFFHQX1 \ram_reg[168][10]  ( .D(n3280), .CK(clk), .Q(\ram[168][10] ) );
  DFFHQX1 \ram_reg[168][9]  ( .D(n3279), .CK(clk), .Q(\ram[168][9] ) );
  DFFHQX1 \ram_reg[168][8]  ( .D(n3278), .CK(clk), .Q(\ram[168][8] ) );
  DFFHQX1 \ram_reg[168][7]  ( .D(n3277), .CK(clk), .Q(\ram[168][7] ) );
  DFFHQX1 \ram_reg[168][6]  ( .D(n3276), .CK(clk), .Q(\ram[168][6] ) );
  DFFHQX1 \ram_reg[168][5]  ( .D(n3275), .CK(clk), .Q(\ram[168][5] ) );
  DFFHQX1 \ram_reg[168][4]  ( .D(n3274), .CK(clk), .Q(\ram[168][4] ) );
  DFFHQX1 \ram_reg[168][3]  ( .D(n3273), .CK(clk), .Q(\ram[168][3] ) );
  DFFHQX1 \ram_reg[168][2]  ( .D(n3272), .CK(clk), .Q(\ram[168][2] ) );
  DFFHQX1 \ram_reg[168][1]  ( .D(n3271), .CK(clk), .Q(\ram[168][1] ) );
  DFFHQX1 \ram_reg[168][0]  ( .D(n3270), .CK(clk), .Q(\ram[168][0] ) );
  DFFHQX1 \ram_reg[164][15]  ( .D(n3221), .CK(clk), .Q(\ram[164][15] ) );
  DFFHQX1 \ram_reg[164][14]  ( .D(n3220), .CK(clk), .Q(\ram[164][14] ) );
  DFFHQX1 \ram_reg[164][13]  ( .D(n3219), .CK(clk), .Q(\ram[164][13] ) );
  DFFHQX1 \ram_reg[164][12]  ( .D(n3218), .CK(clk), .Q(\ram[164][12] ) );
  DFFHQX1 \ram_reg[164][11]  ( .D(n3217), .CK(clk), .Q(\ram[164][11] ) );
  DFFHQX1 \ram_reg[164][10]  ( .D(n3216), .CK(clk), .Q(\ram[164][10] ) );
  DFFHQX1 \ram_reg[164][9]  ( .D(n3215), .CK(clk), .Q(\ram[164][9] ) );
  DFFHQX1 \ram_reg[164][8]  ( .D(n3214), .CK(clk), .Q(\ram[164][8] ) );
  DFFHQX1 \ram_reg[164][7]  ( .D(n3213), .CK(clk), .Q(\ram[164][7] ) );
  DFFHQX1 \ram_reg[164][6]  ( .D(n3212), .CK(clk), .Q(\ram[164][6] ) );
  DFFHQX1 \ram_reg[164][5]  ( .D(n3211), .CK(clk), .Q(\ram[164][5] ) );
  DFFHQX1 \ram_reg[164][4]  ( .D(n3210), .CK(clk), .Q(\ram[164][4] ) );
  DFFHQX1 \ram_reg[164][3]  ( .D(n3209), .CK(clk), .Q(\ram[164][3] ) );
  DFFHQX1 \ram_reg[164][2]  ( .D(n3208), .CK(clk), .Q(\ram[164][2] ) );
  DFFHQX1 \ram_reg[164][1]  ( .D(n3207), .CK(clk), .Q(\ram[164][1] ) );
  DFFHQX1 \ram_reg[164][0]  ( .D(n3206), .CK(clk), .Q(\ram[164][0] ) );
  DFFHQX1 \ram_reg[160][15]  ( .D(n3157), .CK(clk), .Q(\ram[160][15] ) );
  DFFHQX1 \ram_reg[160][14]  ( .D(n3156), .CK(clk), .Q(\ram[160][14] ) );
  DFFHQX1 \ram_reg[160][13]  ( .D(n3155), .CK(clk), .Q(\ram[160][13] ) );
  DFFHQX1 \ram_reg[160][12]  ( .D(n3154), .CK(clk), .Q(\ram[160][12] ) );
  DFFHQX1 \ram_reg[160][11]  ( .D(n3153), .CK(clk), .Q(\ram[160][11] ) );
  DFFHQX1 \ram_reg[160][10]  ( .D(n3152), .CK(clk), .Q(\ram[160][10] ) );
  DFFHQX1 \ram_reg[160][9]  ( .D(n3151), .CK(clk), .Q(\ram[160][9] ) );
  DFFHQX1 \ram_reg[160][8]  ( .D(n3150), .CK(clk), .Q(\ram[160][8] ) );
  DFFHQX1 \ram_reg[160][7]  ( .D(n3149), .CK(clk), .Q(\ram[160][7] ) );
  DFFHQX1 \ram_reg[160][6]  ( .D(n3148), .CK(clk), .Q(\ram[160][6] ) );
  DFFHQX1 \ram_reg[160][5]  ( .D(n3147), .CK(clk), .Q(\ram[160][5] ) );
  DFFHQX1 \ram_reg[160][4]  ( .D(n3146), .CK(clk), .Q(\ram[160][4] ) );
  DFFHQX1 \ram_reg[160][3]  ( .D(n3145), .CK(clk), .Q(\ram[160][3] ) );
  DFFHQX1 \ram_reg[160][2]  ( .D(n3144), .CK(clk), .Q(\ram[160][2] ) );
  DFFHQX1 \ram_reg[160][1]  ( .D(n3143), .CK(clk), .Q(\ram[160][1] ) );
  DFFHQX1 \ram_reg[160][0]  ( .D(n3142), .CK(clk), .Q(\ram[160][0] ) );
  DFFHQX1 \ram_reg[156][15]  ( .D(n3093), .CK(clk), .Q(\ram[156][15] ) );
  DFFHQX1 \ram_reg[156][14]  ( .D(n3092), .CK(clk), .Q(\ram[156][14] ) );
  DFFHQX1 \ram_reg[156][13]  ( .D(n3091), .CK(clk), .Q(\ram[156][13] ) );
  DFFHQX1 \ram_reg[156][12]  ( .D(n3090), .CK(clk), .Q(\ram[156][12] ) );
  DFFHQX1 \ram_reg[156][11]  ( .D(n3089), .CK(clk), .Q(\ram[156][11] ) );
  DFFHQX1 \ram_reg[156][10]  ( .D(n3088), .CK(clk), .Q(\ram[156][10] ) );
  DFFHQX1 \ram_reg[156][9]  ( .D(n3087), .CK(clk), .Q(\ram[156][9] ) );
  DFFHQX1 \ram_reg[156][8]  ( .D(n3086), .CK(clk), .Q(\ram[156][8] ) );
  DFFHQX1 \ram_reg[156][7]  ( .D(n3085), .CK(clk), .Q(\ram[156][7] ) );
  DFFHQX1 \ram_reg[156][6]  ( .D(n3084), .CK(clk), .Q(\ram[156][6] ) );
  DFFHQX1 \ram_reg[156][5]  ( .D(n3083), .CK(clk), .Q(\ram[156][5] ) );
  DFFHQX1 \ram_reg[156][4]  ( .D(n3082), .CK(clk), .Q(\ram[156][4] ) );
  DFFHQX1 \ram_reg[156][3]  ( .D(n3081), .CK(clk), .Q(\ram[156][3] ) );
  DFFHQX1 \ram_reg[156][2]  ( .D(n3080), .CK(clk), .Q(\ram[156][2] ) );
  DFFHQX1 \ram_reg[156][1]  ( .D(n3079), .CK(clk), .Q(\ram[156][1] ) );
  DFFHQX1 \ram_reg[156][0]  ( .D(n3078), .CK(clk), .Q(\ram[156][0] ) );
  DFFHQX1 \ram_reg[152][15]  ( .D(n3029), .CK(clk), .Q(\ram[152][15] ) );
  DFFHQX1 \ram_reg[152][14]  ( .D(n3028), .CK(clk), .Q(\ram[152][14] ) );
  DFFHQX1 \ram_reg[152][13]  ( .D(n3027), .CK(clk), .Q(\ram[152][13] ) );
  DFFHQX1 \ram_reg[152][12]  ( .D(n3026), .CK(clk), .Q(\ram[152][12] ) );
  DFFHQX1 \ram_reg[152][11]  ( .D(n3025), .CK(clk), .Q(\ram[152][11] ) );
  DFFHQX1 \ram_reg[152][10]  ( .D(n3024), .CK(clk), .Q(\ram[152][10] ) );
  DFFHQX1 \ram_reg[152][9]  ( .D(n3023), .CK(clk), .Q(\ram[152][9] ) );
  DFFHQX1 \ram_reg[152][8]  ( .D(n3022), .CK(clk), .Q(\ram[152][8] ) );
  DFFHQX1 \ram_reg[152][7]  ( .D(n3021), .CK(clk), .Q(\ram[152][7] ) );
  DFFHQX1 \ram_reg[152][6]  ( .D(n3020), .CK(clk), .Q(\ram[152][6] ) );
  DFFHQX1 \ram_reg[152][5]  ( .D(n3019), .CK(clk), .Q(\ram[152][5] ) );
  DFFHQX1 \ram_reg[152][4]  ( .D(n3018), .CK(clk), .Q(\ram[152][4] ) );
  DFFHQX1 \ram_reg[152][3]  ( .D(n3017), .CK(clk), .Q(\ram[152][3] ) );
  DFFHQX1 \ram_reg[152][2]  ( .D(n3016), .CK(clk), .Q(\ram[152][2] ) );
  DFFHQX1 \ram_reg[152][1]  ( .D(n3015), .CK(clk), .Q(\ram[152][1] ) );
  DFFHQX1 \ram_reg[152][0]  ( .D(n3014), .CK(clk), .Q(\ram[152][0] ) );
  DFFHQX1 \ram_reg[148][15]  ( .D(n2965), .CK(clk), .Q(\ram[148][15] ) );
  DFFHQX1 \ram_reg[148][14]  ( .D(n2964), .CK(clk), .Q(\ram[148][14] ) );
  DFFHQX1 \ram_reg[148][13]  ( .D(n2963), .CK(clk), .Q(\ram[148][13] ) );
  DFFHQX1 \ram_reg[148][12]  ( .D(n2962), .CK(clk), .Q(\ram[148][12] ) );
  DFFHQX1 \ram_reg[148][11]  ( .D(n2961), .CK(clk), .Q(\ram[148][11] ) );
  DFFHQX1 \ram_reg[148][10]  ( .D(n2960), .CK(clk), .Q(\ram[148][10] ) );
  DFFHQX1 \ram_reg[148][9]  ( .D(n2959), .CK(clk), .Q(\ram[148][9] ) );
  DFFHQX1 \ram_reg[148][8]  ( .D(n2958), .CK(clk), .Q(\ram[148][8] ) );
  DFFHQX1 \ram_reg[148][7]  ( .D(n2957), .CK(clk), .Q(\ram[148][7] ) );
  DFFHQX1 \ram_reg[148][6]  ( .D(n2956), .CK(clk), .Q(\ram[148][6] ) );
  DFFHQX1 \ram_reg[148][5]  ( .D(n2955), .CK(clk), .Q(\ram[148][5] ) );
  DFFHQX1 \ram_reg[148][4]  ( .D(n2954), .CK(clk), .Q(\ram[148][4] ) );
  DFFHQX1 \ram_reg[148][3]  ( .D(n2953), .CK(clk), .Q(\ram[148][3] ) );
  DFFHQX1 \ram_reg[148][2]  ( .D(n2952), .CK(clk), .Q(\ram[148][2] ) );
  DFFHQX1 \ram_reg[148][1]  ( .D(n2951), .CK(clk), .Q(\ram[148][1] ) );
  DFFHQX1 \ram_reg[148][0]  ( .D(n2950), .CK(clk), .Q(\ram[148][0] ) );
  DFFHQX1 \ram_reg[144][15]  ( .D(n2901), .CK(clk), .Q(\ram[144][15] ) );
  DFFHQX1 \ram_reg[144][14]  ( .D(n2900), .CK(clk), .Q(\ram[144][14] ) );
  DFFHQX1 \ram_reg[144][13]  ( .D(n2899), .CK(clk), .Q(\ram[144][13] ) );
  DFFHQX1 \ram_reg[144][12]  ( .D(n2898), .CK(clk), .Q(\ram[144][12] ) );
  DFFHQX1 \ram_reg[144][11]  ( .D(n2897), .CK(clk), .Q(\ram[144][11] ) );
  DFFHQX1 \ram_reg[144][10]  ( .D(n2896), .CK(clk), .Q(\ram[144][10] ) );
  DFFHQX1 \ram_reg[144][9]  ( .D(n2895), .CK(clk), .Q(\ram[144][9] ) );
  DFFHQX1 \ram_reg[144][8]  ( .D(n2894), .CK(clk), .Q(\ram[144][8] ) );
  DFFHQX1 \ram_reg[144][7]  ( .D(n2893), .CK(clk), .Q(\ram[144][7] ) );
  DFFHQX1 \ram_reg[144][6]  ( .D(n2892), .CK(clk), .Q(\ram[144][6] ) );
  DFFHQX1 \ram_reg[144][5]  ( .D(n2891), .CK(clk), .Q(\ram[144][5] ) );
  DFFHQX1 \ram_reg[144][4]  ( .D(n2890), .CK(clk), .Q(\ram[144][4] ) );
  DFFHQX1 \ram_reg[144][3]  ( .D(n2889), .CK(clk), .Q(\ram[144][3] ) );
  DFFHQX1 \ram_reg[144][2]  ( .D(n2888), .CK(clk), .Q(\ram[144][2] ) );
  DFFHQX1 \ram_reg[144][1]  ( .D(n2887), .CK(clk), .Q(\ram[144][1] ) );
  DFFHQX1 \ram_reg[144][0]  ( .D(n2886), .CK(clk), .Q(\ram[144][0] ) );
  DFFHQX1 \ram_reg[140][15]  ( .D(n2837), .CK(clk), .Q(\ram[140][15] ) );
  DFFHQX1 \ram_reg[140][14]  ( .D(n2836), .CK(clk), .Q(\ram[140][14] ) );
  DFFHQX1 \ram_reg[140][13]  ( .D(n2835), .CK(clk), .Q(\ram[140][13] ) );
  DFFHQX1 \ram_reg[140][12]  ( .D(n2834), .CK(clk), .Q(\ram[140][12] ) );
  DFFHQX1 \ram_reg[140][11]  ( .D(n2833), .CK(clk), .Q(\ram[140][11] ) );
  DFFHQX1 \ram_reg[140][10]  ( .D(n2832), .CK(clk), .Q(\ram[140][10] ) );
  DFFHQX1 \ram_reg[140][9]  ( .D(n2831), .CK(clk), .Q(\ram[140][9] ) );
  DFFHQX1 \ram_reg[140][8]  ( .D(n2830), .CK(clk), .Q(\ram[140][8] ) );
  DFFHQX1 \ram_reg[140][7]  ( .D(n2829), .CK(clk), .Q(\ram[140][7] ) );
  DFFHQX1 \ram_reg[140][6]  ( .D(n2828), .CK(clk), .Q(\ram[140][6] ) );
  DFFHQX1 \ram_reg[140][5]  ( .D(n2827), .CK(clk), .Q(\ram[140][5] ) );
  DFFHQX1 \ram_reg[140][4]  ( .D(n2826), .CK(clk), .Q(\ram[140][4] ) );
  DFFHQX1 \ram_reg[140][3]  ( .D(n2825), .CK(clk), .Q(\ram[140][3] ) );
  DFFHQX1 \ram_reg[140][2]  ( .D(n2824), .CK(clk), .Q(\ram[140][2] ) );
  DFFHQX1 \ram_reg[140][1]  ( .D(n2823), .CK(clk), .Q(\ram[140][1] ) );
  DFFHQX1 \ram_reg[140][0]  ( .D(n2822), .CK(clk), .Q(\ram[140][0] ) );
  DFFHQX1 \ram_reg[136][15]  ( .D(n2773), .CK(clk), .Q(\ram[136][15] ) );
  DFFHQX1 \ram_reg[136][14]  ( .D(n2772), .CK(clk), .Q(\ram[136][14] ) );
  DFFHQX1 \ram_reg[136][13]  ( .D(n2771), .CK(clk), .Q(\ram[136][13] ) );
  DFFHQX1 \ram_reg[136][12]  ( .D(n2770), .CK(clk), .Q(\ram[136][12] ) );
  DFFHQX1 \ram_reg[136][11]  ( .D(n2769), .CK(clk), .Q(\ram[136][11] ) );
  DFFHQX1 \ram_reg[136][10]  ( .D(n2768), .CK(clk), .Q(\ram[136][10] ) );
  DFFHQX1 \ram_reg[136][9]  ( .D(n2767), .CK(clk), .Q(\ram[136][9] ) );
  DFFHQX1 \ram_reg[136][8]  ( .D(n2766), .CK(clk), .Q(\ram[136][8] ) );
  DFFHQX1 \ram_reg[136][7]  ( .D(n2765), .CK(clk), .Q(\ram[136][7] ) );
  DFFHQX1 \ram_reg[136][6]  ( .D(n2764), .CK(clk), .Q(\ram[136][6] ) );
  DFFHQX1 \ram_reg[136][5]  ( .D(n2763), .CK(clk), .Q(\ram[136][5] ) );
  DFFHQX1 \ram_reg[136][4]  ( .D(n2762), .CK(clk), .Q(\ram[136][4] ) );
  DFFHQX1 \ram_reg[136][3]  ( .D(n2761), .CK(clk), .Q(\ram[136][3] ) );
  DFFHQX1 \ram_reg[136][2]  ( .D(n2760), .CK(clk), .Q(\ram[136][2] ) );
  DFFHQX1 \ram_reg[136][1]  ( .D(n2759), .CK(clk), .Q(\ram[136][1] ) );
  DFFHQX1 \ram_reg[136][0]  ( .D(n2758), .CK(clk), .Q(\ram[136][0] ) );
  DFFHQX1 \ram_reg[132][15]  ( .D(n2709), .CK(clk), .Q(\ram[132][15] ) );
  DFFHQX1 \ram_reg[132][14]  ( .D(n2708), .CK(clk), .Q(\ram[132][14] ) );
  DFFHQX1 \ram_reg[132][13]  ( .D(n2707), .CK(clk), .Q(\ram[132][13] ) );
  DFFHQX1 \ram_reg[132][12]  ( .D(n2706), .CK(clk), .Q(\ram[132][12] ) );
  DFFHQX1 \ram_reg[132][11]  ( .D(n2705), .CK(clk), .Q(\ram[132][11] ) );
  DFFHQX1 \ram_reg[132][10]  ( .D(n2704), .CK(clk), .Q(\ram[132][10] ) );
  DFFHQX1 \ram_reg[132][9]  ( .D(n2703), .CK(clk), .Q(\ram[132][9] ) );
  DFFHQX1 \ram_reg[132][8]  ( .D(n2702), .CK(clk), .Q(\ram[132][8] ) );
  DFFHQX1 \ram_reg[132][7]  ( .D(n2701), .CK(clk), .Q(\ram[132][7] ) );
  DFFHQX1 \ram_reg[132][6]  ( .D(n2700), .CK(clk), .Q(\ram[132][6] ) );
  DFFHQX1 \ram_reg[132][5]  ( .D(n2699), .CK(clk), .Q(\ram[132][5] ) );
  DFFHQX1 \ram_reg[132][4]  ( .D(n2698), .CK(clk), .Q(\ram[132][4] ) );
  DFFHQX1 \ram_reg[132][3]  ( .D(n2697), .CK(clk), .Q(\ram[132][3] ) );
  DFFHQX1 \ram_reg[132][2]  ( .D(n2696), .CK(clk), .Q(\ram[132][2] ) );
  DFFHQX1 \ram_reg[132][1]  ( .D(n2695), .CK(clk), .Q(\ram[132][1] ) );
  DFFHQX1 \ram_reg[132][0]  ( .D(n2694), .CK(clk), .Q(\ram[132][0] ) );
  DFFHQX1 \ram_reg[128][15]  ( .D(n2645), .CK(clk), .Q(\ram[128][15] ) );
  DFFHQX1 \ram_reg[128][14]  ( .D(n2644), .CK(clk), .Q(\ram[128][14] ) );
  DFFHQX1 \ram_reg[128][13]  ( .D(n2643), .CK(clk), .Q(\ram[128][13] ) );
  DFFHQX1 \ram_reg[128][12]  ( .D(n2642), .CK(clk), .Q(\ram[128][12] ) );
  DFFHQX1 \ram_reg[128][11]  ( .D(n2641), .CK(clk), .Q(\ram[128][11] ) );
  DFFHQX1 \ram_reg[128][10]  ( .D(n2640), .CK(clk), .Q(\ram[128][10] ) );
  DFFHQX1 \ram_reg[128][9]  ( .D(n2639), .CK(clk), .Q(\ram[128][9] ) );
  DFFHQX1 \ram_reg[128][8]  ( .D(n2638), .CK(clk), .Q(\ram[128][8] ) );
  DFFHQX1 \ram_reg[128][7]  ( .D(n2637), .CK(clk), .Q(\ram[128][7] ) );
  DFFHQX1 \ram_reg[128][6]  ( .D(n2636), .CK(clk), .Q(\ram[128][6] ) );
  DFFHQX1 \ram_reg[128][5]  ( .D(n2635), .CK(clk), .Q(\ram[128][5] ) );
  DFFHQX1 \ram_reg[128][4]  ( .D(n2634), .CK(clk), .Q(\ram[128][4] ) );
  DFFHQX1 \ram_reg[128][3]  ( .D(n2633), .CK(clk), .Q(\ram[128][3] ) );
  DFFHQX1 \ram_reg[128][2]  ( .D(n2632), .CK(clk), .Q(\ram[128][2] ) );
  DFFHQX1 \ram_reg[128][1]  ( .D(n2631), .CK(clk), .Q(\ram[128][1] ) );
  DFFHQX1 \ram_reg[128][0]  ( .D(n2630), .CK(clk), .Q(\ram[128][0] ) );
  DFFHQX1 \ram_reg[124][15]  ( .D(n2581), .CK(clk), .Q(\ram[124][15] ) );
  DFFHQX1 \ram_reg[124][14]  ( .D(n2580), .CK(clk), .Q(\ram[124][14] ) );
  DFFHQX1 \ram_reg[124][13]  ( .D(n2579), .CK(clk), .Q(\ram[124][13] ) );
  DFFHQX1 \ram_reg[124][12]  ( .D(n2578), .CK(clk), .Q(\ram[124][12] ) );
  DFFHQX1 \ram_reg[124][11]  ( .D(n2577), .CK(clk), .Q(\ram[124][11] ) );
  DFFHQX1 \ram_reg[124][10]  ( .D(n2576), .CK(clk), .Q(\ram[124][10] ) );
  DFFHQX1 \ram_reg[124][9]  ( .D(n2575), .CK(clk), .Q(\ram[124][9] ) );
  DFFHQX1 \ram_reg[124][8]  ( .D(n2574), .CK(clk), .Q(\ram[124][8] ) );
  DFFHQX1 \ram_reg[124][7]  ( .D(n2573), .CK(clk), .Q(\ram[124][7] ) );
  DFFHQX1 \ram_reg[124][6]  ( .D(n2572), .CK(clk), .Q(\ram[124][6] ) );
  DFFHQX1 \ram_reg[124][5]  ( .D(n2571), .CK(clk), .Q(\ram[124][5] ) );
  DFFHQX1 \ram_reg[124][4]  ( .D(n2570), .CK(clk), .Q(\ram[124][4] ) );
  DFFHQX1 \ram_reg[124][3]  ( .D(n2569), .CK(clk), .Q(\ram[124][3] ) );
  DFFHQX1 \ram_reg[124][2]  ( .D(n2568), .CK(clk), .Q(\ram[124][2] ) );
  DFFHQX1 \ram_reg[124][1]  ( .D(n2567), .CK(clk), .Q(\ram[124][1] ) );
  DFFHQX1 \ram_reg[124][0]  ( .D(n2566), .CK(clk), .Q(\ram[124][0] ) );
  DFFHQX1 \ram_reg[120][15]  ( .D(n2517), .CK(clk), .Q(\ram[120][15] ) );
  DFFHQX1 \ram_reg[120][14]  ( .D(n2516), .CK(clk), .Q(\ram[120][14] ) );
  DFFHQX1 \ram_reg[120][13]  ( .D(n2515), .CK(clk), .Q(\ram[120][13] ) );
  DFFHQX1 \ram_reg[120][12]  ( .D(n2514), .CK(clk), .Q(\ram[120][12] ) );
  DFFHQX1 \ram_reg[120][11]  ( .D(n2513), .CK(clk), .Q(\ram[120][11] ) );
  DFFHQX1 \ram_reg[120][10]  ( .D(n2512), .CK(clk), .Q(\ram[120][10] ) );
  DFFHQX1 \ram_reg[120][9]  ( .D(n2511), .CK(clk), .Q(\ram[120][9] ) );
  DFFHQX1 \ram_reg[120][8]  ( .D(n2510), .CK(clk), .Q(\ram[120][8] ) );
  DFFHQX1 \ram_reg[120][7]  ( .D(n2509), .CK(clk), .Q(\ram[120][7] ) );
  DFFHQX1 \ram_reg[120][6]  ( .D(n2508), .CK(clk), .Q(\ram[120][6] ) );
  DFFHQX1 \ram_reg[120][5]  ( .D(n2507), .CK(clk), .Q(\ram[120][5] ) );
  DFFHQX1 \ram_reg[120][4]  ( .D(n2506), .CK(clk), .Q(\ram[120][4] ) );
  DFFHQX1 \ram_reg[120][3]  ( .D(n2505), .CK(clk), .Q(\ram[120][3] ) );
  DFFHQX1 \ram_reg[120][2]  ( .D(n2504), .CK(clk), .Q(\ram[120][2] ) );
  DFFHQX1 \ram_reg[120][1]  ( .D(n2503), .CK(clk), .Q(\ram[120][1] ) );
  DFFHQX1 \ram_reg[120][0]  ( .D(n2502), .CK(clk), .Q(\ram[120][0] ) );
  DFFHQX1 \ram_reg[116][15]  ( .D(n2453), .CK(clk), .Q(\ram[116][15] ) );
  DFFHQX1 \ram_reg[116][14]  ( .D(n2452), .CK(clk), .Q(\ram[116][14] ) );
  DFFHQX1 \ram_reg[116][13]  ( .D(n2451), .CK(clk), .Q(\ram[116][13] ) );
  DFFHQX1 \ram_reg[116][12]  ( .D(n2450), .CK(clk), .Q(\ram[116][12] ) );
  DFFHQX1 \ram_reg[116][11]  ( .D(n2449), .CK(clk), .Q(\ram[116][11] ) );
  DFFHQX1 \ram_reg[116][10]  ( .D(n2448), .CK(clk), .Q(\ram[116][10] ) );
  DFFHQX1 \ram_reg[116][9]  ( .D(n2447), .CK(clk), .Q(\ram[116][9] ) );
  DFFHQX1 \ram_reg[116][8]  ( .D(n2446), .CK(clk), .Q(\ram[116][8] ) );
  DFFHQX1 \ram_reg[116][7]  ( .D(n2445), .CK(clk), .Q(\ram[116][7] ) );
  DFFHQX1 \ram_reg[116][6]  ( .D(n2444), .CK(clk), .Q(\ram[116][6] ) );
  DFFHQX1 \ram_reg[116][5]  ( .D(n2443), .CK(clk), .Q(\ram[116][5] ) );
  DFFHQX1 \ram_reg[116][4]  ( .D(n2442), .CK(clk), .Q(\ram[116][4] ) );
  DFFHQX1 \ram_reg[116][3]  ( .D(n2441), .CK(clk), .Q(\ram[116][3] ) );
  DFFHQX1 \ram_reg[116][2]  ( .D(n2440), .CK(clk), .Q(\ram[116][2] ) );
  DFFHQX1 \ram_reg[116][1]  ( .D(n2439), .CK(clk), .Q(\ram[116][1] ) );
  DFFHQX1 \ram_reg[116][0]  ( .D(n2438), .CK(clk), .Q(\ram[116][0] ) );
  DFFHQX1 \ram_reg[112][15]  ( .D(n2389), .CK(clk), .Q(\ram[112][15] ) );
  DFFHQX1 \ram_reg[112][14]  ( .D(n2388), .CK(clk), .Q(\ram[112][14] ) );
  DFFHQX1 \ram_reg[112][13]  ( .D(n2387), .CK(clk), .Q(\ram[112][13] ) );
  DFFHQX1 \ram_reg[112][12]  ( .D(n2386), .CK(clk), .Q(\ram[112][12] ) );
  DFFHQX1 \ram_reg[112][11]  ( .D(n2385), .CK(clk), .Q(\ram[112][11] ) );
  DFFHQX1 \ram_reg[112][10]  ( .D(n2384), .CK(clk), .Q(\ram[112][10] ) );
  DFFHQX1 \ram_reg[112][9]  ( .D(n2383), .CK(clk), .Q(\ram[112][9] ) );
  DFFHQX1 \ram_reg[112][8]  ( .D(n2382), .CK(clk), .Q(\ram[112][8] ) );
  DFFHQX1 \ram_reg[112][7]  ( .D(n2381), .CK(clk), .Q(\ram[112][7] ) );
  DFFHQX1 \ram_reg[112][6]  ( .D(n2380), .CK(clk), .Q(\ram[112][6] ) );
  DFFHQX1 \ram_reg[112][5]  ( .D(n2379), .CK(clk), .Q(\ram[112][5] ) );
  DFFHQX1 \ram_reg[112][4]  ( .D(n2378), .CK(clk), .Q(\ram[112][4] ) );
  DFFHQX1 \ram_reg[112][3]  ( .D(n2377), .CK(clk), .Q(\ram[112][3] ) );
  DFFHQX1 \ram_reg[112][2]  ( .D(n2376), .CK(clk), .Q(\ram[112][2] ) );
  DFFHQX1 \ram_reg[112][1]  ( .D(n2375), .CK(clk), .Q(\ram[112][1] ) );
  DFFHQX1 \ram_reg[112][0]  ( .D(n2374), .CK(clk), .Q(\ram[112][0] ) );
  DFFHQX1 \ram_reg[108][15]  ( .D(n2325), .CK(clk), .Q(\ram[108][15] ) );
  DFFHQX1 \ram_reg[108][14]  ( .D(n2324), .CK(clk), .Q(\ram[108][14] ) );
  DFFHQX1 \ram_reg[108][13]  ( .D(n2323), .CK(clk), .Q(\ram[108][13] ) );
  DFFHQX1 \ram_reg[108][12]  ( .D(n2322), .CK(clk), .Q(\ram[108][12] ) );
  DFFHQX1 \ram_reg[108][11]  ( .D(n2321), .CK(clk), .Q(\ram[108][11] ) );
  DFFHQX1 \ram_reg[108][10]  ( .D(n2320), .CK(clk), .Q(\ram[108][10] ) );
  DFFHQX1 \ram_reg[108][9]  ( .D(n2319), .CK(clk), .Q(\ram[108][9] ) );
  DFFHQX1 \ram_reg[108][8]  ( .D(n2318), .CK(clk), .Q(\ram[108][8] ) );
  DFFHQX1 \ram_reg[108][7]  ( .D(n2317), .CK(clk), .Q(\ram[108][7] ) );
  DFFHQX1 \ram_reg[108][6]  ( .D(n2316), .CK(clk), .Q(\ram[108][6] ) );
  DFFHQX1 \ram_reg[108][5]  ( .D(n2315), .CK(clk), .Q(\ram[108][5] ) );
  DFFHQX1 \ram_reg[108][4]  ( .D(n2314), .CK(clk), .Q(\ram[108][4] ) );
  DFFHQX1 \ram_reg[108][3]  ( .D(n2313), .CK(clk), .Q(\ram[108][3] ) );
  DFFHQX1 \ram_reg[108][2]  ( .D(n2312), .CK(clk), .Q(\ram[108][2] ) );
  DFFHQX1 \ram_reg[108][1]  ( .D(n2311), .CK(clk), .Q(\ram[108][1] ) );
  DFFHQX1 \ram_reg[108][0]  ( .D(n2310), .CK(clk), .Q(\ram[108][0] ) );
  DFFHQX1 \ram_reg[104][15]  ( .D(n2261), .CK(clk), .Q(\ram[104][15] ) );
  DFFHQX1 \ram_reg[104][14]  ( .D(n2260), .CK(clk), .Q(\ram[104][14] ) );
  DFFHQX1 \ram_reg[104][13]  ( .D(n2259), .CK(clk), .Q(\ram[104][13] ) );
  DFFHQX1 \ram_reg[104][12]  ( .D(n2258), .CK(clk), .Q(\ram[104][12] ) );
  DFFHQX1 \ram_reg[104][11]  ( .D(n2257), .CK(clk), .Q(\ram[104][11] ) );
  DFFHQX1 \ram_reg[104][10]  ( .D(n2256), .CK(clk), .Q(\ram[104][10] ) );
  DFFHQX1 \ram_reg[104][9]  ( .D(n2255), .CK(clk), .Q(\ram[104][9] ) );
  DFFHQX1 \ram_reg[104][8]  ( .D(n2254), .CK(clk), .Q(\ram[104][8] ) );
  DFFHQX1 \ram_reg[104][7]  ( .D(n2253), .CK(clk), .Q(\ram[104][7] ) );
  DFFHQX1 \ram_reg[104][6]  ( .D(n2252), .CK(clk), .Q(\ram[104][6] ) );
  DFFHQX1 \ram_reg[104][5]  ( .D(n2251), .CK(clk), .Q(\ram[104][5] ) );
  DFFHQX1 \ram_reg[104][4]  ( .D(n2250), .CK(clk), .Q(\ram[104][4] ) );
  DFFHQX1 \ram_reg[104][3]  ( .D(n2249), .CK(clk), .Q(\ram[104][3] ) );
  DFFHQX1 \ram_reg[104][2]  ( .D(n2248), .CK(clk), .Q(\ram[104][2] ) );
  DFFHQX1 \ram_reg[104][1]  ( .D(n2247), .CK(clk), .Q(\ram[104][1] ) );
  DFFHQX1 \ram_reg[104][0]  ( .D(n2246), .CK(clk), .Q(\ram[104][0] ) );
  DFFHQX1 \ram_reg[100][15]  ( .D(n2197), .CK(clk), .Q(\ram[100][15] ) );
  DFFHQX1 \ram_reg[100][14]  ( .D(n2196), .CK(clk), .Q(\ram[100][14] ) );
  DFFHQX1 \ram_reg[100][13]  ( .D(n2195), .CK(clk), .Q(\ram[100][13] ) );
  DFFHQX1 \ram_reg[100][12]  ( .D(n2194), .CK(clk), .Q(\ram[100][12] ) );
  DFFHQX1 \ram_reg[100][11]  ( .D(n2193), .CK(clk), .Q(\ram[100][11] ) );
  DFFHQX1 \ram_reg[100][10]  ( .D(n2192), .CK(clk), .Q(\ram[100][10] ) );
  DFFHQX1 \ram_reg[100][9]  ( .D(n2191), .CK(clk), .Q(\ram[100][9] ) );
  DFFHQX1 \ram_reg[100][8]  ( .D(n2190), .CK(clk), .Q(\ram[100][8] ) );
  DFFHQX1 \ram_reg[100][7]  ( .D(n2189), .CK(clk), .Q(\ram[100][7] ) );
  DFFHQX1 \ram_reg[100][6]  ( .D(n2188), .CK(clk), .Q(\ram[100][6] ) );
  DFFHQX1 \ram_reg[100][5]  ( .D(n2187), .CK(clk), .Q(\ram[100][5] ) );
  DFFHQX1 \ram_reg[100][4]  ( .D(n2186), .CK(clk), .Q(\ram[100][4] ) );
  DFFHQX1 \ram_reg[100][3]  ( .D(n2185), .CK(clk), .Q(\ram[100][3] ) );
  DFFHQX1 \ram_reg[100][2]  ( .D(n2184), .CK(clk), .Q(\ram[100][2] ) );
  DFFHQX1 \ram_reg[100][1]  ( .D(n2183), .CK(clk), .Q(\ram[100][1] ) );
  DFFHQX1 \ram_reg[100][0]  ( .D(n2182), .CK(clk), .Q(\ram[100][0] ) );
  DFFHQX1 \ram_reg[96][15]  ( .D(n2133), .CK(clk), .Q(\ram[96][15] ) );
  DFFHQX1 \ram_reg[96][14]  ( .D(n2132), .CK(clk), .Q(\ram[96][14] ) );
  DFFHQX1 \ram_reg[96][13]  ( .D(n2131), .CK(clk), .Q(\ram[96][13] ) );
  DFFHQX1 \ram_reg[96][12]  ( .D(n2130), .CK(clk), .Q(\ram[96][12] ) );
  DFFHQX1 \ram_reg[96][11]  ( .D(n2129), .CK(clk), .Q(\ram[96][11] ) );
  DFFHQX1 \ram_reg[96][10]  ( .D(n2128), .CK(clk), .Q(\ram[96][10] ) );
  DFFHQX1 \ram_reg[96][9]  ( .D(n2127), .CK(clk), .Q(\ram[96][9] ) );
  DFFHQX1 \ram_reg[96][8]  ( .D(n2126), .CK(clk), .Q(\ram[96][8] ) );
  DFFHQX1 \ram_reg[96][7]  ( .D(n2125), .CK(clk), .Q(\ram[96][7] ) );
  DFFHQX1 \ram_reg[96][6]  ( .D(n2124), .CK(clk), .Q(\ram[96][6] ) );
  DFFHQX1 \ram_reg[96][5]  ( .D(n2123), .CK(clk), .Q(\ram[96][5] ) );
  DFFHQX1 \ram_reg[96][4]  ( .D(n2122), .CK(clk), .Q(\ram[96][4] ) );
  DFFHQX1 \ram_reg[96][3]  ( .D(n2121), .CK(clk), .Q(\ram[96][3] ) );
  DFFHQX1 \ram_reg[96][2]  ( .D(n2120), .CK(clk), .Q(\ram[96][2] ) );
  DFFHQX1 \ram_reg[96][1]  ( .D(n2119), .CK(clk), .Q(\ram[96][1] ) );
  DFFHQX1 \ram_reg[96][0]  ( .D(n2118), .CK(clk), .Q(\ram[96][0] ) );
  DFFHQX1 \ram_reg[92][15]  ( .D(n2069), .CK(clk), .Q(\ram[92][15] ) );
  DFFHQX1 \ram_reg[92][14]  ( .D(n2068), .CK(clk), .Q(\ram[92][14] ) );
  DFFHQX1 \ram_reg[92][13]  ( .D(n2067), .CK(clk), .Q(\ram[92][13] ) );
  DFFHQX1 \ram_reg[92][12]  ( .D(n2066), .CK(clk), .Q(\ram[92][12] ) );
  DFFHQX1 \ram_reg[92][11]  ( .D(n2065), .CK(clk), .Q(\ram[92][11] ) );
  DFFHQX1 \ram_reg[92][10]  ( .D(n2064), .CK(clk), .Q(\ram[92][10] ) );
  DFFHQX1 \ram_reg[92][9]  ( .D(n2063), .CK(clk), .Q(\ram[92][9] ) );
  DFFHQX1 \ram_reg[92][8]  ( .D(n2062), .CK(clk), .Q(\ram[92][8] ) );
  DFFHQX1 \ram_reg[92][7]  ( .D(n2061), .CK(clk), .Q(\ram[92][7] ) );
  DFFHQX1 \ram_reg[92][6]  ( .D(n2060), .CK(clk), .Q(\ram[92][6] ) );
  DFFHQX1 \ram_reg[92][5]  ( .D(n2059), .CK(clk), .Q(\ram[92][5] ) );
  DFFHQX1 \ram_reg[92][4]  ( .D(n2058), .CK(clk), .Q(\ram[92][4] ) );
  DFFHQX1 \ram_reg[92][3]  ( .D(n2057), .CK(clk), .Q(\ram[92][3] ) );
  DFFHQX1 \ram_reg[92][2]  ( .D(n2056), .CK(clk), .Q(\ram[92][2] ) );
  DFFHQX1 \ram_reg[92][1]  ( .D(n2055), .CK(clk), .Q(\ram[92][1] ) );
  DFFHQX1 \ram_reg[92][0]  ( .D(n2054), .CK(clk), .Q(\ram[92][0] ) );
  DFFHQX1 \ram_reg[88][15]  ( .D(n2005), .CK(clk), .Q(\ram[88][15] ) );
  DFFHQX1 \ram_reg[88][14]  ( .D(n2004), .CK(clk), .Q(\ram[88][14] ) );
  DFFHQX1 \ram_reg[88][13]  ( .D(n2003), .CK(clk), .Q(\ram[88][13] ) );
  DFFHQX1 \ram_reg[88][12]  ( .D(n2002), .CK(clk), .Q(\ram[88][12] ) );
  DFFHQX1 \ram_reg[88][11]  ( .D(n2001), .CK(clk), .Q(\ram[88][11] ) );
  DFFHQX1 \ram_reg[88][10]  ( .D(n2000), .CK(clk), .Q(\ram[88][10] ) );
  DFFHQX1 \ram_reg[88][9]  ( .D(n1999), .CK(clk), .Q(\ram[88][9] ) );
  DFFHQX1 \ram_reg[88][8]  ( .D(n1998), .CK(clk), .Q(\ram[88][8] ) );
  DFFHQX1 \ram_reg[88][7]  ( .D(n1997), .CK(clk), .Q(\ram[88][7] ) );
  DFFHQX1 \ram_reg[88][6]  ( .D(n1996), .CK(clk), .Q(\ram[88][6] ) );
  DFFHQX1 \ram_reg[88][5]  ( .D(n1995), .CK(clk), .Q(\ram[88][5] ) );
  DFFHQX1 \ram_reg[88][4]  ( .D(n1994), .CK(clk), .Q(\ram[88][4] ) );
  DFFHQX1 \ram_reg[88][3]  ( .D(n1993), .CK(clk), .Q(\ram[88][3] ) );
  DFFHQX1 \ram_reg[88][2]  ( .D(n1992), .CK(clk), .Q(\ram[88][2] ) );
  DFFHQX1 \ram_reg[88][1]  ( .D(n1991), .CK(clk), .Q(\ram[88][1] ) );
  DFFHQX1 \ram_reg[88][0]  ( .D(n1990), .CK(clk), .Q(\ram[88][0] ) );
  DFFHQX1 \ram_reg[84][15]  ( .D(n1941), .CK(clk), .Q(\ram[84][15] ) );
  DFFHQX1 \ram_reg[84][14]  ( .D(n1940), .CK(clk), .Q(\ram[84][14] ) );
  DFFHQX1 \ram_reg[84][13]  ( .D(n1939), .CK(clk), .Q(\ram[84][13] ) );
  DFFHQX1 \ram_reg[84][12]  ( .D(n1938), .CK(clk), .Q(\ram[84][12] ) );
  DFFHQX1 \ram_reg[84][11]  ( .D(n1937), .CK(clk), .Q(\ram[84][11] ) );
  DFFHQX1 \ram_reg[84][10]  ( .D(n1936), .CK(clk), .Q(\ram[84][10] ) );
  DFFHQX1 \ram_reg[84][9]  ( .D(n1935), .CK(clk), .Q(\ram[84][9] ) );
  DFFHQX1 \ram_reg[84][8]  ( .D(n1934), .CK(clk), .Q(\ram[84][8] ) );
  DFFHQX1 \ram_reg[84][7]  ( .D(n1933), .CK(clk), .Q(\ram[84][7] ) );
  DFFHQX1 \ram_reg[84][6]  ( .D(n1932), .CK(clk), .Q(\ram[84][6] ) );
  DFFHQX1 \ram_reg[84][5]  ( .D(n1931), .CK(clk), .Q(\ram[84][5] ) );
  DFFHQX1 \ram_reg[84][4]  ( .D(n1930), .CK(clk), .Q(\ram[84][4] ) );
  DFFHQX1 \ram_reg[84][3]  ( .D(n1929), .CK(clk), .Q(\ram[84][3] ) );
  DFFHQX1 \ram_reg[84][2]  ( .D(n1928), .CK(clk), .Q(\ram[84][2] ) );
  DFFHQX1 \ram_reg[84][1]  ( .D(n1927), .CK(clk), .Q(\ram[84][1] ) );
  DFFHQX1 \ram_reg[84][0]  ( .D(n1926), .CK(clk), .Q(\ram[84][0] ) );
  DFFHQX1 \ram_reg[80][15]  ( .D(n1877), .CK(clk), .Q(\ram[80][15] ) );
  DFFHQX1 \ram_reg[80][14]  ( .D(n1876), .CK(clk), .Q(\ram[80][14] ) );
  DFFHQX1 \ram_reg[80][13]  ( .D(n1875), .CK(clk), .Q(\ram[80][13] ) );
  DFFHQX1 \ram_reg[80][12]  ( .D(n1874), .CK(clk), .Q(\ram[80][12] ) );
  DFFHQX1 \ram_reg[80][11]  ( .D(n1873), .CK(clk), .Q(\ram[80][11] ) );
  DFFHQX1 \ram_reg[80][10]  ( .D(n1872), .CK(clk), .Q(\ram[80][10] ) );
  DFFHQX1 \ram_reg[80][9]  ( .D(n1871), .CK(clk), .Q(\ram[80][9] ) );
  DFFHQX1 \ram_reg[80][8]  ( .D(n1870), .CK(clk), .Q(\ram[80][8] ) );
  DFFHQX1 \ram_reg[80][7]  ( .D(n1869), .CK(clk), .Q(\ram[80][7] ) );
  DFFHQX1 \ram_reg[80][6]  ( .D(n1868), .CK(clk), .Q(\ram[80][6] ) );
  DFFHQX1 \ram_reg[80][5]  ( .D(n1867), .CK(clk), .Q(\ram[80][5] ) );
  DFFHQX1 \ram_reg[80][4]  ( .D(n1866), .CK(clk), .Q(\ram[80][4] ) );
  DFFHQX1 \ram_reg[80][3]  ( .D(n1865), .CK(clk), .Q(\ram[80][3] ) );
  DFFHQX1 \ram_reg[80][2]  ( .D(n1864), .CK(clk), .Q(\ram[80][2] ) );
  DFFHQX1 \ram_reg[80][1]  ( .D(n1863), .CK(clk), .Q(\ram[80][1] ) );
  DFFHQX1 \ram_reg[80][0]  ( .D(n1862), .CK(clk), .Q(\ram[80][0] ) );
  DFFHQX1 \ram_reg[76][15]  ( .D(n1813), .CK(clk), .Q(\ram[76][15] ) );
  DFFHQX1 \ram_reg[76][14]  ( .D(n1812), .CK(clk), .Q(\ram[76][14] ) );
  DFFHQX1 \ram_reg[76][13]  ( .D(n1811), .CK(clk), .Q(\ram[76][13] ) );
  DFFHQX1 \ram_reg[76][12]  ( .D(n1810), .CK(clk), .Q(\ram[76][12] ) );
  DFFHQX1 \ram_reg[76][11]  ( .D(n1809), .CK(clk), .Q(\ram[76][11] ) );
  DFFHQX1 \ram_reg[76][10]  ( .D(n1808), .CK(clk), .Q(\ram[76][10] ) );
  DFFHQX1 \ram_reg[76][9]  ( .D(n1807), .CK(clk), .Q(\ram[76][9] ) );
  DFFHQX1 \ram_reg[76][8]  ( .D(n1806), .CK(clk), .Q(\ram[76][8] ) );
  DFFHQX1 \ram_reg[76][7]  ( .D(n1805), .CK(clk), .Q(\ram[76][7] ) );
  DFFHQX1 \ram_reg[76][6]  ( .D(n1804), .CK(clk), .Q(\ram[76][6] ) );
  DFFHQX1 \ram_reg[76][5]  ( .D(n1803), .CK(clk), .Q(\ram[76][5] ) );
  DFFHQX1 \ram_reg[76][4]  ( .D(n1802), .CK(clk), .Q(\ram[76][4] ) );
  DFFHQX1 \ram_reg[76][3]  ( .D(n1801), .CK(clk), .Q(\ram[76][3] ) );
  DFFHQX1 \ram_reg[76][2]  ( .D(n1800), .CK(clk), .Q(\ram[76][2] ) );
  DFFHQX1 \ram_reg[76][1]  ( .D(n1799), .CK(clk), .Q(\ram[76][1] ) );
  DFFHQX1 \ram_reg[76][0]  ( .D(n1798), .CK(clk), .Q(\ram[76][0] ) );
  DFFHQX1 \ram_reg[72][15]  ( .D(n1749), .CK(clk), .Q(\ram[72][15] ) );
  DFFHQX1 \ram_reg[72][14]  ( .D(n1748), .CK(clk), .Q(\ram[72][14] ) );
  DFFHQX1 \ram_reg[72][13]  ( .D(n1747), .CK(clk), .Q(\ram[72][13] ) );
  DFFHQX1 \ram_reg[72][12]  ( .D(n1746), .CK(clk), .Q(\ram[72][12] ) );
  DFFHQX1 \ram_reg[72][11]  ( .D(n1745), .CK(clk), .Q(\ram[72][11] ) );
  DFFHQX1 \ram_reg[72][10]  ( .D(n1744), .CK(clk), .Q(\ram[72][10] ) );
  DFFHQX1 \ram_reg[72][9]  ( .D(n1743), .CK(clk), .Q(\ram[72][9] ) );
  DFFHQX1 \ram_reg[72][8]  ( .D(n1742), .CK(clk), .Q(\ram[72][8] ) );
  DFFHQX1 \ram_reg[72][7]  ( .D(n1741), .CK(clk), .Q(\ram[72][7] ) );
  DFFHQX1 \ram_reg[72][6]  ( .D(n1740), .CK(clk), .Q(\ram[72][6] ) );
  DFFHQX1 \ram_reg[72][5]  ( .D(n1739), .CK(clk), .Q(\ram[72][5] ) );
  DFFHQX1 \ram_reg[72][4]  ( .D(n1738), .CK(clk), .Q(\ram[72][4] ) );
  DFFHQX1 \ram_reg[72][3]  ( .D(n1737), .CK(clk), .Q(\ram[72][3] ) );
  DFFHQX1 \ram_reg[72][2]  ( .D(n1736), .CK(clk), .Q(\ram[72][2] ) );
  DFFHQX1 \ram_reg[72][1]  ( .D(n1735), .CK(clk), .Q(\ram[72][1] ) );
  DFFHQX1 \ram_reg[72][0]  ( .D(n1734), .CK(clk), .Q(\ram[72][0] ) );
  DFFHQX1 \ram_reg[68][15]  ( .D(n1685), .CK(clk), .Q(\ram[68][15] ) );
  DFFHQX1 \ram_reg[68][14]  ( .D(n1684), .CK(clk), .Q(\ram[68][14] ) );
  DFFHQX1 \ram_reg[68][13]  ( .D(n1683), .CK(clk), .Q(\ram[68][13] ) );
  DFFHQX1 \ram_reg[68][12]  ( .D(n1682), .CK(clk), .Q(\ram[68][12] ) );
  DFFHQX1 \ram_reg[68][11]  ( .D(n1681), .CK(clk), .Q(\ram[68][11] ) );
  DFFHQX1 \ram_reg[68][10]  ( .D(n1680), .CK(clk), .Q(\ram[68][10] ) );
  DFFHQX1 \ram_reg[68][9]  ( .D(n1679), .CK(clk), .Q(\ram[68][9] ) );
  DFFHQX1 \ram_reg[68][8]  ( .D(n1678), .CK(clk), .Q(\ram[68][8] ) );
  DFFHQX1 \ram_reg[68][7]  ( .D(n1677), .CK(clk), .Q(\ram[68][7] ) );
  DFFHQX1 \ram_reg[68][6]  ( .D(n1676), .CK(clk), .Q(\ram[68][6] ) );
  DFFHQX1 \ram_reg[68][5]  ( .D(n1675), .CK(clk), .Q(\ram[68][5] ) );
  DFFHQX1 \ram_reg[68][4]  ( .D(n1674), .CK(clk), .Q(\ram[68][4] ) );
  DFFHQX1 \ram_reg[68][3]  ( .D(n1673), .CK(clk), .Q(\ram[68][3] ) );
  DFFHQX1 \ram_reg[68][2]  ( .D(n1672), .CK(clk), .Q(\ram[68][2] ) );
  DFFHQX1 \ram_reg[68][1]  ( .D(n1671), .CK(clk), .Q(\ram[68][1] ) );
  DFFHQX1 \ram_reg[68][0]  ( .D(n1670), .CK(clk), .Q(\ram[68][0] ) );
  DFFHQX1 \ram_reg[64][15]  ( .D(n1621), .CK(clk), .Q(\ram[64][15] ) );
  DFFHQX1 \ram_reg[64][14]  ( .D(n1620), .CK(clk), .Q(\ram[64][14] ) );
  DFFHQX1 \ram_reg[64][13]  ( .D(n1619), .CK(clk), .Q(\ram[64][13] ) );
  DFFHQX1 \ram_reg[64][12]  ( .D(n1618), .CK(clk), .Q(\ram[64][12] ) );
  DFFHQX1 \ram_reg[64][11]  ( .D(n1617), .CK(clk), .Q(\ram[64][11] ) );
  DFFHQX1 \ram_reg[64][10]  ( .D(n1616), .CK(clk), .Q(\ram[64][10] ) );
  DFFHQX1 \ram_reg[64][9]  ( .D(n1615), .CK(clk), .Q(\ram[64][9] ) );
  DFFHQX1 \ram_reg[64][8]  ( .D(n1614), .CK(clk), .Q(\ram[64][8] ) );
  DFFHQX1 \ram_reg[64][7]  ( .D(n1613), .CK(clk), .Q(\ram[64][7] ) );
  DFFHQX1 \ram_reg[64][6]  ( .D(n1612), .CK(clk), .Q(\ram[64][6] ) );
  DFFHQX1 \ram_reg[64][5]  ( .D(n1611), .CK(clk), .Q(\ram[64][5] ) );
  DFFHQX1 \ram_reg[64][4]  ( .D(n1610), .CK(clk), .Q(\ram[64][4] ) );
  DFFHQX1 \ram_reg[64][3]  ( .D(n1609), .CK(clk), .Q(\ram[64][3] ) );
  DFFHQX1 \ram_reg[64][2]  ( .D(n1608), .CK(clk), .Q(\ram[64][2] ) );
  DFFHQX1 \ram_reg[64][1]  ( .D(n1607), .CK(clk), .Q(\ram[64][1] ) );
  DFFHQX1 \ram_reg[64][0]  ( .D(n1606), .CK(clk), .Q(\ram[64][0] ) );
  DFFHQX1 \ram_reg[60][15]  ( .D(n1557), .CK(clk), .Q(\ram[60][15] ) );
  DFFHQX1 \ram_reg[60][14]  ( .D(n1556), .CK(clk), .Q(\ram[60][14] ) );
  DFFHQX1 \ram_reg[60][13]  ( .D(n1555), .CK(clk), .Q(\ram[60][13] ) );
  DFFHQX1 \ram_reg[60][12]  ( .D(n1554), .CK(clk), .Q(\ram[60][12] ) );
  DFFHQX1 \ram_reg[60][11]  ( .D(n1553), .CK(clk), .Q(\ram[60][11] ) );
  DFFHQX1 \ram_reg[60][10]  ( .D(n1552), .CK(clk), .Q(\ram[60][10] ) );
  DFFHQX1 \ram_reg[60][9]  ( .D(n1551), .CK(clk), .Q(\ram[60][9] ) );
  DFFHQX1 \ram_reg[60][8]  ( .D(n1550), .CK(clk), .Q(\ram[60][8] ) );
  DFFHQX1 \ram_reg[60][7]  ( .D(n1549), .CK(clk), .Q(\ram[60][7] ) );
  DFFHQX1 \ram_reg[60][6]  ( .D(n1548), .CK(clk), .Q(\ram[60][6] ) );
  DFFHQX1 \ram_reg[60][5]  ( .D(n1547), .CK(clk), .Q(\ram[60][5] ) );
  DFFHQX1 \ram_reg[60][4]  ( .D(n1546), .CK(clk), .Q(\ram[60][4] ) );
  DFFHQX1 \ram_reg[60][3]  ( .D(n1545), .CK(clk), .Q(\ram[60][3] ) );
  DFFHQX1 \ram_reg[60][2]  ( .D(n1544), .CK(clk), .Q(\ram[60][2] ) );
  DFFHQX1 \ram_reg[60][1]  ( .D(n1543), .CK(clk), .Q(\ram[60][1] ) );
  DFFHQX1 \ram_reg[60][0]  ( .D(n1542), .CK(clk), .Q(\ram[60][0] ) );
  DFFHQX1 \ram_reg[56][15]  ( .D(n1493), .CK(clk), .Q(\ram[56][15] ) );
  DFFHQX1 \ram_reg[56][14]  ( .D(n1492), .CK(clk), .Q(\ram[56][14] ) );
  DFFHQX1 \ram_reg[56][13]  ( .D(n1491), .CK(clk), .Q(\ram[56][13] ) );
  DFFHQX1 \ram_reg[56][12]  ( .D(n1490), .CK(clk), .Q(\ram[56][12] ) );
  DFFHQX1 \ram_reg[56][11]  ( .D(n1489), .CK(clk), .Q(\ram[56][11] ) );
  DFFHQX1 \ram_reg[56][10]  ( .D(n1488), .CK(clk), .Q(\ram[56][10] ) );
  DFFHQX1 \ram_reg[56][9]  ( .D(n1487), .CK(clk), .Q(\ram[56][9] ) );
  DFFHQX1 \ram_reg[56][8]  ( .D(n1486), .CK(clk), .Q(\ram[56][8] ) );
  DFFHQX1 \ram_reg[56][7]  ( .D(n1485), .CK(clk), .Q(\ram[56][7] ) );
  DFFHQX1 \ram_reg[56][6]  ( .D(n1484), .CK(clk), .Q(\ram[56][6] ) );
  DFFHQX1 \ram_reg[56][5]  ( .D(n1483), .CK(clk), .Q(\ram[56][5] ) );
  DFFHQX1 \ram_reg[56][4]  ( .D(n1482), .CK(clk), .Q(\ram[56][4] ) );
  DFFHQX1 \ram_reg[56][3]  ( .D(n1481), .CK(clk), .Q(\ram[56][3] ) );
  DFFHQX1 \ram_reg[56][2]  ( .D(n1480), .CK(clk), .Q(\ram[56][2] ) );
  DFFHQX1 \ram_reg[56][1]  ( .D(n1479), .CK(clk), .Q(\ram[56][1] ) );
  DFFHQX1 \ram_reg[56][0]  ( .D(n1478), .CK(clk), .Q(\ram[56][0] ) );
  DFFHQX1 \ram_reg[52][15]  ( .D(n1429), .CK(clk), .Q(\ram[52][15] ) );
  DFFHQX1 \ram_reg[52][14]  ( .D(n1428), .CK(clk), .Q(\ram[52][14] ) );
  DFFHQX1 \ram_reg[52][13]  ( .D(n1427), .CK(clk), .Q(\ram[52][13] ) );
  DFFHQX1 \ram_reg[52][12]  ( .D(n1426), .CK(clk), .Q(\ram[52][12] ) );
  DFFHQX1 \ram_reg[52][11]  ( .D(n1425), .CK(clk), .Q(\ram[52][11] ) );
  DFFHQX1 \ram_reg[52][10]  ( .D(n1424), .CK(clk), .Q(\ram[52][10] ) );
  DFFHQX1 \ram_reg[52][9]  ( .D(n1423), .CK(clk), .Q(\ram[52][9] ) );
  DFFHQX1 \ram_reg[52][8]  ( .D(n1422), .CK(clk), .Q(\ram[52][8] ) );
  DFFHQX1 \ram_reg[52][7]  ( .D(n1421), .CK(clk), .Q(\ram[52][7] ) );
  DFFHQX1 \ram_reg[52][6]  ( .D(n1420), .CK(clk), .Q(\ram[52][6] ) );
  DFFHQX1 \ram_reg[52][5]  ( .D(n1419), .CK(clk), .Q(\ram[52][5] ) );
  DFFHQX1 \ram_reg[52][4]  ( .D(n1418), .CK(clk), .Q(\ram[52][4] ) );
  DFFHQX1 \ram_reg[52][3]  ( .D(n1417), .CK(clk), .Q(\ram[52][3] ) );
  DFFHQX1 \ram_reg[52][2]  ( .D(n1416), .CK(clk), .Q(\ram[52][2] ) );
  DFFHQX1 \ram_reg[52][1]  ( .D(n1415), .CK(clk), .Q(\ram[52][1] ) );
  DFFHQX1 \ram_reg[52][0]  ( .D(n1414), .CK(clk), .Q(\ram[52][0] ) );
  DFFHQX1 \ram_reg[48][15]  ( .D(n1365), .CK(clk), .Q(\ram[48][15] ) );
  DFFHQX1 \ram_reg[48][14]  ( .D(n1364), .CK(clk), .Q(\ram[48][14] ) );
  DFFHQX1 \ram_reg[48][13]  ( .D(n1363), .CK(clk), .Q(\ram[48][13] ) );
  DFFHQX1 \ram_reg[48][12]  ( .D(n1362), .CK(clk), .Q(\ram[48][12] ) );
  DFFHQX1 \ram_reg[48][11]  ( .D(n1361), .CK(clk), .Q(\ram[48][11] ) );
  DFFHQX1 \ram_reg[48][10]  ( .D(n1360), .CK(clk), .Q(\ram[48][10] ) );
  DFFHQX1 \ram_reg[48][9]  ( .D(n1359), .CK(clk), .Q(\ram[48][9] ) );
  DFFHQX1 \ram_reg[48][8]  ( .D(n1358), .CK(clk), .Q(\ram[48][8] ) );
  DFFHQX1 \ram_reg[48][7]  ( .D(n1357), .CK(clk), .Q(\ram[48][7] ) );
  DFFHQX1 \ram_reg[48][6]  ( .D(n1356), .CK(clk), .Q(\ram[48][6] ) );
  DFFHQX1 \ram_reg[48][5]  ( .D(n1355), .CK(clk), .Q(\ram[48][5] ) );
  DFFHQX1 \ram_reg[48][4]  ( .D(n1354), .CK(clk), .Q(\ram[48][4] ) );
  DFFHQX1 \ram_reg[48][3]  ( .D(n1353), .CK(clk), .Q(\ram[48][3] ) );
  DFFHQX1 \ram_reg[48][2]  ( .D(n1352), .CK(clk), .Q(\ram[48][2] ) );
  DFFHQX1 \ram_reg[48][1]  ( .D(n1351), .CK(clk), .Q(\ram[48][1] ) );
  DFFHQX1 \ram_reg[48][0]  ( .D(n1350), .CK(clk), .Q(\ram[48][0] ) );
  DFFHQX1 \ram_reg[44][15]  ( .D(n1301), .CK(clk), .Q(\ram[44][15] ) );
  DFFHQX1 \ram_reg[44][14]  ( .D(n1300), .CK(clk), .Q(\ram[44][14] ) );
  DFFHQX1 \ram_reg[44][13]  ( .D(n1299), .CK(clk), .Q(\ram[44][13] ) );
  DFFHQX1 \ram_reg[44][12]  ( .D(n1298), .CK(clk), .Q(\ram[44][12] ) );
  DFFHQX1 \ram_reg[44][11]  ( .D(n1297), .CK(clk), .Q(\ram[44][11] ) );
  DFFHQX1 \ram_reg[44][10]  ( .D(n1296), .CK(clk), .Q(\ram[44][10] ) );
  DFFHQX1 \ram_reg[44][9]  ( .D(n1295), .CK(clk), .Q(\ram[44][9] ) );
  DFFHQX1 \ram_reg[44][8]  ( .D(n1294), .CK(clk), .Q(\ram[44][8] ) );
  DFFHQX1 \ram_reg[44][7]  ( .D(n1293), .CK(clk), .Q(\ram[44][7] ) );
  DFFHQX1 \ram_reg[44][6]  ( .D(n1292), .CK(clk), .Q(\ram[44][6] ) );
  DFFHQX1 \ram_reg[44][5]  ( .D(n1291), .CK(clk), .Q(\ram[44][5] ) );
  DFFHQX1 \ram_reg[44][4]  ( .D(n1290), .CK(clk), .Q(\ram[44][4] ) );
  DFFHQX1 \ram_reg[44][3]  ( .D(n1289), .CK(clk), .Q(\ram[44][3] ) );
  DFFHQX1 \ram_reg[44][2]  ( .D(n1288), .CK(clk), .Q(\ram[44][2] ) );
  DFFHQX1 \ram_reg[44][1]  ( .D(n1287), .CK(clk), .Q(\ram[44][1] ) );
  DFFHQX1 \ram_reg[44][0]  ( .D(n1286), .CK(clk), .Q(\ram[44][0] ) );
  DFFHQX1 \ram_reg[40][15]  ( .D(n1237), .CK(clk), .Q(\ram[40][15] ) );
  DFFHQX1 \ram_reg[40][14]  ( .D(n1236), .CK(clk), .Q(\ram[40][14] ) );
  DFFHQX1 \ram_reg[40][13]  ( .D(n1235), .CK(clk), .Q(\ram[40][13] ) );
  DFFHQX1 \ram_reg[40][12]  ( .D(n1234), .CK(clk), .Q(\ram[40][12] ) );
  DFFHQX1 \ram_reg[40][11]  ( .D(n1233), .CK(clk), .Q(\ram[40][11] ) );
  DFFHQX1 \ram_reg[40][10]  ( .D(n1232), .CK(clk), .Q(\ram[40][10] ) );
  DFFHQX1 \ram_reg[40][9]  ( .D(n1231), .CK(clk), .Q(\ram[40][9] ) );
  DFFHQX1 \ram_reg[40][8]  ( .D(n1230), .CK(clk), .Q(\ram[40][8] ) );
  DFFHQX1 \ram_reg[40][7]  ( .D(n1229), .CK(clk), .Q(\ram[40][7] ) );
  DFFHQX1 \ram_reg[40][6]  ( .D(n1228), .CK(clk), .Q(\ram[40][6] ) );
  DFFHQX1 \ram_reg[40][5]  ( .D(n1227), .CK(clk), .Q(\ram[40][5] ) );
  DFFHQX1 \ram_reg[40][4]  ( .D(n1226), .CK(clk), .Q(\ram[40][4] ) );
  DFFHQX1 \ram_reg[40][3]  ( .D(n1225), .CK(clk), .Q(\ram[40][3] ) );
  DFFHQX1 \ram_reg[40][2]  ( .D(n1224), .CK(clk), .Q(\ram[40][2] ) );
  DFFHQX1 \ram_reg[40][1]  ( .D(n1223), .CK(clk), .Q(\ram[40][1] ) );
  DFFHQX1 \ram_reg[40][0]  ( .D(n1222), .CK(clk), .Q(\ram[40][0] ) );
  DFFHQX1 \ram_reg[36][15]  ( .D(n1173), .CK(clk), .Q(\ram[36][15] ) );
  DFFHQX1 \ram_reg[36][14]  ( .D(n1172), .CK(clk), .Q(\ram[36][14] ) );
  DFFHQX1 \ram_reg[36][13]  ( .D(n1171), .CK(clk), .Q(\ram[36][13] ) );
  DFFHQX1 \ram_reg[36][12]  ( .D(n1170), .CK(clk), .Q(\ram[36][12] ) );
  DFFHQX1 \ram_reg[36][11]  ( .D(n1169), .CK(clk), .Q(\ram[36][11] ) );
  DFFHQX1 \ram_reg[36][10]  ( .D(n1168), .CK(clk), .Q(\ram[36][10] ) );
  DFFHQX1 \ram_reg[36][9]  ( .D(n1167), .CK(clk), .Q(\ram[36][9] ) );
  DFFHQX1 \ram_reg[36][8]  ( .D(n1166), .CK(clk), .Q(\ram[36][8] ) );
  DFFHQX1 \ram_reg[36][7]  ( .D(n1165), .CK(clk), .Q(\ram[36][7] ) );
  DFFHQX1 \ram_reg[36][6]  ( .D(n1164), .CK(clk), .Q(\ram[36][6] ) );
  DFFHQX1 \ram_reg[36][5]  ( .D(n1163), .CK(clk), .Q(\ram[36][5] ) );
  DFFHQX1 \ram_reg[36][4]  ( .D(n1162), .CK(clk), .Q(\ram[36][4] ) );
  DFFHQX1 \ram_reg[36][3]  ( .D(n1161), .CK(clk), .Q(\ram[36][3] ) );
  DFFHQX1 \ram_reg[36][2]  ( .D(n1160), .CK(clk), .Q(\ram[36][2] ) );
  DFFHQX1 \ram_reg[36][1]  ( .D(n1159), .CK(clk), .Q(\ram[36][1] ) );
  DFFHQX1 \ram_reg[36][0]  ( .D(n1158), .CK(clk), .Q(\ram[36][0] ) );
  DFFHQX1 \ram_reg[32][15]  ( .D(n1109), .CK(clk), .Q(\ram[32][15] ) );
  DFFHQX1 \ram_reg[32][14]  ( .D(n1108), .CK(clk), .Q(\ram[32][14] ) );
  DFFHQX1 \ram_reg[32][13]  ( .D(n1107), .CK(clk), .Q(\ram[32][13] ) );
  DFFHQX1 \ram_reg[32][12]  ( .D(n1106), .CK(clk), .Q(\ram[32][12] ) );
  DFFHQX1 \ram_reg[32][11]  ( .D(n1105), .CK(clk), .Q(\ram[32][11] ) );
  DFFHQX1 \ram_reg[32][10]  ( .D(n1104), .CK(clk), .Q(\ram[32][10] ) );
  DFFHQX1 \ram_reg[32][9]  ( .D(n1103), .CK(clk), .Q(\ram[32][9] ) );
  DFFHQX1 \ram_reg[32][8]  ( .D(n1102), .CK(clk), .Q(\ram[32][8] ) );
  DFFHQX1 \ram_reg[32][7]  ( .D(n1101), .CK(clk), .Q(\ram[32][7] ) );
  DFFHQX1 \ram_reg[32][6]  ( .D(n1100), .CK(clk), .Q(\ram[32][6] ) );
  DFFHQX1 \ram_reg[32][5]  ( .D(n1099), .CK(clk), .Q(\ram[32][5] ) );
  DFFHQX1 \ram_reg[32][4]  ( .D(n1098), .CK(clk), .Q(\ram[32][4] ) );
  DFFHQX1 \ram_reg[32][3]  ( .D(n1097), .CK(clk), .Q(\ram[32][3] ) );
  DFFHQX1 \ram_reg[32][2]  ( .D(n1096), .CK(clk), .Q(\ram[32][2] ) );
  DFFHQX1 \ram_reg[32][1]  ( .D(n1095), .CK(clk), .Q(\ram[32][1] ) );
  DFFHQX1 \ram_reg[32][0]  ( .D(n1094), .CK(clk), .Q(\ram[32][0] ) );
  DFFHQX1 \ram_reg[28][15]  ( .D(n1045), .CK(clk), .Q(\ram[28][15] ) );
  DFFHQX1 \ram_reg[28][14]  ( .D(n1044), .CK(clk), .Q(\ram[28][14] ) );
  DFFHQX1 \ram_reg[28][13]  ( .D(n1043), .CK(clk), .Q(\ram[28][13] ) );
  DFFHQX1 \ram_reg[28][12]  ( .D(n1042), .CK(clk), .Q(\ram[28][12] ) );
  DFFHQX1 \ram_reg[28][11]  ( .D(n1041), .CK(clk), .Q(\ram[28][11] ) );
  DFFHQX1 \ram_reg[28][10]  ( .D(n1040), .CK(clk), .Q(\ram[28][10] ) );
  DFFHQX1 \ram_reg[28][9]  ( .D(n1039), .CK(clk), .Q(\ram[28][9] ) );
  DFFHQX1 \ram_reg[28][8]  ( .D(n1038), .CK(clk), .Q(\ram[28][8] ) );
  DFFHQX1 \ram_reg[28][7]  ( .D(n1037), .CK(clk), .Q(\ram[28][7] ) );
  DFFHQX1 \ram_reg[28][6]  ( .D(n1036), .CK(clk), .Q(\ram[28][6] ) );
  DFFHQX1 \ram_reg[28][5]  ( .D(n1035), .CK(clk), .Q(\ram[28][5] ) );
  DFFHQX1 \ram_reg[28][4]  ( .D(n1034), .CK(clk), .Q(\ram[28][4] ) );
  DFFHQX1 \ram_reg[28][3]  ( .D(n1033), .CK(clk), .Q(\ram[28][3] ) );
  DFFHQX1 \ram_reg[28][2]  ( .D(n1032), .CK(clk), .Q(\ram[28][2] ) );
  DFFHQX1 \ram_reg[28][1]  ( .D(n1031), .CK(clk), .Q(\ram[28][1] ) );
  DFFHQX1 \ram_reg[28][0]  ( .D(n1030), .CK(clk), .Q(\ram[28][0] ) );
  DFFHQX1 \ram_reg[24][15]  ( .D(n981), .CK(clk), .Q(\ram[24][15] ) );
  DFFHQX1 \ram_reg[24][14]  ( .D(n980), .CK(clk), .Q(\ram[24][14] ) );
  DFFHQX1 \ram_reg[24][13]  ( .D(n979), .CK(clk), .Q(\ram[24][13] ) );
  DFFHQX1 \ram_reg[24][12]  ( .D(n978), .CK(clk), .Q(\ram[24][12] ) );
  DFFHQX1 \ram_reg[24][11]  ( .D(n977), .CK(clk), .Q(\ram[24][11] ) );
  DFFHQX1 \ram_reg[24][10]  ( .D(n976), .CK(clk), .Q(\ram[24][10] ) );
  DFFHQX1 \ram_reg[24][9]  ( .D(n975), .CK(clk), .Q(\ram[24][9] ) );
  DFFHQX1 \ram_reg[24][8]  ( .D(n974), .CK(clk), .Q(\ram[24][8] ) );
  DFFHQX1 \ram_reg[24][7]  ( .D(n973), .CK(clk), .Q(\ram[24][7] ) );
  DFFHQX1 \ram_reg[24][6]  ( .D(n972), .CK(clk), .Q(\ram[24][6] ) );
  DFFHQX1 \ram_reg[24][5]  ( .D(n971), .CK(clk), .Q(\ram[24][5] ) );
  DFFHQX1 \ram_reg[24][4]  ( .D(n970), .CK(clk), .Q(\ram[24][4] ) );
  DFFHQX1 \ram_reg[24][3]  ( .D(n969), .CK(clk), .Q(\ram[24][3] ) );
  DFFHQX1 \ram_reg[24][2]  ( .D(n968), .CK(clk), .Q(\ram[24][2] ) );
  DFFHQX1 \ram_reg[24][1]  ( .D(n967), .CK(clk), .Q(\ram[24][1] ) );
  DFFHQX1 \ram_reg[24][0]  ( .D(n966), .CK(clk), .Q(\ram[24][0] ) );
  DFFHQX1 \ram_reg[20][15]  ( .D(n917), .CK(clk), .Q(\ram[20][15] ) );
  DFFHQX1 \ram_reg[20][14]  ( .D(n916), .CK(clk), .Q(\ram[20][14] ) );
  DFFHQX1 \ram_reg[20][13]  ( .D(n915), .CK(clk), .Q(\ram[20][13] ) );
  DFFHQX1 \ram_reg[20][12]  ( .D(n914), .CK(clk), .Q(\ram[20][12] ) );
  DFFHQX1 \ram_reg[20][11]  ( .D(n913), .CK(clk), .Q(\ram[20][11] ) );
  DFFHQX1 \ram_reg[20][10]  ( .D(n912), .CK(clk), .Q(\ram[20][10] ) );
  DFFHQX1 \ram_reg[20][9]  ( .D(n911), .CK(clk), .Q(\ram[20][9] ) );
  DFFHQX1 \ram_reg[20][8]  ( .D(n910), .CK(clk), .Q(\ram[20][8] ) );
  DFFHQX1 \ram_reg[20][7]  ( .D(n909), .CK(clk), .Q(\ram[20][7] ) );
  DFFHQX1 \ram_reg[20][6]  ( .D(n908), .CK(clk), .Q(\ram[20][6] ) );
  DFFHQX1 \ram_reg[20][5]  ( .D(n907), .CK(clk), .Q(\ram[20][5] ) );
  DFFHQX1 \ram_reg[20][4]  ( .D(n906), .CK(clk), .Q(\ram[20][4] ) );
  DFFHQX1 \ram_reg[20][3]  ( .D(n905), .CK(clk), .Q(\ram[20][3] ) );
  DFFHQX1 \ram_reg[20][2]  ( .D(n904), .CK(clk), .Q(\ram[20][2] ) );
  DFFHQX1 \ram_reg[20][1]  ( .D(n903), .CK(clk), .Q(\ram[20][1] ) );
  DFFHQX1 \ram_reg[20][0]  ( .D(n902), .CK(clk), .Q(\ram[20][0] ) );
  DFFHQX1 \ram_reg[16][15]  ( .D(n853), .CK(clk), .Q(\ram[16][15] ) );
  DFFHQX1 \ram_reg[16][14]  ( .D(n852), .CK(clk), .Q(\ram[16][14] ) );
  DFFHQX1 \ram_reg[16][13]  ( .D(n851), .CK(clk), .Q(\ram[16][13] ) );
  DFFHQX1 \ram_reg[16][12]  ( .D(n850), .CK(clk), .Q(\ram[16][12] ) );
  DFFHQX1 \ram_reg[16][11]  ( .D(n849), .CK(clk), .Q(\ram[16][11] ) );
  DFFHQX1 \ram_reg[16][10]  ( .D(n848), .CK(clk), .Q(\ram[16][10] ) );
  DFFHQX1 \ram_reg[16][9]  ( .D(n847), .CK(clk), .Q(\ram[16][9] ) );
  DFFHQX1 \ram_reg[16][8]  ( .D(n846), .CK(clk), .Q(\ram[16][8] ) );
  DFFHQX1 \ram_reg[16][7]  ( .D(n845), .CK(clk), .Q(\ram[16][7] ) );
  DFFHQX1 \ram_reg[16][6]  ( .D(n844), .CK(clk), .Q(\ram[16][6] ) );
  DFFHQX1 \ram_reg[16][5]  ( .D(n843), .CK(clk), .Q(\ram[16][5] ) );
  DFFHQX1 \ram_reg[16][4]  ( .D(n842), .CK(clk), .Q(\ram[16][4] ) );
  DFFHQX1 \ram_reg[16][3]  ( .D(n841), .CK(clk), .Q(\ram[16][3] ) );
  DFFHQX1 \ram_reg[16][2]  ( .D(n840), .CK(clk), .Q(\ram[16][2] ) );
  DFFHQX1 \ram_reg[16][1]  ( .D(n839), .CK(clk), .Q(\ram[16][1] ) );
  DFFHQX1 \ram_reg[16][0]  ( .D(n838), .CK(clk), .Q(\ram[16][0] ) );
  DFFHQX1 \ram_reg[12][15]  ( .D(n789), .CK(clk), .Q(\ram[12][15] ) );
  DFFHQX1 \ram_reg[12][14]  ( .D(n788), .CK(clk), .Q(\ram[12][14] ) );
  DFFHQX1 \ram_reg[12][13]  ( .D(n787), .CK(clk), .Q(\ram[12][13] ) );
  DFFHQX1 \ram_reg[12][12]  ( .D(n786), .CK(clk), .Q(\ram[12][12] ) );
  DFFHQX1 \ram_reg[12][11]  ( .D(n785), .CK(clk), .Q(\ram[12][11] ) );
  DFFHQX1 \ram_reg[12][10]  ( .D(n784), .CK(clk), .Q(\ram[12][10] ) );
  DFFHQX1 \ram_reg[12][9]  ( .D(n783), .CK(clk), .Q(\ram[12][9] ) );
  DFFHQX1 \ram_reg[12][8]  ( .D(n782), .CK(clk), .Q(\ram[12][8] ) );
  DFFHQX1 \ram_reg[12][7]  ( .D(n781), .CK(clk), .Q(\ram[12][7] ) );
  DFFHQX1 \ram_reg[12][6]  ( .D(n780), .CK(clk), .Q(\ram[12][6] ) );
  DFFHQX1 \ram_reg[12][5]  ( .D(n779), .CK(clk), .Q(\ram[12][5] ) );
  DFFHQX1 \ram_reg[12][4]  ( .D(n778), .CK(clk), .Q(\ram[12][4] ) );
  DFFHQX1 \ram_reg[12][3]  ( .D(n777), .CK(clk), .Q(\ram[12][3] ) );
  DFFHQX1 \ram_reg[12][2]  ( .D(n776), .CK(clk), .Q(\ram[12][2] ) );
  DFFHQX1 \ram_reg[12][1]  ( .D(n775), .CK(clk), .Q(\ram[12][1] ) );
  DFFHQX1 \ram_reg[12][0]  ( .D(n774), .CK(clk), .Q(\ram[12][0] ) );
  DFFHQX1 \ram_reg[8][15]  ( .D(n725), .CK(clk), .Q(\ram[8][15] ) );
  DFFHQX1 \ram_reg[8][14]  ( .D(n724), .CK(clk), .Q(\ram[8][14] ) );
  DFFHQX1 \ram_reg[8][13]  ( .D(n723), .CK(clk), .Q(\ram[8][13] ) );
  DFFHQX1 \ram_reg[8][12]  ( .D(n722), .CK(clk), .Q(\ram[8][12] ) );
  DFFHQX1 \ram_reg[8][11]  ( .D(n721), .CK(clk), .Q(\ram[8][11] ) );
  DFFHQX1 \ram_reg[8][10]  ( .D(n720), .CK(clk), .Q(\ram[8][10] ) );
  DFFHQX1 \ram_reg[8][9]  ( .D(n719), .CK(clk), .Q(\ram[8][9] ) );
  DFFHQX1 \ram_reg[8][8]  ( .D(n718), .CK(clk), .Q(\ram[8][8] ) );
  DFFHQX1 \ram_reg[8][7]  ( .D(n717), .CK(clk), .Q(\ram[8][7] ) );
  DFFHQX1 \ram_reg[8][6]  ( .D(n716), .CK(clk), .Q(\ram[8][6] ) );
  DFFHQX1 \ram_reg[8][5]  ( .D(n715), .CK(clk), .Q(\ram[8][5] ) );
  DFFHQX1 \ram_reg[8][4]  ( .D(n714), .CK(clk), .Q(\ram[8][4] ) );
  DFFHQX1 \ram_reg[8][3]  ( .D(n713), .CK(clk), .Q(\ram[8][3] ) );
  DFFHQX1 \ram_reg[8][2]  ( .D(n712), .CK(clk), .Q(\ram[8][2] ) );
  DFFHQX1 \ram_reg[8][1]  ( .D(n711), .CK(clk), .Q(\ram[8][1] ) );
  DFFHQX1 \ram_reg[8][0]  ( .D(n710), .CK(clk), .Q(\ram[8][0] ) );
  DFFHQX1 \ram_reg[4][15]  ( .D(n661), .CK(clk), .Q(\ram[4][15] ) );
  DFFHQX1 \ram_reg[4][14]  ( .D(n660), .CK(clk), .Q(\ram[4][14] ) );
  DFFHQX1 \ram_reg[4][13]  ( .D(n659), .CK(clk), .Q(\ram[4][13] ) );
  DFFHQX1 \ram_reg[4][12]  ( .D(n658), .CK(clk), .Q(\ram[4][12] ) );
  DFFHQX1 \ram_reg[4][11]  ( .D(n657), .CK(clk), .Q(\ram[4][11] ) );
  DFFHQX1 \ram_reg[4][10]  ( .D(n656), .CK(clk), .Q(\ram[4][10] ) );
  DFFHQX1 \ram_reg[4][9]  ( .D(n655), .CK(clk), .Q(\ram[4][9] ) );
  DFFHQX1 \ram_reg[4][8]  ( .D(n654), .CK(clk), .Q(\ram[4][8] ) );
  DFFHQX1 \ram_reg[4][7]  ( .D(n653), .CK(clk), .Q(\ram[4][7] ) );
  DFFHQX1 \ram_reg[4][6]  ( .D(n652), .CK(clk), .Q(\ram[4][6] ) );
  DFFHQX1 \ram_reg[4][5]  ( .D(n651), .CK(clk), .Q(\ram[4][5] ) );
  DFFHQX1 \ram_reg[4][4]  ( .D(n650), .CK(clk), .Q(\ram[4][4] ) );
  DFFHQX1 \ram_reg[4][3]  ( .D(n649), .CK(clk), .Q(\ram[4][3] ) );
  DFFHQX1 \ram_reg[4][2]  ( .D(n648), .CK(clk), .Q(\ram[4][2] ) );
  DFFHQX1 \ram_reg[4][1]  ( .D(n647), .CK(clk), .Q(\ram[4][1] ) );
  DFFHQX1 \ram_reg[4][0]  ( .D(n646), .CK(clk), .Q(\ram[4][0] ) );
  DFFHQX1 \ram_reg[0][15]  ( .D(n597), .CK(clk), .Q(\ram[0][15] ) );
  DFFHQX1 \ram_reg[0][14]  ( .D(n596), .CK(clk), .Q(\ram[0][14] ) );
  DFFHQX1 \ram_reg[0][13]  ( .D(n595), .CK(clk), .Q(\ram[0][13] ) );
  DFFHQX1 \ram_reg[0][12]  ( .D(n594), .CK(clk), .Q(\ram[0][12] ) );
  DFFHQX1 \ram_reg[0][11]  ( .D(n593), .CK(clk), .Q(\ram[0][11] ) );
  DFFHQX1 \ram_reg[0][10]  ( .D(n592), .CK(clk), .Q(\ram[0][10] ) );
  DFFHQX1 \ram_reg[0][9]  ( .D(n591), .CK(clk), .Q(\ram[0][9] ) );
  DFFHQX1 \ram_reg[0][8]  ( .D(n590), .CK(clk), .Q(\ram[0][8] ) );
  DFFHQX1 \ram_reg[0][7]  ( .D(n589), .CK(clk), .Q(\ram[0][7] ) );
  DFFHQX1 \ram_reg[0][6]  ( .D(n588), .CK(clk), .Q(\ram[0][6] ) );
  DFFHQX1 \ram_reg[0][5]  ( .D(n587), .CK(clk), .Q(\ram[0][5] ) );
  DFFHQX1 \ram_reg[0][4]  ( .D(n586), .CK(clk), .Q(\ram[0][4] ) );
  DFFHQX1 \ram_reg[0][3]  ( .D(n585), .CK(clk), .Q(\ram[0][3] ) );
  DFFHQX1 \ram_reg[0][2]  ( .D(n584), .CK(clk), .Q(\ram[0][2] ) );
  DFFHQX1 \ram_reg[0][1]  ( .D(n583), .CK(clk), .Q(\ram[0][1] ) );
  DFFHQX1 \ram_reg[0][0]  ( .D(n582), .CK(clk), .Q(\ram[0][0] ) );
  DFFHQX1 \ram_reg[254][15]  ( .D(n4661), .CK(clk), .Q(\ram[254][15] ) );
  DFFHQX1 \ram_reg[254][14]  ( .D(n4660), .CK(clk), .Q(\ram[254][14] ) );
  DFFHQX1 \ram_reg[254][13]  ( .D(n4659), .CK(clk), .Q(\ram[254][13] ) );
  DFFHQX1 \ram_reg[254][12]  ( .D(n4658), .CK(clk), .Q(\ram[254][12] ) );
  DFFHQX1 \ram_reg[254][11]  ( .D(n4657), .CK(clk), .Q(\ram[254][11] ) );
  DFFHQX1 \ram_reg[254][10]  ( .D(n4656), .CK(clk), .Q(\ram[254][10] ) );
  DFFHQX1 \ram_reg[254][9]  ( .D(n4655), .CK(clk), .Q(\ram[254][9] ) );
  DFFHQX1 \ram_reg[254][8]  ( .D(n4654), .CK(clk), .Q(\ram[254][8] ) );
  DFFHQX1 \ram_reg[254][7]  ( .D(n4653), .CK(clk), .Q(\ram[254][7] ) );
  DFFHQX1 \ram_reg[254][6]  ( .D(n4652), .CK(clk), .Q(\ram[254][6] ) );
  DFFHQX1 \ram_reg[254][5]  ( .D(n4651), .CK(clk), .Q(\ram[254][5] ) );
  DFFHQX1 \ram_reg[254][4]  ( .D(n4650), .CK(clk), .Q(\ram[254][4] ) );
  DFFHQX1 \ram_reg[254][3]  ( .D(n4649), .CK(clk), .Q(\ram[254][3] ) );
  DFFHQX1 \ram_reg[254][2]  ( .D(n4648), .CK(clk), .Q(\ram[254][2] ) );
  DFFHQX1 \ram_reg[254][1]  ( .D(n4647), .CK(clk), .Q(\ram[254][1] ) );
  DFFHQX1 \ram_reg[254][0]  ( .D(n4646), .CK(clk), .Q(\ram[254][0] ) );
  DFFHQX1 \ram_reg[250][15]  ( .D(n4597), .CK(clk), .Q(\ram[250][15] ) );
  DFFHQX1 \ram_reg[250][14]  ( .D(n4596), .CK(clk), .Q(\ram[250][14] ) );
  DFFHQX1 \ram_reg[250][13]  ( .D(n4595), .CK(clk), .Q(\ram[250][13] ) );
  DFFHQX1 \ram_reg[250][12]  ( .D(n4594), .CK(clk), .Q(\ram[250][12] ) );
  DFFHQX1 \ram_reg[250][11]  ( .D(n4593), .CK(clk), .Q(\ram[250][11] ) );
  DFFHQX1 \ram_reg[250][10]  ( .D(n4592), .CK(clk), .Q(\ram[250][10] ) );
  DFFHQX1 \ram_reg[250][9]  ( .D(n4591), .CK(clk), .Q(\ram[250][9] ) );
  DFFHQX1 \ram_reg[250][8]  ( .D(n4590), .CK(clk), .Q(\ram[250][8] ) );
  DFFHQX1 \ram_reg[250][7]  ( .D(n4589), .CK(clk), .Q(\ram[250][7] ) );
  DFFHQX1 \ram_reg[250][6]  ( .D(n4588), .CK(clk), .Q(\ram[250][6] ) );
  DFFHQX1 \ram_reg[250][5]  ( .D(n4587), .CK(clk), .Q(\ram[250][5] ) );
  DFFHQX1 \ram_reg[250][4]  ( .D(n4586), .CK(clk), .Q(\ram[250][4] ) );
  DFFHQX1 \ram_reg[250][3]  ( .D(n4585), .CK(clk), .Q(\ram[250][3] ) );
  DFFHQX1 \ram_reg[250][2]  ( .D(n4584), .CK(clk), .Q(\ram[250][2] ) );
  DFFHQX1 \ram_reg[250][1]  ( .D(n4583), .CK(clk), .Q(\ram[250][1] ) );
  DFFHQX1 \ram_reg[250][0]  ( .D(n4582), .CK(clk), .Q(\ram[250][0] ) );
  DFFHQX1 \ram_reg[246][15]  ( .D(n4533), .CK(clk), .Q(\ram[246][15] ) );
  DFFHQX1 \ram_reg[246][14]  ( .D(n4532), .CK(clk), .Q(\ram[246][14] ) );
  DFFHQX1 \ram_reg[246][13]  ( .D(n4531), .CK(clk), .Q(\ram[246][13] ) );
  DFFHQX1 \ram_reg[246][12]  ( .D(n4530), .CK(clk), .Q(\ram[246][12] ) );
  DFFHQX1 \ram_reg[246][11]  ( .D(n4529), .CK(clk), .Q(\ram[246][11] ) );
  DFFHQX1 \ram_reg[246][10]  ( .D(n4528), .CK(clk), .Q(\ram[246][10] ) );
  DFFHQX1 \ram_reg[246][9]  ( .D(n4527), .CK(clk), .Q(\ram[246][9] ) );
  DFFHQX1 \ram_reg[246][8]  ( .D(n4526), .CK(clk), .Q(\ram[246][8] ) );
  DFFHQX1 \ram_reg[246][7]  ( .D(n4525), .CK(clk), .Q(\ram[246][7] ) );
  DFFHQX1 \ram_reg[246][6]  ( .D(n4524), .CK(clk), .Q(\ram[246][6] ) );
  DFFHQX1 \ram_reg[246][5]  ( .D(n4523), .CK(clk), .Q(\ram[246][5] ) );
  DFFHQX1 \ram_reg[246][4]  ( .D(n4522), .CK(clk), .Q(\ram[246][4] ) );
  DFFHQX1 \ram_reg[246][3]  ( .D(n4521), .CK(clk), .Q(\ram[246][3] ) );
  DFFHQX1 \ram_reg[246][2]  ( .D(n4520), .CK(clk), .Q(\ram[246][2] ) );
  DFFHQX1 \ram_reg[246][1]  ( .D(n4519), .CK(clk), .Q(\ram[246][1] ) );
  DFFHQX1 \ram_reg[246][0]  ( .D(n4518), .CK(clk), .Q(\ram[246][0] ) );
  DFFHQX1 \ram_reg[242][15]  ( .D(n4469), .CK(clk), .Q(\ram[242][15] ) );
  DFFHQX1 \ram_reg[242][14]  ( .D(n4468), .CK(clk), .Q(\ram[242][14] ) );
  DFFHQX1 \ram_reg[242][13]  ( .D(n4467), .CK(clk), .Q(\ram[242][13] ) );
  DFFHQX1 \ram_reg[242][12]  ( .D(n4466), .CK(clk), .Q(\ram[242][12] ) );
  DFFHQX1 \ram_reg[242][11]  ( .D(n4465), .CK(clk), .Q(\ram[242][11] ) );
  DFFHQX1 \ram_reg[242][10]  ( .D(n4464), .CK(clk), .Q(\ram[242][10] ) );
  DFFHQX1 \ram_reg[242][9]  ( .D(n4463), .CK(clk), .Q(\ram[242][9] ) );
  DFFHQX1 \ram_reg[242][8]  ( .D(n4462), .CK(clk), .Q(\ram[242][8] ) );
  DFFHQX1 \ram_reg[242][7]  ( .D(n4461), .CK(clk), .Q(\ram[242][7] ) );
  DFFHQX1 \ram_reg[242][6]  ( .D(n4460), .CK(clk), .Q(\ram[242][6] ) );
  DFFHQX1 \ram_reg[242][5]  ( .D(n4459), .CK(clk), .Q(\ram[242][5] ) );
  DFFHQX1 \ram_reg[242][4]  ( .D(n4458), .CK(clk), .Q(\ram[242][4] ) );
  DFFHQX1 \ram_reg[242][3]  ( .D(n4457), .CK(clk), .Q(\ram[242][3] ) );
  DFFHQX1 \ram_reg[242][2]  ( .D(n4456), .CK(clk), .Q(\ram[242][2] ) );
  DFFHQX1 \ram_reg[242][1]  ( .D(n4455), .CK(clk), .Q(\ram[242][1] ) );
  DFFHQX1 \ram_reg[242][0]  ( .D(n4454), .CK(clk), .Q(\ram[242][0] ) );
  DFFHQX1 \ram_reg[238][15]  ( .D(n4405), .CK(clk), .Q(\ram[238][15] ) );
  DFFHQX1 \ram_reg[238][14]  ( .D(n4404), .CK(clk), .Q(\ram[238][14] ) );
  DFFHQX1 \ram_reg[238][13]  ( .D(n4403), .CK(clk), .Q(\ram[238][13] ) );
  DFFHQX1 \ram_reg[238][12]  ( .D(n4402), .CK(clk), .Q(\ram[238][12] ) );
  DFFHQX1 \ram_reg[238][11]  ( .D(n4401), .CK(clk), .Q(\ram[238][11] ) );
  DFFHQX1 \ram_reg[238][10]  ( .D(n4400), .CK(clk), .Q(\ram[238][10] ) );
  DFFHQX1 \ram_reg[238][9]  ( .D(n4399), .CK(clk), .Q(\ram[238][9] ) );
  DFFHQX1 \ram_reg[238][8]  ( .D(n4398), .CK(clk), .Q(\ram[238][8] ) );
  DFFHQX1 \ram_reg[238][7]  ( .D(n4397), .CK(clk), .Q(\ram[238][7] ) );
  DFFHQX1 \ram_reg[238][6]  ( .D(n4396), .CK(clk), .Q(\ram[238][6] ) );
  DFFHQX1 \ram_reg[238][5]  ( .D(n4395), .CK(clk), .Q(\ram[238][5] ) );
  DFFHQX1 \ram_reg[238][4]  ( .D(n4394), .CK(clk), .Q(\ram[238][4] ) );
  DFFHQX1 \ram_reg[238][3]  ( .D(n4393), .CK(clk), .Q(\ram[238][3] ) );
  DFFHQX1 \ram_reg[238][2]  ( .D(n4392), .CK(clk), .Q(\ram[238][2] ) );
  DFFHQX1 \ram_reg[238][1]  ( .D(n4391), .CK(clk), .Q(\ram[238][1] ) );
  DFFHQX1 \ram_reg[238][0]  ( .D(n4390), .CK(clk), .Q(\ram[238][0] ) );
  DFFHQX1 \ram_reg[234][15]  ( .D(n4341), .CK(clk), .Q(\ram[234][15] ) );
  DFFHQX1 \ram_reg[234][14]  ( .D(n4340), .CK(clk), .Q(\ram[234][14] ) );
  DFFHQX1 \ram_reg[234][13]  ( .D(n4339), .CK(clk), .Q(\ram[234][13] ) );
  DFFHQX1 \ram_reg[234][12]  ( .D(n4338), .CK(clk), .Q(\ram[234][12] ) );
  DFFHQX1 \ram_reg[234][11]  ( .D(n4337), .CK(clk), .Q(\ram[234][11] ) );
  DFFHQX1 \ram_reg[234][10]  ( .D(n4336), .CK(clk), .Q(\ram[234][10] ) );
  DFFHQX1 \ram_reg[234][9]  ( .D(n4335), .CK(clk), .Q(\ram[234][9] ) );
  DFFHQX1 \ram_reg[234][8]  ( .D(n4334), .CK(clk), .Q(\ram[234][8] ) );
  DFFHQX1 \ram_reg[234][7]  ( .D(n4333), .CK(clk), .Q(\ram[234][7] ) );
  DFFHQX1 \ram_reg[234][6]  ( .D(n4332), .CK(clk), .Q(\ram[234][6] ) );
  DFFHQX1 \ram_reg[234][5]  ( .D(n4331), .CK(clk), .Q(\ram[234][5] ) );
  DFFHQX1 \ram_reg[234][4]  ( .D(n4330), .CK(clk), .Q(\ram[234][4] ) );
  DFFHQX1 \ram_reg[234][3]  ( .D(n4329), .CK(clk), .Q(\ram[234][3] ) );
  DFFHQX1 \ram_reg[234][2]  ( .D(n4328), .CK(clk), .Q(\ram[234][2] ) );
  DFFHQX1 \ram_reg[234][1]  ( .D(n4327), .CK(clk), .Q(\ram[234][1] ) );
  DFFHQX1 \ram_reg[234][0]  ( .D(n4326), .CK(clk), .Q(\ram[234][0] ) );
  DFFHQX1 \ram_reg[230][15]  ( .D(n4277), .CK(clk), .Q(\ram[230][15] ) );
  DFFHQX1 \ram_reg[230][14]  ( .D(n4276), .CK(clk), .Q(\ram[230][14] ) );
  DFFHQX1 \ram_reg[230][13]  ( .D(n4275), .CK(clk), .Q(\ram[230][13] ) );
  DFFHQX1 \ram_reg[230][12]  ( .D(n4274), .CK(clk), .Q(\ram[230][12] ) );
  DFFHQX1 \ram_reg[230][11]  ( .D(n4273), .CK(clk), .Q(\ram[230][11] ) );
  DFFHQX1 \ram_reg[230][10]  ( .D(n4272), .CK(clk), .Q(\ram[230][10] ) );
  DFFHQX1 \ram_reg[230][9]  ( .D(n4271), .CK(clk), .Q(\ram[230][9] ) );
  DFFHQX1 \ram_reg[230][8]  ( .D(n4270), .CK(clk), .Q(\ram[230][8] ) );
  DFFHQX1 \ram_reg[230][7]  ( .D(n4269), .CK(clk), .Q(\ram[230][7] ) );
  DFFHQX1 \ram_reg[230][6]  ( .D(n4268), .CK(clk), .Q(\ram[230][6] ) );
  DFFHQX1 \ram_reg[230][5]  ( .D(n4267), .CK(clk), .Q(\ram[230][5] ) );
  DFFHQX1 \ram_reg[230][4]  ( .D(n4266), .CK(clk), .Q(\ram[230][4] ) );
  DFFHQX1 \ram_reg[230][3]  ( .D(n4265), .CK(clk), .Q(\ram[230][3] ) );
  DFFHQX1 \ram_reg[230][2]  ( .D(n4264), .CK(clk), .Q(\ram[230][2] ) );
  DFFHQX1 \ram_reg[230][1]  ( .D(n4263), .CK(clk), .Q(\ram[230][1] ) );
  DFFHQX1 \ram_reg[230][0]  ( .D(n4262), .CK(clk), .Q(\ram[230][0] ) );
  DFFHQX1 \ram_reg[226][15]  ( .D(n4213), .CK(clk), .Q(\ram[226][15] ) );
  DFFHQX1 \ram_reg[226][14]  ( .D(n4212), .CK(clk), .Q(\ram[226][14] ) );
  DFFHQX1 \ram_reg[226][13]  ( .D(n4211), .CK(clk), .Q(\ram[226][13] ) );
  DFFHQX1 \ram_reg[226][12]  ( .D(n4210), .CK(clk), .Q(\ram[226][12] ) );
  DFFHQX1 \ram_reg[226][11]  ( .D(n4209), .CK(clk), .Q(\ram[226][11] ) );
  DFFHQX1 \ram_reg[226][10]  ( .D(n4208), .CK(clk), .Q(\ram[226][10] ) );
  DFFHQX1 \ram_reg[226][9]  ( .D(n4207), .CK(clk), .Q(\ram[226][9] ) );
  DFFHQX1 \ram_reg[226][8]  ( .D(n4206), .CK(clk), .Q(\ram[226][8] ) );
  DFFHQX1 \ram_reg[226][7]  ( .D(n4205), .CK(clk), .Q(\ram[226][7] ) );
  DFFHQX1 \ram_reg[226][6]  ( .D(n4204), .CK(clk), .Q(\ram[226][6] ) );
  DFFHQX1 \ram_reg[226][5]  ( .D(n4203), .CK(clk), .Q(\ram[226][5] ) );
  DFFHQX1 \ram_reg[226][4]  ( .D(n4202), .CK(clk), .Q(\ram[226][4] ) );
  DFFHQX1 \ram_reg[226][3]  ( .D(n4201), .CK(clk), .Q(\ram[226][3] ) );
  DFFHQX1 \ram_reg[226][2]  ( .D(n4200), .CK(clk), .Q(\ram[226][2] ) );
  DFFHQX1 \ram_reg[226][1]  ( .D(n4199), .CK(clk), .Q(\ram[226][1] ) );
  DFFHQX1 \ram_reg[226][0]  ( .D(n4198), .CK(clk), .Q(\ram[226][0] ) );
  DFFHQX1 \ram_reg[222][15]  ( .D(n4149), .CK(clk), .Q(\ram[222][15] ) );
  DFFHQX1 \ram_reg[222][14]  ( .D(n4148), .CK(clk), .Q(\ram[222][14] ) );
  DFFHQX1 \ram_reg[222][13]  ( .D(n4147), .CK(clk), .Q(\ram[222][13] ) );
  DFFHQX1 \ram_reg[222][12]  ( .D(n4146), .CK(clk), .Q(\ram[222][12] ) );
  DFFHQX1 \ram_reg[222][11]  ( .D(n4145), .CK(clk), .Q(\ram[222][11] ) );
  DFFHQX1 \ram_reg[222][10]  ( .D(n4144), .CK(clk), .Q(\ram[222][10] ) );
  DFFHQX1 \ram_reg[222][9]  ( .D(n4143), .CK(clk), .Q(\ram[222][9] ) );
  DFFHQX1 \ram_reg[222][8]  ( .D(n4142), .CK(clk), .Q(\ram[222][8] ) );
  DFFHQX1 \ram_reg[222][7]  ( .D(n4141), .CK(clk), .Q(\ram[222][7] ) );
  DFFHQX1 \ram_reg[222][6]  ( .D(n4140), .CK(clk), .Q(\ram[222][6] ) );
  DFFHQX1 \ram_reg[222][5]  ( .D(n4139), .CK(clk), .Q(\ram[222][5] ) );
  DFFHQX1 \ram_reg[222][4]  ( .D(n4138), .CK(clk), .Q(\ram[222][4] ) );
  DFFHQX1 \ram_reg[222][3]  ( .D(n4137), .CK(clk), .Q(\ram[222][3] ) );
  DFFHQX1 \ram_reg[222][2]  ( .D(n4136), .CK(clk), .Q(\ram[222][2] ) );
  DFFHQX1 \ram_reg[222][1]  ( .D(n4135), .CK(clk), .Q(\ram[222][1] ) );
  DFFHQX1 \ram_reg[222][0]  ( .D(n4134), .CK(clk), .Q(\ram[222][0] ) );
  DFFHQX1 \ram_reg[218][15]  ( .D(n4085), .CK(clk), .Q(\ram[218][15] ) );
  DFFHQX1 \ram_reg[218][14]  ( .D(n4084), .CK(clk), .Q(\ram[218][14] ) );
  DFFHQX1 \ram_reg[218][13]  ( .D(n4083), .CK(clk), .Q(\ram[218][13] ) );
  DFFHQX1 \ram_reg[218][12]  ( .D(n4082), .CK(clk), .Q(\ram[218][12] ) );
  DFFHQX1 \ram_reg[218][11]  ( .D(n4081), .CK(clk), .Q(\ram[218][11] ) );
  DFFHQX1 \ram_reg[218][10]  ( .D(n4080), .CK(clk), .Q(\ram[218][10] ) );
  DFFHQX1 \ram_reg[218][9]  ( .D(n4079), .CK(clk), .Q(\ram[218][9] ) );
  DFFHQX1 \ram_reg[218][8]  ( .D(n4078), .CK(clk), .Q(\ram[218][8] ) );
  DFFHQX1 \ram_reg[218][7]  ( .D(n4077), .CK(clk), .Q(\ram[218][7] ) );
  DFFHQX1 \ram_reg[218][6]  ( .D(n4076), .CK(clk), .Q(\ram[218][6] ) );
  DFFHQX1 \ram_reg[218][5]  ( .D(n4075), .CK(clk), .Q(\ram[218][5] ) );
  DFFHQX1 \ram_reg[218][4]  ( .D(n4074), .CK(clk), .Q(\ram[218][4] ) );
  DFFHQX1 \ram_reg[218][3]  ( .D(n4073), .CK(clk), .Q(\ram[218][3] ) );
  DFFHQX1 \ram_reg[218][2]  ( .D(n4072), .CK(clk), .Q(\ram[218][2] ) );
  DFFHQX1 \ram_reg[218][1]  ( .D(n4071), .CK(clk), .Q(\ram[218][1] ) );
  DFFHQX1 \ram_reg[218][0]  ( .D(n4070), .CK(clk), .Q(\ram[218][0] ) );
  DFFHQX1 \ram_reg[214][15]  ( .D(n4021), .CK(clk), .Q(\ram[214][15] ) );
  DFFHQX1 \ram_reg[214][14]  ( .D(n4020), .CK(clk), .Q(\ram[214][14] ) );
  DFFHQX1 \ram_reg[214][13]  ( .D(n4019), .CK(clk), .Q(\ram[214][13] ) );
  DFFHQX1 \ram_reg[214][12]  ( .D(n4018), .CK(clk), .Q(\ram[214][12] ) );
  DFFHQX1 \ram_reg[214][11]  ( .D(n4017), .CK(clk), .Q(\ram[214][11] ) );
  DFFHQX1 \ram_reg[214][10]  ( .D(n4016), .CK(clk), .Q(\ram[214][10] ) );
  DFFHQX1 \ram_reg[214][9]  ( .D(n4015), .CK(clk), .Q(\ram[214][9] ) );
  DFFHQX1 \ram_reg[214][8]  ( .D(n4014), .CK(clk), .Q(\ram[214][8] ) );
  DFFHQX1 \ram_reg[214][7]  ( .D(n4013), .CK(clk), .Q(\ram[214][7] ) );
  DFFHQX1 \ram_reg[214][6]  ( .D(n4012), .CK(clk), .Q(\ram[214][6] ) );
  DFFHQX1 \ram_reg[214][5]  ( .D(n4011), .CK(clk), .Q(\ram[214][5] ) );
  DFFHQX1 \ram_reg[214][4]  ( .D(n4010), .CK(clk), .Q(\ram[214][4] ) );
  DFFHQX1 \ram_reg[214][3]  ( .D(n4009), .CK(clk), .Q(\ram[214][3] ) );
  DFFHQX1 \ram_reg[214][2]  ( .D(n4008), .CK(clk), .Q(\ram[214][2] ) );
  DFFHQX1 \ram_reg[214][1]  ( .D(n4007), .CK(clk), .Q(\ram[214][1] ) );
  DFFHQX1 \ram_reg[214][0]  ( .D(n4006), .CK(clk), .Q(\ram[214][0] ) );
  DFFHQX1 \ram_reg[210][15]  ( .D(n3957), .CK(clk), .Q(\ram[210][15] ) );
  DFFHQX1 \ram_reg[210][14]  ( .D(n3956), .CK(clk), .Q(\ram[210][14] ) );
  DFFHQX1 \ram_reg[210][13]  ( .D(n3955), .CK(clk), .Q(\ram[210][13] ) );
  DFFHQX1 \ram_reg[210][12]  ( .D(n3954), .CK(clk), .Q(\ram[210][12] ) );
  DFFHQX1 \ram_reg[210][11]  ( .D(n3953), .CK(clk), .Q(\ram[210][11] ) );
  DFFHQX1 \ram_reg[210][10]  ( .D(n3952), .CK(clk), .Q(\ram[210][10] ) );
  DFFHQX1 \ram_reg[210][9]  ( .D(n3951), .CK(clk), .Q(\ram[210][9] ) );
  DFFHQX1 \ram_reg[210][8]  ( .D(n3950), .CK(clk), .Q(\ram[210][8] ) );
  DFFHQX1 \ram_reg[210][7]  ( .D(n3949), .CK(clk), .Q(\ram[210][7] ) );
  DFFHQX1 \ram_reg[210][6]  ( .D(n3948), .CK(clk), .Q(\ram[210][6] ) );
  DFFHQX1 \ram_reg[210][5]  ( .D(n3947), .CK(clk), .Q(\ram[210][5] ) );
  DFFHQX1 \ram_reg[210][4]  ( .D(n3946), .CK(clk), .Q(\ram[210][4] ) );
  DFFHQX1 \ram_reg[210][3]  ( .D(n3945), .CK(clk), .Q(\ram[210][3] ) );
  DFFHQX1 \ram_reg[210][2]  ( .D(n3944), .CK(clk), .Q(\ram[210][2] ) );
  DFFHQX1 \ram_reg[210][1]  ( .D(n3943), .CK(clk), .Q(\ram[210][1] ) );
  DFFHQX1 \ram_reg[210][0]  ( .D(n3942), .CK(clk), .Q(\ram[210][0] ) );
  DFFHQX1 \ram_reg[206][15]  ( .D(n3893), .CK(clk), .Q(\ram[206][15] ) );
  DFFHQX1 \ram_reg[206][14]  ( .D(n3892), .CK(clk), .Q(\ram[206][14] ) );
  DFFHQX1 \ram_reg[206][13]  ( .D(n3891), .CK(clk), .Q(\ram[206][13] ) );
  DFFHQX1 \ram_reg[206][12]  ( .D(n3890), .CK(clk), .Q(\ram[206][12] ) );
  DFFHQX1 \ram_reg[206][11]  ( .D(n3889), .CK(clk), .Q(\ram[206][11] ) );
  DFFHQX1 \ram_reg[206][10]  ( .D(n3888), .CK(clk), .Q(\ram[206][10] ) );
  DFFHQX1 \ram_reg[206][9]  ( .D(n3887), .CK(clk), .Q(\ram[206][9] ) );
  DFFHQX1 \ram_reg[206][8]  ( .D(n3886), .CK(clk), .Q(\ram[206][8] ) );
  DFFHQX1 \ram_reg[206][7]  ( .D(n3885), .CK(clk), .Q(\ram[206][7] ) );
  DFFHQX1 \ram_reg[206][6]  ( .D(n3884), .CK(clk), .Q(\ram[206][6] ) );
  DFFHQX1 \ram_reg[206][5]  ( .D(n3883), .CK(clk), .Q(\ram[206][5] ) );
  DFFHQX1 \ram_reg[206][4]  ( .D(n3882), .CK(clk), .Q(\ram[206][4] ) );
  DFFHQX1 \ram_reg[206][3]  ( .D(n3881), .CK(clk), .Q(\ram[206][3] ) );
  DFFHQX1 \ram_reg[206][2]  ( .D(n3880), .CK(clk), .Q(\ram[206][2] ) );
  DFFHQX1 \ram_reg[206][1]  ( .D(n3879), .CK(clk), .Q(\ram[206][1] ) );
  DFFHQX1 \ram_reg[206][0]  ( .D(n3878), .CK(clk), .Q(\ram[206][0] ) );
  DFFHQX1 \ram_reg[202][15]  ( .D(n3829), .CK(clk), .Q(\ram[202][15] ) );
  DFFHQX1 \ram_reg[202][14]  ( .D(n3828), .CK(clk), .Q(\ram[202][14] ) );
  DFFHQX1 \ram_reg[202][13]  ( .D(n3827), .CK(clk), .Q(\ram[202][13] ) );
  DFFHQX1 \ram_reg[202][12]  ( .D(n3826), .CK(clk), .Q(\ram[202][12] ) );
  DFFHQX1 \ram_reg[202][11]  ( .D(n3825), .CK(clk), .Q(\ram[202][11] ) );
  DFFHQX1 \ram_reg[202][10]  ( .D(n3824), .CK(clk), .Q(\ram[202][10] ) );
  DFFHQX1 \ram_reg[202][9]  ( .D(n3823), .CK(clk), .Q(\ram[202][9] ) );
  DFFHQX1 \ram_reg[202][8]  ( .D(n3822), .CK(clk), .Q(\ram[202][8] ) );
  DFFHQX1 \ram_reg[202][7]  ( .D(n3821), .CK(clk), .Q(\ram[202][7] ) );
  DFFHQX1 \ram_reg[202][6]  ( .D(n3820), .CK(clk), .Q(\ram[202][6] ) );
  DFFHQX1 \ram_reg[202][5]  ( .D(n3819), .CK(clk), .Q(\ram[202][5] ) );
  DFFHQX1 \ram_reg[202][4]  ( .D(n3818), .CK(clk), .Q(\ram[202][4] ) );
  DFFHQX1 \ram_reg[202][3]  ( .D(n3817), .CK(clk), .Q(\ram[202][3] ) );
  DFFHQX1 \ram_reg[202][2]  ( .D(n3816), .CK(clk), .Q(\ram[202][2] ) );
  DFFHQX1 \ram_reg[202][1]  ( .D(n3815), .CK(clk), .Q(\ram[202][1] ) );
  DFFHQX1 \ram_reg[202][0]  ( .D(n3814), .CK(clk), .Q(\ram[202][0] ) );
  DFFHQX1 \ram_reg[198][15]  ( .D(n3765), .CK(clk), .Q(\ram[198][15] ) );
  DFFHQX1 \ram_reg[198][14]  ( .D(n3764), .CK(clk), .Q(\ram[198][14] ) );
  DFFHQX1 \ram_reg[198][13]  ( .D(n3763), .CK(clk), .Q(\ram[198][13] ) );
  DFFHQX1 \ram_reg[198][12]  ( .D(n3762), .CK(clk), .Q(\ram[198][12] ) );
  DFFHQX1 \ram_reg[198][11]  ( .D(n3761), .CK(clk), .Q(\ram[198][11] ) );
  DFFHQX1 \ram_reg[198][10]  ( .D(n3760), .CK(clk), .Q(\ram[198][10] ) );
  DFFHQX1 \ram_reg[198][9]  ( .D(n3759), .CK(clk), .Q(\ram[198][9] ) );
  DFFHQX1 \ram_reg[198][8]  ( .D(n3758), .CK(clk), .Q(\ram[198][8] ) );
  DFFHQX1 \ram_reg[198][7]  ( .D(n3757), .CK(clk), .Q(\ram[198][7] ) );
  DFFHQX1 \ram_reg[198][6]  ( .D(n3756), .CK(clk), .Q(\ram[198][6] ) );
  DFFHQX1 \ram_reg[198][5]  ( .D(n3755), .CK(clk), .Q(\ram[198][5] ) );
  DFFHQX1 \ram_reg[198][4]  ( .D(n3754), .CK(clk), .Q(\ram[198][4] ) );
  DFFHQX1 \ram_reg[198][3]  ( .D(n3753), .CK(clk), .Q(\ram[198][3] ) );
  DFFHQX1 \ram_reg[198][2]  ( .D(n3752), .CK(clk), .Q(\ram[198][2] ) );
  DFFHQX1 \ram_reg[198][1]  ( .D(n3751), .CK(clk), .Q(\ram[198][1] ) );
  DFFHQX1 \ram_reg[198][0]  ( .D(n3750), .CK(clk), .Q(\ram[198][0] ) );
  DFFHQX1 \ram_reg[194][15]  ( .D(n3701), .CK(clk), .Q(\ram[194][15] ) );
  DFFHQX1 \ram_reg[194][14]  ( .D(n3700), .CK(clk), .Q(\ram[194][14] ) );
  DFFHQX1 \ram_reg[194][13]  ( .D(n3699), .CK(clk), .Q(\ram[194][13] ) );
  DFFHQX1 \ram_reg[194][12]  ( .D(n3698), .CK(clk), .Q(\ram[194][12] ) );
  DFFHQX1 \ram_reg[194][11]  ( .D(n3697), .CK(clk), .Q(\ram[194][11] ) );
  DFFHQX1 \ram_reg[194][10]  ( .D(n3696), .CK(clk), .Q(\ram[194][10] ) );
  DFFHQX1 \ram_reg[194][9]  ( .D(n3695), .CK(clk), .Q(\ram[194][9] ) );
  DFFHQX1 \ram_reg[194][8]  ( .D(n3694), .CK(clk), .Q(\ram[194][8] ) );
  DFFHQX1 \ram_reg[194][7]  ( .D(n3693), .CK(clk), .Q(\ram[194][7] ) );
  DFFHQX1 \ram_reg[194][6]  ( .D(n3692), .CK(clk), .Q(\ram[194][6] ) );
  DFFHQX1 \ram_reg[194][5]  ( .D(n3691), .CK(clk), .Q(\ram[194][5] ) );
  DFFHQX1 \ram_reg[194][4]  ( .D(n3690), .CK(clk), .Q(\ram[194][4] ) );
  DFFHQX1 \ram_reg[194][3]  ( .D(n3689), .CK(clk), .Q(\ram[194][3] ) );
  DFFHQX1 \ram_reg[194][2]  ( .D(n3688), .CK(clk), .Q(\ram[194][2] ) );
  DFFHQX1 \ram_reg[194][1]  ( .D(n3687), .CK(clk), .Q(\ram[194][1] ) );
  DFFHQX1 \ram_reg[194][0]  ( .D(n3686), .CK(clk), .Q(\ram[194][0] ) );
  DFFHQX1 \ram_reg[190][15]  ( .D(n3637), .CK(clk), .Q(\ram[190][15] ) );
  DFFHQX1 \ram_reg[190][14]  ( .D(n3636), .CK(clk), .Q(\ram[190][14] ) );
  DFFHQX1 \ram_reg[190][13]  ( .D(n3635), .CK(clk), .Q(\ram[190][13] ) );
  DFFHQX1 \ram_reg[190][12]  ( .D(n3634), .CK(clk), .Q(\ram[190][12] ) );
  DFFHQX1 \ram_reg[190][11]  ( .D(n3633), .CK(clk), .Q(\ram[190][11] ) );
  DFFHQX1 \ram_reg[190][10]  ( .D(n3632), .CK(clk), .Q(\ram[190][10] ) );
  DFFHQX1 \ram_reg[190][9]  ( .D(n3631), .CK(clk), .Q(\ram[190][9] ) );
  DFFHQX1 \ram_reg[190][8]  ( .D(n3630), .CK(clk), .Q(\ram[190][8] ) );
  DFFHQX1 \ram_reg[190][7]  ( .D(n3629), .CK(clk), .Q(\ram[190][7] ) );
  DFFHQX1 \ram_reg[190][6]  ( .D(n3628), .CK(clk), .Q(\ram[190][6] ) );
  DFFHQX1 \ram_reg[190][5]  ( .D(n3627), .CK(clk), .Q(\ram[190][5] ) );
  DFFHQX1 \ram_reg[190][4]  ( .D(n3626), .CK(clk), .Q(\ram[190][4] ) );
  DFFHQX1 \ram_reg[190][3]  ( .D(n3625), .CK(clk), .Q(\ram[190][3] ) );
  DFFHQX1 \ram_reg[190][2]  ( .D(n3624), .CK(clk), .Q(\ram[190][2] ) );
  DFFHQX1 \ram_reg[190][1]  ( .D(n3623), .CK(clk), .Q(\ram[190][1] ) );
  DFFHQX1 \ram_reg[190][0]  ( .D(n3622), .CK(clk), .Q(\ram[190][0] ) );
  DFFHQX1 \ram_reg[186][15]  ( .D(n3573), .CK(clk), .Q(\ram[186][15] ) );
  DFFHQX1 \ram_reg[186][14]  ( .D(n3572), .CK(clk), .Q(\ram[186][14] ) );
  DFFHQX1 \ram_reg[186][13]  ( .D(n3571), .CK(clk), .Q(\ram[186][13] ) );
  DFFHQX1 \ram_reg[186][12]  ( .D(n3570), .CK(clk), .Q(\ram[186][12] ) );
  DFFHQX1 \ram_reg[186][11]  ( .D(n3569), .CK(clk), .Q(\ram[186][11] ) );
  DFFHQX1 \ram_reg[186][10]  ( .D(n3568), .CK(clk), .Q(\ram[186][10] ) );
  DFFHQX1 \ram_reg[186][9]  ( .D(n3567), .CK(clk), .Q(\ram[186][9] ) );
  DFFHQX1 \ram_reg[186][8]  ( .D(n3566), .CK(clk), .Q(\ram[186][8] ) );
  DFFHQX1 \ram_reg[186][7]  ( .D(n3565), .CK(clk), .Q(\ram[186][7] ) );
  DFFHQX1 \ram_reg[186][6]  ( .D(n3564), .CK(clk), .Q(\ram[186][6] ) );
  DFFHQX1 \ram_reg[186][5]  ( .D(n3563), .CK(clk), .Q(\ram[186][5] ) );
  DFFHQX1 \ram_reg[186][4]  ( .D(n3562), .CK(clk), .Q(\ram[186][4] ) );
  DFFHQX1 \ram_reg[186][3]  ( .D(n3561), .CK(clk), .Q(\ram[186][3] ) );
  DFFHQX1 \ram_reg[186][2]  ( .D(n3560), .CK(clk), .Q(\ram[186][2] ) );
  DFFHQX1 \ram_reg[186][1]  ( .D(n3559), .CK(clk), .Q(\ram[186][1] ) );
  DFFHQX1 \ram_reg[186][0]  ( .D(n3558), .CK(clk), .Q(\ram[186][0] ) );
  DFFHQX1 \ram_reg[182][15]  ( .D(n3509), .CK(clk), .Q(\ram[182][15] ) );
  DFFHQX1 \ram_reg[182][14]  ( .D(n3508), .CK(clk), .Q(\ram[182][14] ) );
  DFFHQX1 \ram_reg[182][13]  ( .D(n3507), .CK(clk), .Q(\ram[182][13] ) );
  DFFHQX1 \ram_reg[182][12]  ( .D(n3506), .CK(clk), .Q(\ram[182][12] ) );
  DFFHQX1 \ram_reg[182][11]  ( .D(n3505), .CK(clk), .Q(\ram[182][11] ) );
  DFFHQX1 \ram_reg[182][10]  ( .D(n3504), .CK(clk), .Q(\ram[182][10] ) );
  DFFHQX1 \ram_reg[182][9]  ( .D(n3503), .CK(clk), .Q(\ram[182][9] ) );
  DFFHQX1 \ram_reg[182][8]  ( .D(n3502), .CK(clk), .Q(\ram[182][8] ) );
  DFFHQX1 \ram_reg[182][7]  ( .D(n3501), .CK(clk), .Q(\ram[182][7] ) );
  DFFHQX1 \ram_reg[182][6]  ( .D(n3500), .CK(clk), .Q(\ram[182][6] ) );
  DFFHQX1 \ram_reg[182][5]  ( .D(n3499), .CK(clk), .Q(\ram[182][5] ) );
  DFFHQX1 \ram_reg[182][4]  ( .D(n3498), .CK(clk), .Q(\ram[182][4] ) );
  DFFHQX1 \ram_reg[182][3]  ( .D(n3497), .CK(clk), .Q(\ram[182][3] ) );
  DFFHQX1 \ram_reg[182][2]  ( .D(n3496), .CK(clk), .Q(\ram[182][2] ) );
  DFFHQX1 \ram_reg[182][1]  ( .D(n3495), .CK(clk), .Q(\ram[182][1] ) );
  DFFHQX1 \ram_reg[182][0]  ( .D(n3494), .CK(clk), .Q(\ram[182][0] ) );
  DFFHQX1 \ram_reg[178][15]  ( .D(n3445), .CK(clk), .Q(\ram[178][15] ) );
  DFFHQX1 \ram_reg[178][14]  ( .D(n3444), .CK(clk), .Q(\ram[178][14] ) );
  DFFHQX1 \ram_reg[178][13]  ( .D(n3443), .CK(clk), .Q(\ram[178][13] ) );
  DFFHQX1 \ram_reg[178][12]  ( .D(n3442), .CK(clk), .Q(\ram[178][12] ) );
  DFFHQX1 \ram_reg[178][11]  ( .D(n3441), .CK(clk), .Q(\ram[178][11] ) );
  DFFHQX1 \ram_reg[178][10]  ( .D(n3440), .CK(clk), .Q(\ram[178][10] ) );
  DFFHQX1 \ram_reg[178][9]  ( .D(n3439), .CK(clk), .Q(\ram[178][9] ) );
  DFFHQX1 \ram_reg[178][8]  ( .D(n3438), .CK(clk), .Q(\ram[178][8] ) );
  DFFHQX1 \ram_reg[178][7]  ( .D(n3437), .CK(clk), .Q(\ram[178][7] ) );
  DFFHQX1 \ram_reg[178][6]  ( .D(n3436), .CK(clk), .Q(\ram[178][6] ) );
  DFFHQX1 \ram_reg[178][5]  ( .D(n3435), .CK(clk), .Q(\ram[178][5] ) );
  DFFHQX1 \ram_reg[178][4]  ( .D(n3434), .CK(clk), .Q(\ram[178][4] ) );
  DFFHQX1 \ram_reg[178][3]  ( .D(n3433), .CK(clk), .Q(\ram[178][3] ) );
  DFFHQX1 \ram_reg[178][2]  ( .D(n3432), .CK(clk), .Q(\ram[178][2] ) );
  DFFHQX1 \ram_reg[178][1]  ( .D(n3431), .CK(clk), .Q(\ram[178][1] ) );
  DFFHQX1 \ram_reg[178][0]  ( .D(n3430), .CK(clk), .Q(\ram[178][0] ) );
  DFFHQX1 \ram_reg[174][15]  ( .D(n3381), .CK(clk), .Q(\ram[174][15] ) );
  DFFHQX1 \ram_reg[174][14]  ( .D(n3380), .CK(clk), .Q(\ram[174][14] ) );
  DFFHQX1 \ram_reg[174][13]  ( .D(n3379), .CK(clk), .Q(\ram[174][13] ) );
  DFFHQX1 \ram_reg[174][12]  ( .D(n3378), .CK(clk), .Q(\ram[174][12] ) );
  DFFHQX1 \ram_reg[174][11]  ( .D(n3377), .CK(clk), .Q(\ram[174][11] ) );
  DFFHQX1 \ram_reg[174][10]  ( .D(n3376), .CK(clk), .Q(\ram[174][10] ) );
  DFFHQX1 \ram_reg[174][9]  ( .D(n3375), .CK(clk), .Q(\ram[174][9] ) );
  DFFHQX1 \ram_reg[174][8]  ( .D(n3374), .CK(clk), .Q(\ram[174][8] ) );
  DFFHQX1 \ram_reg[174][7]  ( .D(n3373), .CK(clk), .Q(\ram[174][7] ) );
  DFFHQX1 \ram_reg[174][6]  ( .D(n3372), .CK(clk), .Q(\ram[174][6] ) );
  DFFHQX1 \ram_reg[174][5]  ( .D(n3371), .CK(clk), .Q(\ram[174][5] ) );
  DFFHQX1 \ram_reg[174][4]  ( .D(n3370), .CK(clk), .Q(\ram[174][4] ) );
  DFFHQX1 \ram_reg[174][3]  ( .D(n3369), .CK(clk), .Q(\ram[174][3] ) );
  DFFHQX1 \ram_reg[174][2]  ( .D(n3368), .CK(clk), .Q(\ram[174][2] ) );
  DFFHQX1 \ram_reg[174][1]  ( .D(n3367), .CK(clk), .Q(\ram[174][1] ) );
  DFFHQX1 \ram_reg[174][0]  ( .D(n3366), .CK(clk), .Q(\ram[174][0] ) );
  DFFHQX1 \ram_reg[170][15]  ( .D(n3317), .CK(clk), .Q(\ram[170][15] ) );
  DFFHQX1 \ram_reg[170][14]  ( .D(n3316), .CK(clk), .Q(\ram[170][14] ) );
  DFFHQX1 \ram_reg[170][13]  ( .D(n3315), .CK(clk), .Q(\ram[170][13] ) );
  DFFHQX1 \ram_reg[170][12]  ( .D(n3314), .CK(clk), .Q(\ram[170][12] ) );
  DFFHQX1 \ram_reg[170][11]  ( .D(n3313), .CK(clk), .Q(\ram[170][11] ) );
  DFFHQX1 \ram_reg[170][10]  ( .D(n3312), .CK(clk), .Q(\ram[170][10] ) );
  DFFHQX1 \ram_reg[170][9]  ( .D(n3311), .CK(clk), .Q(\ram[170][9] ) );
  DFFHQX1 \ram_reg[170][8]  ( .D(n3310), .CK(clk), .Q(\ram[170][8] ) );
  DFFHQX1 \ram_reg[170][7]  ( .D(n3309), .CK(clk), .Q(\ram[170][7] ) );
  DFFHQX1 \ram_reg[170][6]  ( .D(n3308), .CK(clk), .Q(\ram[170][6] ) );
  DFFHQX1 \ram_reg[170][5]  ( .D(n3307), .CK(clk), .Q(\ram[170][5] ) );
  DFFHQX1 \ram_reg[170][4]  ( .D(n3306), .CK(clk), .Q(\ram[170][4] ) );
  DFFHQX1 \ram_reg[170][3]  ( .D(n3305), .CK(clk), .Q(\ram[170][3] ) );
  DFFHQX1 \ram_reg[170][2]  ( .D(n3304), .CK(clk), .Q(\ram[170][2] ) );
  DFFHQX1 \ram_reg[170][1]  ( .D(n3303), .CK(clk), .Q(\ram[170][1] ) );
  DFFHQX1 \ram_reg[170][0]  ( .D(n3302), .CK(clk), .Q(\ram[170][0] ) );
  DFFHQX1 \ram_reg[166][15]  ( .D(n3253), .CK(clk), .Q(\ram[166][15] ) );
  DFFHQX1 \ram_reg[166][14]  ( .D(n3252), .CK(clk), .Q(\ram[166][14] ) );
  DFFHQX1 \ram_reg[166][13]  ( .D(n3251), .CK(clk), .Q(\ram[166][13] ) );
  DFFHQX1 \ram_reg[166][12]  ( .D(n3250), .CK(clk), .Q(\ram[166][12] ) );
  DFFHQX1 \ram_reg[166][11]  ( .D(n3249), .CK(clk), .Q(\ram[166][11] ) );
  DFFHQX1 \ram_reg[166][10]  ( .D(n3248), .CK(clk), .Q(\ram[166][10] ) );
  DFFHQX1 \ram_reg[166][9]  ( .D(n3247), .CK(clk), .Q(\ram[166][9] ) );
  DFFHQX1 \ram_reg[166][8]  ( .D(n3246), .CK(clk), .Q(\ram[166][8] ) );
  DFFHQX1 \ram_reg[166][7]  ( .D(n3245), .CK(clk), .Q(\ram[166][7] ) );
  DFFHQX1 \ram_reg[166][6]  ( .D(n3244), .CK(clk), .Q(\ram[166][6] ) );
  DFFHQX1 \ram_reg[166][5]  ( .D(n3243), .CK(clk), .Q(\ram[166][5] ) );
  DFFHQX1 \ram_reg[166][4]  ( .D(n3242), .CK(clk), .Q(\ram[166][4] ) );
  DFFHQX1 \ram_reg[166][3]  ( .D(n3241), .CK(clk), .Q(\ram[166][3] ) );
  DFFHQX1 \ram_reg[166][2]  ( .D(n3240), .CK(clk), .Q(\ram[166][2] ) );
  DFFHQX1 \ram_reg[166][1]  ( .D(n3239), .CK(clk), .Q(\ram[166][1] ) );
  DFFHQX1 \ram_reg[166][0]  ( .D(n3238), .CK(clk), .Q(\ram[166][0] ) );
  DFFHQX1 \ram_reg[162][15]  ( .D(n3189), .CK(clk), .Q(\ram[162][15] ) );
  DFFHQX1 \ram_reg[162][14]  ( .D(n3188), .CK(clk), .Q(\ram[162][14] ) );
  DFFHQX1 \ram_reg[162][13]  ( .D(n3187), .CK(clk), .Q(\ram[162][13] ) );
  DFFHQX1 \ram_reg[162][12]  ( .D(n3186), .CK(clk), .Q(\ram[162][12] ) );
  DFFHQX1 \ram_reg[162][11]  ( .D(n3185), .CK(clk), .Q(\ram[162][11] ) );
  DFFHQX1 \ram_reg[162][10]  ( .D(n3184), .CK(clk), .Q(\ram[162][10] ) );
  DFFHQX1 \ram_reg[162][9]  ( .D(n3183), .CK(clk), .Q(\ram[162][9] ) );
  DFFHQX1 \ram_reg[162][8]  ( .D(n3182), .CK(clk), .Q(\ram[162][8] ) );
  DFFHQX1 \ram_reg[162][7]  ( .D(n3181), .CK(clk), .Q(\ram[162][7] ) );
  DFFHQX1 \ram_reg[162][6]  ( .D(n3180), .CK(clk), .Q(\ram[162][6] ) );
  DFFHQX1 \ram_reg[162][5]  ( .D(n3179), .CK(clk), .Q(\ram[162][5] ) );
  DFFHQX1 \ram_reg[162][4]  ( .D(n3178), .CK(clk), .Q(\ram[162][4] ) );
  DFFHQX1 \ram_reg[162][3]  ( .D(n3177), .CK(clk), .Q(\ram[162][3] ) );
  DFFHQX1 \ram_reg[162][2]  ( .D(n3176), .CK(clk), .Q(\ram[162][2] ) );
  DFFHQX1 \ram_reg[162][1]  ( .D(n3175), .CK(clk), .Q(\ram[162][1] ) );
  DFFHQX1 \ram_reg[162][0]  ( .D(n3174), .CK(clk), .Q(\ram[162][0] ) );
  DFFHQX1 \ram_reg[158][15]  ( .D(n3125), .CK(clk), .Q(\ram[158][15] ) );
  DFFHQX1 \ram_reg[158][14]  ( .D(n3124), .CK(clk), .Q(\ram[158][14] ) );
  DFFHQX1 \ram_reg[158][13]  ( .D(n3123), .CK(clk), .Q(\ram[158][13] ) );
  DFFHQX1 \ram_reg[158][12]  ( .D(n3122), .CK(clk), .Q(\ram[158][12] ) );
  DFFHQX1 \ram_reg[158][11]  ( .D(n3121), .CK(clk), .Q(\ram[158][11] ) );
  DFFHQX1 \ram_reg[158][10]  ( .D(n3120), .CK(clk), .Q(\ram[158][10] ) );
  DFFHQX1 \ram_reg[158][9]  ( .D(n3119), .CK(clk), .Q(\ram[158][9] ) );
  DFFHQX1 \ram_reg[158][8]  ( .D(n3118), .CK(clk), .Q(\ram[158][8] ) );
  DFFHQX1 \ram_reg[158][7]  ( .D(n3117), .CK(clk), .Q(\ram[158][7] ) );
  DFFHQX1 \ram_reg[158][6]  ( .D(n3116), .CK(clk), .Q(\ram[158][6] ) );
  DFFHQX1 \ram_reg[158][5]  ( .D(n3115), .CK(clk), .Q(\ram[158][5] ) );
  DFFHQX1 \ram_reg[158][4]  ( .D(n3114), .CK(clk), .Q(\ram[158][4] ) );
  DFFHQX1 \ram_reg[158][3]  ( .D(n3113), .CK(clk), .Q(\ram[158][3] ) );
  DFFHQX1 \ram_reg[158][2]  ( .D(n3112), .CK(clk), .Q(\ram[158][2] ) );
  DFFHQX1 \ram_reg[158][1]  ( .D(n3111), .CK(clk), .Q(\ram[158][1] ) );
  DFFHQX1 \ram_reg[158][0]  ( .D(n3110), .CK(clk), .Q(\ram[158][0] ) );
  DFFHQX1 \ram_reg[154][15]  ( .D(n3061), .CK(clk), .Q(\ram[154][15] ) );
  DFFHQX1 \ram_reg[154][14]  ( .D(n3060), .CK(clk), .Q(\ram[154][14] ) );
  DFFHQX1 \ram_reg[154][13]  ( .D(n3059), .CK(clk), .Q(\ram[154][13] ) );
  DFFHQX1 \ram_reg[154][12]  ( .D(n3058), .CK(clk), .Q(\ram[154][12] ) );
  DFFHQX1 \ram_reg[154][11]  ( .D(n3057), .CK(clk), .Q(\ram[154][11] ) );
  DFFHQX1 \ram_reg[154][10]  ( .D(n3056), .CK(clk), .Q(\ram[154][10] ) );
  DFFHQX1 \ram_reg[154][9]  ( .D(n3055), .CK(clk), .Q(\ram[154][9] ) );
  DFFHQX1 \ram_reg[154][8]  ( .D(n3054), .CK(clk), .Q(\ram[154][8] ) );
  DFFHQX1 \ram_reg[154][7]  ( .D(n3053), .CK(clk), .Q(\ram[154][7] ) );
  DFFHQX1 \ram_reg[154][6]  ( .D(n3052), .CK(clk), .Q(\ram[154][6] ) );
  DFFHQX1 \ram_reg[154][5]  ( .D(n3051), .CK(clk), .Q(\ram[154][5] ) );
  DFFHQX1 \ram_reg[154][4]  ( .D(n3050), .CK(clk), .Q(\ram[154][4] ) );
  DFFHQX1 \ram_reg[154][3]  ( .D(n3049), .CK(clk), .Q(\ram[154][3] ) );
  DFFHQX1 \ram_reg[154][2]  ( .D(n3048), .CK(clk), .Q(\ram[154][2] ) );
  DFFHQX1 \ram_reg[154][1]  ( .D(n3047), .CK(clk), .Q(\ram[154][1] ) );
  DFFHQX1 \ram_reg[154][0]  ( .D(n3046), .CK(clk), .Q(\ram[154][0] ) );
  DFFHQX1 \ram_reg[150][15]  ( .D(n2997), .CK(clk), .Q(\ram[150][15] ) );
  DFFHQX1 \ram_reg[150][14]  ( .D(n2996), .CK(clk), .Q(\ram[150][14] ) );
  DFFHQX1 \ram_reg[150][13]  ( .D(n2995), .CK(clk), .Q(\ram[150][13] ) );
  DFFHQX1 \ram_reg[150][12]  ( .D(n2994), .CK(clk), .Q(\ram[150][12] ) );
  DFFHQX1 \ram_reg[150][11]  ( .D(n2993), .CK(clk), .Q(\ram[150][11] ) );
  DFFHQX1 \ram_reg[150][10]  ( .D(n2992), .CK(clk), .Q(\ram[150][10] ) );
  DFFHQX1 \ram_reg[150][9]  ( .D(n2991), .CK(clk), .Q(\ram[150][9] ) );
  DFFHQX1 \ram_reg[150][8]  ( .D(n2990), .CK(clk), .Q(\ram[150][8] ) );
  DFFHQX1 \ram_reg[150][7]  ( .D(n2989), .CK(clk), .Q(\ram[150][7] ) );
  DFFHQX1 \ram_reg[150][6]  ( .D(n2988), .CK(clk), .Q(\ram[150][6] ) );
  DFFHQX1 \ram_reg[150][5]  ( .D(n2987), .CK(clk), .Q(\ram[150][5] ) );
  DFFHQX1 \ram_reg[150][4]  ( .D(n2986), .CK(clk), .Q(\ram[150][4] ) );
  DFFHQX1 \ram_reg[150][3]  ( .D(n2985), .CK(clk), .Q(\ram[150][3] ) );
  DFFHQX1 \ram_reg[150][2]  ( .D(n2984), .CK(clk), .Q(\ram[150][2] ) );
  DFFHQX1 \ram_reg[150][1]  ( .D(n2983), .CK(clk), .Q(\ram[150][1] ) );
  DFFHQX1 \ram_reg[150][0]  ( .D(n2982), .CK(clk), .Q(\ram[150][0] ) );
  DFFHQX1 \ram_reg[146][15]  ( .D(n2933), .CK(clk), .Q(\ram[146][15] ) );
  DFFHQX1 \ram_reg[146][14]  ( .D(n2932), .CK(clk), .Q(\ram[146][14] ) );
  DFFHQX1 \ram_reg[146][13]  ( .D(n2931), .CK(clk), .Q(\ram[146][13] ) );
  DFFHQX1 \ram_reg[146][12]  ( .D(n2930), .CK(clk), .Q(\ram[146][12] ) );
  DFFHQX1 \ram_reg[146][11]  ( .D(n2929), .CK(clk), .Q(\ram[146][11] ) );
  DFFHQX1 \ram_reg[146][10]  ( .D(n2928), .CK(clk), .Q(\ram[146][10] ) );
  DFFHQX1 \ram_reg[146][9]  ( .D(n2927), .CK(clk), .Q(\ram[146][9] ) );
  DFFHQX1 \ram_reg[146][8]  ( .D(n2926), .CK(clk), .Q(\ram[146][8] ) );
  DFFHQX1 \ram_reg[146][7]  ( .D(n2925), .CK(clk), .Q(\ram[146][7] ) );
  DFFHQX1 \ram_reg[146][6]  ( .D(n2924), .CK(clk), .Q(\ram[146][6] ) );
  DFFHQX1 \ram_reg[146][5]  ( .D(n2923), .CK(clk), .Q(\ram[146][5] ) );
  DFFHQX1 \ram_reg[146][4]  ( .D(n2922), .CK(clk), .Q(\ram[146][4] ) );
  DFFHQX1 \ram_reg[146][3]  ( .D(n2921), .CK(clk), .Q(\ram[146][3] ) );
  DFFHQX1 \ram_reg[146][2]  ( .D(n2920), .CK(clk), .Q(\ram[146][2] ) );
  DFFHQX1 \ram_reg[146][1]  ( .D(n2919), .CK(clk), .Q(\ram[146][1] ) );
  DFFHQX1 \ram_reg[146][0]  ( .D(n2918), .CK(clk), .Q(\ram[146][0] ) );
  DFFHQX1 \ram_reg[142][15]  ( .D(n2869), .CK(clk), .Q(\ram[142][15] ) );
  DFFHQX1 \ram_reg[142][14]  ( .D(n2868), .CK(clk), .Q(\ram[142][14] ) );
  DFFHQX1 \ram_reg[142][13]  ( .D(n2867), .CK(clk), .Q(\ram[142][13] ) );
  DFFHQX1 \ram_reg[142][12]  ( .D(n2866), .CK(clk), .Q(\ram[142][12] ) );
  DFFHQX1 \ram_reg[142][11]  ( .D(n2865), .CK(clk), .Q(\ram[142][11] ) );
  DFFHQX1 \ram_reg[142][10]  ( .D(n2864), .CK(clk), .Q(\ram[142][10] ) );
  DFFHQX1 \ram_reg[142][9]  ( .D(n2863), .CK(clk), .Q(\ram[142][9] ) );
  DFFHQX1 \ram_reg[142][8]  ( .D(n2862), .CK(clk), .Q(\ram[142][8] ) );
  DFFHQX1 \ram_reg[142][7]  ( .D(n2861), .CK(clk), .Q(\ram[142][7] ) );
  DFFHQX1 \ram_reg[142][6]  ( .D(n2860), .CK(clk), .Q(\ram[142][6] ) );
  DFFHQX1 \ram_reg[142][5]  ( .D(n2859), .CK(clk), .Q(\ram[142][5] ) );
  DFFHQX1 \ram_reg[142][4]  ( .D(n2858), .CK(clk), .Q(\ram[142][4] ) );
  DFFHQX1 \ram_reg[142][3]  ( .D(n2857), .CK(clk), .Q(\ram[142][3] ) );
  DFFHQX1 \ram_reg[142][2]  ( .D(n2856), .CK(clk), .Q(\ram[142][2] ) );
  DFFHQX1 \ram_reg[142][1]  ( .D(n2855), .CK(clk), .Q(\ram[142][1] ) );
  DFFHQX1 \ram_reg[142][0]  ( .D(n2854), .CK(clk), .Q(\ram[142][0] ) );
  DFFHQX1 \ram_reg[138][15]  ( .D(n2805), .CK(clk), .Q(\ram[138][15] ) );
  DFFHQX1 \ram_reg[138][14]  ( .D(n2804), .CK(clk), .Q(\ram[138][14] ) );
  DFFHQX1 \ram_reg[138][13]  ( .D(n2803), .CK(clk), .Q(\ram[138][13] ) );
  DFFHQX1 \ram_reg[138][12]  ( .D(n2802), .CK(clk), .Q(\ram[138][12] ) );
  DFFHQX1 \ram_reg[138][11]  ( .D(n2801), .CK(clk), .Q(\ram[138][11] ) );
  DFFHQX1 \ram_reg[138][10]  ( .D(n2800), .CK(clk), .Q(\ram[138][10] ) );
  DFFHQX1 \ram_reg[138][9]  ( .D(n2799), .CK(clk), .Q(\ram[138][9] ) );
  DFFHQX1 \ram_reg[138][8]  ( .D(n2798), .CK(clk), .Q(\ram[138][8] ) );
  DFFHQX1 \ram_reg[138][7]  ( .D(n2797), .CK(clk), .Q(\ram[138][7] ) );
  DFFHQX1 \ram_reg[138][6]  ( .D(n2796), .CK(clk), .Q(\ram[138][6] ) );
  DFFHQX1 \ram_reg[138][5]  ( .D(n2795), .CK(clk), .Q(\ram[138][5] ) );
  DFFHQX1 \ram_reg[138][4]  ( .D(n2794), .CK(clk), .Q(\ram[138][4] ) );
  DFFHQX1 \ram_reg[138][3]  ( .D(n2793), .CK(clk), .Q(\ram[138][3] ) );
  DFFHQX1 \ram_reg[138][2]  ( .D(n2792), .CK(clk), .Q(\ram[138][2] ) );
  DFFHQX1 \ram_reg[138][1]  ( .D(n2791), .CK(clk), .Q(\ram[138][1] ) );
  DFFHQX1 \ram_reg[138][0]  ( .D(n2790), .CK(clk), .Q(\ram[138][0] ) );
  DFFHQX1 \ram_reg[134][15]  ( .D(n2741), .CK(clk), .Q(\ram[134][15] ) );
  DFFHQX1 \ram_reg[134][14]  ( .D(n2740), .CK(clk), .Q(\ram[134][14] ) );
  DFFHQX1 \ram_reg[134][13]  ( .D(n2739), .CK(clk), .Q(\ram[134][13] ) );
  DFFHQX1 \ram_reg[134][12]  ( .D(n2738), .CK(clk), .Q(\ram[134][12] ) );
  DFFHQX1 \ram_reg[134][11]  ( .D(n2737), .CK(clk), .Q(\ram[134][11] ) );
  DFFHQX1 \ram_reg[134][10]  ( .D(n2736), .CK(clk), .Q(\ram[134][10] ) );
  DFFHQX1 \ram_reg[134][9]  ( .D(n2735), .CK(clk), .Q(\ram[134][9] ) );
  DFFHQX1 \ram_reg[134][8]  ( .D(n2734), .CK(clk), .Q(\ram[134][8] ) );
  DFFHQX1 \ram_reg[134][7]  ( .D(n2733), .CK(clk), .Q(\ram[134][7] ) );
  DFFHQX1 \ram_reg[134][6]  ( .D(n2732), .CK(clk), .Q(\ram[134][6] ) );
  DFFHQX1 \ram_reg[134][5]  ( .D(n2731), .CK(clk), .Q(\ram[134][5] ) );
  DFFHQX1 \ram_reg[134][4]  ( .D(n2730), .CK(clk), .Q(\ram[134][4] ) );
  DFFHQX1 \ram_reg[134][3]  ( .D(n2729), .CK(clk), .Q(\ram[134][3] ) );
  DFFHQX1 \ram_reg[134][2]  ( .D(n2728), .CK(clk), .Q(\ram[134][2] ) );
  DFFHQX1 \ram_reg[134][1]  ( .D(n2727), .CK(clk), .Q(\ram[134][1] ) );
  DFFHQX1 \ram_reg[134][0]  ( .D(n2726), .CK(clk), .Q(\ram[134][0] ) );
  DFFHQX1 \ram_reg[130][15]  ( .D(n2677), .CK(clk), .Q(\ram[130][15] ) );
  DFFHQX1 \ram_reg[130][14]  ( .D(n2676), .CK(clk), .Q(\ram[130][14] ) );
  DFFHQX1 \ram_reg[130][13]  ( .D(n2675), .CK(clk), .Q(\ram[130][13] ) );
  DFFHQX1 \ram_reg[130][12]  ( .D(n2674), .CK(clk), .Q(\ram[130][12] ) );
  DFFHQX1 \ram_reg[130][11]  ( .D(n2673), .CK(clk), .Q(\ram[130][11] ) );
  DFFHQX1 \ram_reg[130][10]  ( .D(n2672), .CK(clk), .Q(\ram[130][10] ) );
  DFFHQX1 \ram_reg[130][9]  ( .D(n2671), .CK(clk), .Q(\ram[130][9] ) );
  DFFHQX1 \ram_reg[130][8]  ( .D(n2670), .CK(clk), .Q(\ram[130][8] ) );
  DFFHQX1 \ram_reg[130][7]  ( .D(n2669), .CK(clk), .Q(\ram[130][7] ) );
  DFFHQX1 \ram_reg[130][6]  ( .D(n2668), .CK(clk), .Q(\ram[130][6] ) );
  DFFHQX1 \ram_reg[130][5]  ( .D(n2667), .CK(clk), .Q(\ram[130][5] ) );
  DFFHQX1 \ram_reg[130][4]  ( .D(n2666), .CK(clk), .Q(\ram[130][4] ) );
  DFFHQX1 \ram_reg[130][3]  ( .D(n2665), .CK(clk), .Q(\ram[130][3] ) );
  DFFHQX1 \ram_reg[130][2]  ( .D(n2664), .CK(clk), .Q(\ram[130][2] ) );
  DFFHQX1 \ram_reg[130][1]  ( .D(n2663), .CK(clk), .Q(\ram[130][1] ) );
  DFFHQX1 \ram_reg[130][0]  ( .D(n2662), .CK(clk), .Q(\ram[130][0] ) );
  DFFHQX1 \ram_reg[126][15]  ( .D(n2613), .CK(clk), .Q(\ram[126][15] ) );
  DFFHQX1 \ram_reg[126][14]  ( .D(n2612), .CK(clk), .Q(\ram[126][14] ) );
  DFFHQX1 \ram_reg[126][13]  ( .D(n2611), .CK(clk), .Q(\ram[126][13] ) );
  DFFHQX1 \ram_reg[126][12]  ( .D(n2610), .CK(clk), .Q(\ram[126][12] ) );
  DFFHQX1 \ram_reg[126][11]  ( .D(n2609), .CK(clk), .Q(\ram[126][11] ) );
  DFFHQX1 \ram_reg[126][10]  ( .D(n2608), .CK(clk), .Q(\ram[126][10] ) );
  DFFHQX1 \ram_reg[126][9]  ( .D(n2607), .CK(clk), .Q(\ram[126][9] ) );
  DFFHQX1 \ram_reg[126][8]  ( .D(n2606), .CK(clk), .Q(\ram[126][8] ) );
  DFFHQX1 \ram_reg[126][7]  ( .D(n2605), .CK(clk), .Q(\ram[126][7] ) );
  DFFHQX1 \ram_reg[126][6]  ( .D(n2604), .CK(clk), .Q(\ram[126][6] ) );
  DFFHQX1 \ram_reg[126][5]  ( .D(n2603), .CK(clk), .Q(\ram[126][5] ) );
  DFFHQX1 \ram_reg[126][4]  ( .D(n2602), .CK(clk), .Q(\ram[126][4] ) );
  DFFHQX1 \ram_reg[126][3]  ( .D(n2601), .CK(clk), .Q(\ram[126][3] ) );
  DFFHQX1 \ram_reg[126][2]  ( .D(n2600), .CK(clk), .Q(\ram[126][2] ) );
  DFFHQX1 \ram_reg[126][1]  ( .D(n2599), .CK(clk), .Q(\ram[126][1] ) );
  DFFHQX1 \ram_reg[126][0]  ( .D(n2598), .CK(clk), .Q(\ram[126][0] ) );
  DFFHQX1 \ram_reg[122][15]  ( .D(n2549), .CK(clk), .Q(\ram[122][15] ) );
  DFFHQX1 \ram_reg[122][14]  ( .D(n2548), .CK(clk), .Q(\ram[122][14] ) );
  DFFHQX1 \ram_reg[122][13]  ( .D(n2547), .CK(clk), .Q(\ram[122][13] ) );
  DFFHQX1 \ram_reg[122][12]  ( .D(n2546), .CK(clk), .Q(\ram[122][12] ) );
  DFFHQX1 \ram_reg[122][11]  ( .D(n2545), .CK(clk), .Q(\ram[122][11] ) );
  DFFHQX1 \ram_reg[122][10]  ( .D(n2544), .CK(clk), .Q(\ram[122][10] ) );
  DFFHQX1 \ram_reg[122][9]  ( .D(n2543), .CK(clk), .Q(\ram[122][9] ) );
  DFFHQX1 \ram_reg[122][8]  ( .D(n2542), .CK(clk), .Q(\ram[122][8] ) );
  DFFHQX1 \ram_reg[122][7]  ( .D(n2541), .CK(clk), .Q(\ram[122][7] ) );
  DFFHQX1 \ram_reg[122][6]  ( .D(n2540), .CK(clk), .Q(\ram[122][6] ) );
  DFFHQX1 \ram_reg[122][5]  ( .D(n2539), .CK(clk), .Q(\ram[122][5] ) );
  DFFHQX1 \ram_reg[122][4]  ( .D(n2538), .CK(clk), .Q(\ram[122][4] ) );
  DFFHQX1 \ram_reg[122][3]  ( .D(n2537), .CK(clk), .Q(\ram[122][3] ) );
  DFFHQX1 \ram_reg[122][2]  ( .D(n2536), .CK(clk), .Q(\ram[122][2] ) );
  DFFHQX1 \ram_reg[122][1]  ( .D(n2535), .CK(clk), .Q(\ram[122][1] ) );
  DFFHQX1 \ram_reg[122][0]  ( .D(n2534), .CK(clk), .Q(\ram[122][0] ) );
  DFFHQX1 \ram_reg[118][15]  ( .D(n2485), .CK(clk), .Q(\ram[118][15] ) );
  DFFHQX1 \ram_reg[118][14]  ( .D(n2484), .CK(clk), .Q(\ram[118][14] ) );
  DFFHQX1 \ram_reg[118][13]  ( .D(n2483), .CK(clk), .Q(\ram[118][13] ) );
  DFFHQX1 \ram_reg[118][12]  ( .D(n2482), .CK(clk), .Q(\ram[118][12] ) );
  DFFHQX1 \ram_reg[118][11]  ( .D(n2481), .CK(clk), .Q(\ram[118][11] ) );
  DFFHQX1 \ram_reg[118][10]  ( .D(n2480), .CK(clk), .Q(\ram[118][10] ) );
  DFFHQX1 \ram_reg[118][9]  ( .D(n2479), .CK(clk), .Q(\ram[118][9] ) );
  DFFHQX1 \ram_reg[118][8]  ( .D(n2478), .CK(clk), .Q(\ram[118][8] ) );
  DFFHQX1 \ram_reg[118][7]  ( .D(n2477), .CK(clk), .Q(\ram[118][7] ) );
  DFFHQX1 \ram_reg[118][6]  ( .D(n2476), .CK(clk), .Q(\ram[118][6] ) );
  DFFHQX1 \ram_reg[118][5]  ( .D(n2475), .CK(clk), .Q(\ram[118][5] ) );
  DFFHQX1 \ram_reg[118][4]  ( .D(n2474), .CK(clk), .Q(\ram[118][4] ) );
  DFFHQX1 \ram_reg[118][3]  ( .D(n2473), .CK(clk), .Q(\ram[118][3] ) );
  DFFHQX1 \ram_reg[118][2]  ( .D(n2472), .CK(clk), .Q(\ram[118][2] ) );
  DFFHQX1 \ram_reg[118][1]  ( .D(n2471), .CK(clk), .Q(\ram[118][1] ) );
  DFFHQX1 \ram_reg[118][0]  ( .D(n2470), .CK(clk), .Q(\ram[118][0] ) );
  DFFHQX1 \ram_reg[114][15]  ( .D(n2421), .CK(clk), .Q(\ram[114][15] ) );
  DFFHQX1 \ram_reg[114][14]  ( .D(n2420), .CK(clk), .Q(\ram[114][14] ) );
  DFFHQX1 \ram_reg[114][13]  ( .D(n2419), .CK(clk), .Q(\ram[114][13] ) );
  DFFHQX1 \ram_reg[114][12]  ( .D(n2418), .CK(clk), .Q(\ram[114][12] ) );
  DFFHQX1 \ram_reg[114][11]  ( .D(n2417), .CK(clk), .Q(\ram[114][11] ) );
  DFFHQX1 \ram_reg[114][10]  ( .D(n2416), .CK(clk), .Q(\ram[114][10] ) );
  DFFHQX1 \ram_reg[114][9]  ( .D(n2415), .CK(clk), .Q(\ram[114][9] ) );
  DFFHQX1 \ram_reg[114][8]  ( .D(n2414), .CK(clk), .Q(\ram[114][8] ) );
  DFFHQX1 \ram_reg[114][7]  ( .D(n2413), .CK(clk), .Q(\ram[114][7] ) );
  DFFHQX1 \ram_reg[114][6]  ( .D(n2412), .CK(clk), .Q(\ram[114][6] ) );
  DFFHQX1 \ram_reg[114][5]  ( .D(n2411), .CK(clk), .Q(\ram[114][5] ) );
  DFFHQX1 \ram_reg[114][4]  ( .D(n2410), .CK(clk), .Q(\ram[114][4] ) );
  DFFHQX1 \ram_reg[114][3]  ( .D(n2409), .CK(clk), .Q(\ram[114][3] ) );
  DFFHQX1 \ram_reg[114][2]  ( .D(n2408), .CK(clk), .Q(\ram[114][2] ) );
  DFFHQX1 \ram_reg[114][1]  ( .D(n2407), .CK(clk), .Q(\ram[114][1] ) );
  DFFHQX1 \ram_reg[114][0]  ( .D(n2406), .CK(clk), .Q(\ram[114][0] ) );
  DFFHQX1 \ram_reg[110][15]  ( .D(n2357), .CK(clk), .Q(\ram[110][15] ) );
  DFFHQX1 \ram_reg[110][14]  ( .D(n2356), .CK(clk), .Q(\ram[110][14] ) );
  DFFHQX1 \ram_reg[110][13]  ( .D(n2355), .CK(clk), .Q(\ram[110][13] ) );
  DFFHQX1 \ram_reg[110][12]  ( .D(n2354), .CK(clk), .Q(\ram[110][12] ) );
  DFFHQX1 \ram_reg[110][11]  ( .D(n2353), .CK(clk), .Q(\ram[110][11] ) );
  DFFHQX1 \ram_reg[110][10]  ( .D(n2352), .CK(clk), .Q(\ram[110][10] ) );
  DFFHQX1 \ram_reg[110][9]  ( .D(n2351), .CK(clk), .Q(\ram[110][9] ) );
  DFFHQX1 \ram_reg[110][8]  ( .D(n2350), .CK(clk), .Q(\ram[110][8] ) );
  DFFHQX1 \ram_reg[110][7]  ( .D(n2349), .CK(clk), .Q(\ram[110][7] ) );
  DFFHQX1 \ram_reg[110][6]  ( .D(n2348), .CK(clk), .Q(\ram[110][6] ) );
  DFFHQX1 \ram_reg[110][5]  ( .D(n2347), .CK(clk), .Q(\ram[110][5] ) );
  DFFHQX1 \ram_reg[110][4]  ( .D(n2346), .CK(clk), .Q(\ram[110][4] ) );
  DFFHQX1 \ram_reg[110][3]  ( .D(n2345), .CK(clk), .Q(\ram[110][3] ) );
  DFFHQX1 \ram_reg[110][2]  ( .D(n2344), .CK(clk), .Q(\ram[110][2] ) );
  DFFHQX1 \ram_reg[110][1]  ( .D(n2343), .CK(clk), .Q(\ram[110][1] ) );
  DFFHQX1 \ram_reg[110][0]  ( .D(n2342), .CK(clk), .Q(\ram[110][0] ) );
  DFFHQX1 \ram_reg[106][15]  ( .D(n2293), .CK(clk), .Q(\ram[106][15] ) );
  DFFHQX1 \ram_reg[106][14]  ( .D(n2292), .CK(clk), .Q(\ram[106][14] ) );
  DFFHQX1 \ram_reg[106][13]  ( .D(n2291), .CK(clk), .Q(\ram[106][13] ) );
  DFFHQX1 \ram_reg[106][12]  ( .D(n2290), .CK(clk), .Q(\ram[106][12] ) );
  DFFHQX1 \ram_reg[106][11]  ( .D(n2289), .CK(clk), .Q(\ram[106][11] ) );
  DFFHQX1 \ram_reg[106][10]  ( .D(n2288), .CK(clk), .Q(\ram[106][10] ) );
  DFFHQX1 \ram_reg[106][9]  ( .D(n2287), .CK(clk), .Q(\ram[106][9] ) );
  DFFHQX1 \ram_reg[106][8]  ( .D(n2286), .CK(clk), .Q(\ram[106][8] ) );
  DFFHQX1 \ram_reg[106][7]  ( .D(n2285), .CK(clk), .Q(\ram[106][7] ) );
  DFFHQX1 \ram_reg[106][6]  ( .D(n2284), .CK(clk), .Q(\ram[106][6] ) );
  DFFHQX1 \ram_reg[106][5]  ( .D(n2283), .CK(clk), .Q(\ram[106][5] ) );
  DFFHQX1 \ram_reg[106][4]  ( .D(n2282), .CK(clk), .Q(\ram[106][4] ) );
  DFFHQX1 \ram_reg[106][3]  ( .D(n2281), .CK(clk), .Q(\ram[106][3] ) );
  DFFHQX1 \ram_reg[106][2]  ( .D(n2280), .CK(clk), .Q(\ram[106][2] ) );
  DFFHQX1 \ram_reg[106][1]  ( .D(n2279), .CK(clk), .Q(\ram[106][1] ) );
  DFFHQX1 \ram_reg[106][0]  ( .D(n2278), .CK(clk), .Q(\ram[106][0] ) );
  DFFHQX1 \ram_reg[102][15]  ( .D(n2229), .CK(clk), .Q(\ram[102][15] ) );
  DFFHQX1 \ram_reg[102][14]  ( .D(n2228), .CK(clk), .Q(\ram[102][14] ) );
  DFFHQX1 \ram_reg[102][13]  ( .D(n2227), .CK(clk), .Q(\ram[102][13] ) );
  DFFHQX1 \ram_reg[102][12]  ( .D(n2226), .CK(clk), .Q(\ram[102][12] ) );
  DFFHQX1 \ram_reg[102][11]  ( .D(n2225), .CK(clk), .Q(\ram[102][11] ) );
  DFFHQX1 \ram_reg[102][10]  ( .D(n2224), .CK(clk), .Q(\ram[102][10] ) );
  DFFHQX1 \ram_reg[102][9]  ( .D(n2223), .CK(clk), .Q(\ram[102][9] ) );
  DFFHQX1 \ram_reg[102][8]  ( .D(n2222), .CK(clk), .Q(\ram[102][8] ) );
  DFFHQX1 \ram_reg[102][7]  ( .D(n2221), .CK(clk), .Q(\ram[102][7] ) );
  DFFHQX1 \ram_reg[102][6]  ( .D(n2220), .CK(clk), .Q(\ram[102][6] ) );
  DFFHQX1 \ram_reg[102][5]  ( .D(n2219), .CK(clk), .Q(\ram[102][5] ) );
  DFFHQX1 \ram_reg[102][4]  ( .D(n2218), .CK(clk), .Q(\ram[102][4] ) );
  DFFHQX1 \ram_reg[102][3]  ( .D(n2217), .CK(clk), .Q(\ram[102][3] ) );
  DFFHQX1 \ram_reg[102][2]  ( .D(n2216), .CK(clk), .Q(\ram[102][2] ) );
  DFFHQX1 \ram_reg[102][1]  ( .D(n2215), .CK(clk), .Q(\ram[102][1] ) );
  DFFHQX1 \ram_reg[102][0]  ( .D(n2214), .CK(clk), .Q(\ram[102][0] ) );
  DFFHQX1 \ram_reg[98][15]  ( .D(n2165), .CK(clk), .Q(\ram[98][15] ) );
  DFFHQX1 \ram_reg[98][14]  ( .D(n2164), .CK(clk), .Q(\ram[98][14] ) );
  DFFHQX1 \ram_reg[98][13]  ( .D(n2163), .CK(clk), .Q(\ram[98][13] ) );
  DFFHQX1 \ram_reg[98][12]  ( .D(n2162), .CK(clk), .Q(\ram[98][12] ) );
  DFFHQX1 \ram_reg[98][11]  ( .D(n2161), .CK(clk), .Q(\ram[98][11] ) );
  DFFHQX1 \ram_reg[98][10]  ( .D(n2160), .CK(clk), .Q(\ram[98][10] ) );
  DFFHQX1 \ram_reg[98][9]  ( .D(n2159), .CK(clk), .Q(\ram[98][9] ) );
  DFFHQX1 \ram_reg[98][8]  ( .D(n2158), .CK(clk), .Q(\ram[98][8] ) );
  DFFHQX1 \ram_reg[98][7]  ( .D(n2157), .CK(clk), .Q(\ram[98][7] ) );
  DFFHQX1 \ram_reg[98][6]  ( .D(n2156), .CK(clk), .Q(\ram[98][6] ) );
  DFFHQX1 \ram_reg[98][5]  ( .D(n2155), .CK(clk), .Q(\ram[98][5] ) );
  DFFHQX1 \ram_reg[98][4]  ( .D(n2154), .CK(clk), .Q(\ram[98][4] ) );
  DFFHQX1 \ram_reg[98][3]  ( .D(n2153), .CK(clk), .Q(\ram[98][3] ) );
  DFFHQX1 \ram_reg[98][2]  ( .D(n2152), .CK(clk), .Q(\ram[98][2] ) );
  DFFHQX1 \ram_reg[98][1]  ( .D(n2151), .CK(clk), .Q(\ram[98][1] ) );
  DFFHQX1 \ram_reg[98][0]  ( .D(n2150), .CK(clk), .Q(\ram[98][0] ) );
  DFFHQX1 \ram_reg[94][15]  ( .D(n2101), .CK(clk), .Q(\ram[94][15] ) );
  DFFHQX1 \ram_reg[94][14]  ( .D(n2100), .CK(clk), .Q(\ram[94][14] ) );
  DFFHQX1 \ram_reg[94][13]  ( .D(n2099), .CK(clk), .Q(\ram[94][13] ) );
  DFFHQX1 \ram_reg[94][12]  ( .D(n2098), .CK(clk), .Q(\ram[94][12] ) );
  DFFHQX1 \ram_reg[94][11]  ( .D(n2097), .CK(clk), .Q(\ram[94][11] ) );
  DFFHQX1 \ram_reg[94][10]  ( .D(n2096), .CK(clk), .Q(\ram[94][10] ) );
  DFFHQX1 \ram_reg[94][9]  ( .D(n2095), .CK(clk), .Q(\ram[94][9] ) );
  DFFHQX1 \ram_reg[94][8]  ( .D(n2094), .CK(clk), .Q(\ram[94][8] ) );
  DFFHQX1 \ram_reg[94][7]  ( .D(n2093), .CK(clk), .Q(\ram[94][7] ) );
  DFFHQX1 \ram_reg[94][6]  ( .D(n2092), .CK(clk), .Q(\ram[94][6] ) );
  DFFHQX1 \ram_reg[94][5]  ( .D(n2091), .CK(clk), .Q(\ram[94][5] ) );
  DFFHQX1 \ram_reg[94][4]  ( .D(n2090), .CK(clk), .Q(\ram[94][4] ) );
  DFFHQX1 \ram_reg[94][3]  ( .D(n2089), .CK(clk), .Q(\ram[94][3] ) );
  DFFHQX1 \ram_reg[94][2]  ( .D(n2088), .CK(clk), .Q(\ram[94][2] ) );
  DFFHQX1 \ram_reg[94][1]  ( .D(n2087), .CK(clk), .Q(\ram[94][1] ) );
  DFFHQX1 \ram_reg[94][0]  ( .D(n2086), .CK(clk), .Q(\ram[94][0] ) );
  DFFHQX1 \ram_reg[90][15]  ( .D(n2037), .CK(clk), .Q(\ram[90][15] ) );
  DFFHQX1 \ram_reg[90][14]  ( .D(n2036), .CK(clk), .Q(\ram[90][14] ) );
  DFFHQX1 \ram_reg[90][13]  ( .D(n2035), .CK(clk), .Q(\ram[90][13] ) );
  DFFHQX1 \ram_reg[90][12]  ( .D(n2034), .CK(clk), .Q(\ram[90][12] ) );
  DFFHQX1 \ram_reg[90][11]  ( .D(n2033), .CK(clk), .Q(\ram[90][11] ) );
  DFFHQX1 \ram_reg[90][10]  ( .D(n2032), .CK(clk), .Q(\ram[90][10] ) );
  DFFHQX1 \ram_reg[90][9]  ( .D(n2031), .CK(clk), .Q(\ram[90][9] ) );
  DFFHQX1 \ram_reg[90][8]  ( .D(n2030), .CK(clk), .Q(\ram[90][8] ) );
  DFFHQX1 \ram_reg[90][7]  ( .D(n2029), .CK(clk), .Q(\ram[90][7] ) );
  DFFHQX1 \ram_reg[90][6]  ( .D(n2028), .CK(clk), .Q(\ram[90][6] ) );
  DFFHQX1 \ram_reg[90][5]  ( .D(n2027), .CK(clk), .Q(\ram[90][5] ) );
  DFFHQX1 \ram_reg[90][4]  ( .D(n2026), .CK(clk), .Q(\ram[90][4] ) );
  DFFHQX1 \ram_reg[90][3]  ( .D(n2025), .CK(clk), .Q(\ram[90][3] ) );
  DFFHQX1 \ram_reg[90][2]  ( .D(n2024), .CK(clk), .Q(\ram[90][2] ) );
  DFFHQX1 \ram_reg[90][1]  ( .D(n2023), .CK(clk), .Q(\ram[90][1] ) );
  DFFHQX1 \ram_reg[90][0]  ( .D(n2022), .CK(clk), .Q(\ram[90][0] ) );
  DFFHQX1 \ram_reg[86][15]  ( .D(n1973), .CK(clk), .Q(\ram[86][15] ) );
  DFFHQX1 \ram_reg[86][14]  ( .D(n1972), .CK(clk), .Q(\ram[86][14] ) );
  DFFHQX1 \ram_reg[86][13]  ( .D(n1971), .CK(clk), .Q(\ram[86][13] ) );
  DFFHQX1 \ram_reg[86][12]  ( .D(n1970), .CK(clk), .Q(\ram[86][12] ) );
  DFFHQX1 \ram_reg[86][11]  ( .D(n1969), .CK(clk), .Q(\ram[86][11] ) );
  DFFHQX1 \ram_reg[86][10]  ( .D(n1968), .CK(clk), .Q(\ram[86][10] ) );
  DFFHQX1 \ram_reg[86][9]  ( .D(n1967), .CK(clk), .Q(\ram[86][9] ) );
  DFFHQX1 \ram_reg[86][8]  ( .D(n1966), .CK(clk), .Q(\ram[86][8] ) );
  DFFHQX1 \ram_reg[86][7]  ( .D(n1965), .CK(clk), .Q(\ram[86][7] ) );
  DFFHQX1 \ram_reg[86][6]  ( .D(n1964), .CK(clk), .Q(\ram[86][6] ) );
  DFFHQX1 \ram_reg[86][5]  ( .D(n1963), .CK(clk), .Q(\ram[86][5] ) );
  DFFHQX1 \ram_reg[86][4]  ( .D(n1962), .CK(clk), .Q(\ram[86][4] ) );
  DFFHQX1 \ram_reg[86][3]  ( .D(n1961), .CK(clk), .Q(\ram[86][3] ) );
  DFFHQX1 \ram_reg[86][2]  ( .D(n1960), .CK(clk), .Q(\ram[86][2] ) );
  DFFHQX1 \ram_reg[86][1]  ( .D(n1959), .CK(clk), .Q(\ram[86][1] ) );
  DFFHQX1 \ram_reg[86][0]  ( .D(n1958), .CK(clk), .Q(\ram[86][0] ) );
  DFFHQX1 \ram_reg[82][15]  ( .D(n1909), .CK(clk), .Q(\ram[82][15] ) );
  DFFHQX1 \ram_reg[82][14]  ( .D(n1908), .CK(clk), .Q(\ram[82][14] ) );
  DFFHQX1 \ram_reg[82][13]  ( .D(n1907), .CK(clk), .Q(\ram[82][13] ) );
  DFFHQX1 \ram_reg[82][12]  ( .D(n1906), .CK(clk), .Q(\ram[82][12] ) );
  DFFHQX1 \ram_reg[82][11]  ( .D(n1905), .CK(clk), .Q(\ram[82][11] ) );
  DFFHQX1 \ram_reg[82][10]  ( .D(n1904), .CK(clk), .Q(\ram[82][10] ) );
  DFFHQX1 \ram_reg[82][9]  ( .D(n1903), .CK(clk), .Q(\ram[82][9] ) );
  DFFHQX1 \ram_reg[82][8]  ( .D(n1902), .CK(clk), .Q(\ram[82][8] ) );
  DFFHQX1 \ram_reg[82][7]  ( .D(n1901), .CK(clk), .Q(\ram[82][7] ) );
  DFFHQX1 \ram_reg[82][6]  ( .D(n1900), .CK(clk), .Q(\ram[82][6] ) );
  DFFHQX1 \ram_reg[82][5]  ( .D(n1899), .CK(clk), .Q(\ram[82][5] ) );
  DFFHQX1 \ram_reg[82][4]  ( .D(n1898), .CK(clk), .Q(\ram[82][4] ) );
  DFFHQX1 \ram_reg[82][3]  ( .D(n1897), .CK(clk), .Q(\ram[82][3] ) );
  DFFHQX1 \ram_reg[82][2]  ( .D(n1896), .CK(clk), .Q(\ram[82][2] ) );
  DFFHQX1 \ram_reg[82][1]  ( .D(n1895), .CK(clk), .Q(\ram[82][1] ) );
  DFFHQX1 \ram_reg[82][0]  ( .D(n1894), .CK(clk), .Q(\ram[82][0] ) );
  DFFHQX1 \ram_reg[78][15]  ( .D(n1845), .CK(clk), .Q(\ram[78][15] ) );
  DFFHQX1 \ram_reg[78][14]  ( .D(n1844), .CK(clk), .Q(\ram[78][14] ) );
  DFFHQX1 \ram_reg[78][13]  ( .D(n1843), .CK(clk), .Q(\ram[78][13] ) );
  DFFHQX1 \ram_reg[78][12]  ( .D(n1842), .CK(clk), .Q(\ram[78][12] ) );
  DFFHQX1 \ram_reg[78][11]  ( .D(n1841), .CK(clk), .Q(\ram[78][11] ) );
  DFFHQX1 \ram_reg[78][10]  ( .D(n1840), .CK(clk), .Q(\ram[78][10] ) );
  DFFHQX1 \ram_reg[78][9]  ( .D(n1839), .CK(clk), .Q(\ram[78][9] ) );
  DFFHQX1 \ram_reg[78][8]  ( .D(n1838), .CK(clk), .Q(\ram[78][8] ) );
  DFFHQX1 \ram_reg[78][7]  ( .D(n1837), .CK(clk), .Q(\ram[78][7] ) );
  DFFHQX1 \ram_reg[78][6]  ( .D(n1836), .CK(clk), .Q(\ram[78][6] ) );
  DFFHQX1 \ram_reg[78][5]  ( .D(n1835), .CK(clk), .Q(\ram[78][5] ) );
  DFFHQX1 \ram_reg[78][4]  ( .D(n1834), .CK(clk), .Q(\ram[78][4] ) );
  DFFHQX1 \ram_reg[78][3]  ( .D(n1833), .CK(clk), .Q(\ram[78][3] ) );
  DFFHQX1 \ram_reg[78][2]  ( .D(n1832), .CK(clk), .Q(\ram[78][2] ) );
  DFFHQX1 \ram_reg[78][1]  ( .D(n1831), .CK(clk), .Q(\ram[78][1] ) );
  DFFHQX1 \ram_reg[78][0]  ( .D(n1830), .CK(clk), .Q(\ram[78][0] ) );
  DFFHQX1 \ram_reg[74][15]  ( .D(n1781), .CK(clk), .Q(\ram[74][15] ) );
  DFFHQX1 \ram_reg[74][14]  ( .D(n1780), .CK(clk), .Q(\ram[74][14] ) );
  DFFHQX1 \ram_reg[74][13]  ( .D(n1779), .CK(clk), .Q(\ram[74][13] ) );
  DFFHQX1 \ram_reg[74][12]  ( .D(n1778), .CK(clk), .Q(\ram[74][12] ) );
  DFFHQX1 \ram_reg[74][11]  ( .D(n1777), .CK(clk), .Q(\ram[74][11] ) );
  DFFHQX1 \ram_reg[74][10]  ( .D(n1776), .CK(clk), .Q(\ram[74][10] ) );
  DFFHQX1 \ram_reg[74][9]  ( .D(n1775), .CK(clk), .Q(\ram[74][9] ) );
  DFFHQX1 \ram_reg[74][8]  ( .D(n1774), .CK(clk), .Q(\ram[74][8] ) );
  DFFHQX1 \ram_reg[74][7]  ( .D(n1773), .CK(clk), .Q(\ram[74][7] ) );
  DFFHQX1 \ram_reg[74][6]  ( .D(n1772), .CK(clk), .Q(\ram[74][6] ) );
  DFFHQX1 \ram_reg[74][5]  ( .D(n1771), .CK(clk), .Q(\ram[74][5] ) );
  DFFHQX1 \ram_reg[74][4]  ( .D(n1770), .CK(clk), .Q(\ram[74][4] ) );
  DFFHQX1 \ram_reg[74][3]  ( .D(n1769), .CK(clk), .Q(\ram[74][3] ) );
  DFFHQX1 \ram_reg[74][2]  ( .D(n1768), .CK(clk), .Q(\ram[74][2] ) );
  DFFHQX1 \ram_reg[74][1]  ( .D(n1767), .CK(clk), .Q(\ram[74][1] ) );
  DFFHQX1 \ram_reg[74][0]  ( .D(n1766), .CK(clk), .Q(\ram[74][0] ) );
  DFFHQX1 \ram_reg[70][15]  ( .D(n1717), .CK(clk), .Q(\ram[70][15] ) );
  DFFHQX1 \ram_reg[70][14]  ( .D(n1716), .CK(clk), .Q(\ram[70][14] ) );
  DFFHQX1 \ram_reg[70][13]  ( .D(n1715), .CK(clk), .Q(\ram[70][13] ) );
  DFFHQX1 \ram_reg[70][12]  ( .D(n1714), .CK(clk), .Q(\ram[70][12] ) );
  DFFHQX1 \ram_reg[70][11]  ( .D(n1713), .CK(clk), .Q(\ram[70][11] ) );
  DFFHQX1 \ram_reg[70][10]  ( .D(n1712), .CK(clk), .Q(\ram[70][10] ) );
  DFFHQX1 \ram_reg[70][9]  ( .D(n1711), .CK(clk), .Q(\ram[70][9] ) );
  DFFHQX1 \ram_reg[70][8]  ( .D(n1710), .CK(clk), .Q(\ram[70][8] ) );
  DFFHQX1 \ram_reg[70][7]  ( .D(n1709), .CK(clk), .Q(\ram[70][7] ) );
  DFFHQX1 \ram_reg[70][6]  ( .D(n1708), .CK(clk), .Q(\ram[70][6] ) );
  DFFHQX1 \ram_reg[70][5]  ( .D(n1707), .CK(clk), .Q(\ram[70][5] ) );
  DFFHQX1 \ram_reg[70][4]  ( .D(n1706), .CK(clk), .Q(\ram[70][4] ) );
  DFFHQX1 \ram_reg[70][3]  ( .D(n1705), .CK(clk), .Q(\ram[70][3] ) );
  DFFHQX1 \ram_reg[70][2]  ( .D(n1704), .CK(clk), .Q(\ram[70][2] ) );
  DFFHQX1 \ram_reg[70][1]  ( .D(n1703), .CK(clk), .Q(\ram[70][1] ) );
  DFFHQX1 \ram_reg[70][0]  ( .D(n1702), .CK(clk), .Q(\ram[70][0] ) );
  DFFHQX1 \ram_reg[66][15]  ( .D(n1653), .CK(clk), .Q(\ram[66][15] ) );
  DFFHQX1 \ram_reg[66][14]  ( .D(n1652), .CK(clk), .Q(\ram[66][14] ) );
  DFFHQX1 \ram_reg[66][13]  ( .D(n1651), .CK(clk), .Q(\ram[66][13] ) );
  DFFHQX1 \ram_reg[66][12]  ( .D(n1650), .CK(clk), .Q(\ram[66][12] ) );
  DFFHQX1 \ram_reg[66][11]  ( .D(n1649), .CK(clk), .Q(\ram[66][11] ) );
  DFFHQX1 \ram_reg[66][10]  ( .D(n1648), .CK(clk), .Q(\ram[66][10] ) );
  DFFHQX1 \ram_reg[66][9]  ( .D(n1647), .CK(clk), .Q(\ram[66][9] ) );
  DFFHQX1 \ram_reg[66][8]  ( .D(n1646), .CK(clk), .Q(\ram[66][8] ) );
  DFFHQX1 \ram_reg[66][7]  ( .D(n1645), .CK(clk), .Q(\ram[66][7] ) );
  DFFHQX1 \ram_reg[66][6]  ( .D(n1644), .CK(clk), .Q(\ram[66][6] ) );
  DFFHQX1 \ram_reg[66][5]  ( .D(n1643), .CK(clk), .Q(\ram[66][5] ) );
  DFFHQX1 \ram_reg[66][4]  ( .D(n1642), .CK(clk), .Q(\ram[66][4] ) );
  DFFHQX1 \ram_reg[66][3]  ( .D(n1641), .CK(clk), .Q(\ram[66][3] ) );
  DFFHQX1 \ram_reg[66][2]  ( .D(n1640), .CK(clk), .Q(\ram[66][2] ) );
  DFFHQX1 \ram_reg[66][1]  ( .D(n1639), .CK(clk), .Q(\ram[66][1] ) );
  DFFHQX1 \ram_reg[66][0]  ( .D(n1638), .CK(clk), .Q(\ram[66][0] ) );
  DFFHQX1 \ram_reg[62][15]  ( .D(n1589), .CK(clk), .Q(\ram[62][15] ) );
  DFFHQX1 \ram_reg[62][14]  ( .D(n1588), .CK(clk), .Q(\ram[62][14] ) );
  DFFHQX1 \ram_reg[62][13]  ( .D(n1587), .CK(clk), .Q(\ram[62][13] ) );
  DFFHQX1 \ram_reg[62][12]  ( .D(n1586), .CK(clk), .Q(\ram[62][12] ) );
  DFFHQX1 \ram_reg[62][11]  ( .D(n1585), .CK(clk), .Q(\ram[62][11] ) );
  DFFHQX1 \ram_reg[62][10]  ( .D(n1584), .CK(clk), .Q(\ram[62][10] ) );
  DFFHQX1 \ram_reg[62][9]  ( .D(n1583), .CK(clk), .Q(\ram[62][9] ) );
  DFFHQX1 \ram_reg[62][8]  ( .D(n1582), .CK(clk), .Q(\ram[62][8] ) );
  DFFHQX1 \ram_reg[62][7]  ( .D(n1581), .CK(clk), .Q(\ram[62][7] ) );
  DFFHQX1 \ram_reg[62][6]  ( .D(n1580), .CK(clk), .Q(\ram[62][6] ) );
  DFFHQX1 \ram_reg[62][5]  ( .D(n1579), .CK(clk), .Q(\ram[62][5] ) );
  DFFHQX1 \ram_reg[62][4]  ( .D(n1578), .CK(clk), .Q(\ram[62][4] ) );
  DFFHQX1 \ram_reg[62][3]  ( .D(n1577), .CK(clk), .Q(\ram[62][3] ) );
  DFFHQX1 \ram_reg[62][2]  ( .D(n1576), .CK(clk), .Q(\ram[62][2] ) );
  DFFHQX1 \ram_reg[62][1]  ( .D(n1575), .CK(clk), .Q(\ram[62][1] ) );
  DFFHQX1 \ram_reg[62][0]  ( .D(n1574), .CK(clk), .Q(\ram[62][0] ) );
  DFFHQX1 \ram_reg[58][15]  ( .D(n1525), .CK(clk), .Q(\ram[58][15] ) );
  DFFHQX1 \ram_reg[58][14]  ( .D(n1524), .CK(clk), .Q(\ram[58][14] ) );
  DFFHQX1 \ram_reg[58][13]  ( .D(n1523), .CK(clk), .Q(\ram[58][13] ) );
  DFFHQX1 \ram_reg[58][12]  ( .D(n1522), .CK(clk), .Q(\ram[58][12] ) );
  DFFHQX1 \ram_reg[58][11]  ( .D(n1521), .CK(clk), .Q(\ram[58][11] ) );
  DFFHQX1 \ram_reg[58][10]  ( .D(n1520), .CK(clk), .Q(\ram[58][10] ) );
  DFFHQX1 \ram_reg[58][9]  ( .D(n1519), .CK(clk), .Q(\ram[58][9] ) );
  DFFHQX1 \ram_reg[58][8]  ( .D(n1518), .CK(clk), .Q(\ram[58][8] ) );
  DFFHQX1 \ram_reg[58][7]  ( .D(n1517), .CK(clk), .Q(\ram[58][7] ) );
  DFFHQX1 \ram_reg[58][6]  ( .D(n1516), .CK(clk), .Q(\ram[58][6] ) );
  DFFHQX1 \ram_reg[58][5]  ( .D(n1515), .CK(clk), .Q(\ram[58][5] ) );
  DFFHQX1 \ram_reg[58][4]  ( .D(n1514), .CK(clk), .Q(\ram[58][4] ) );
  DFFHQX1 \ram_reg[58][3]  ( .D(n1513), .CK(clk), .Q(\ram[58][3] ) );
  DFFHQX1 \ram_reg[58][2]  ( .D(n1512), .CK(clk), .Q(\ram[58][2] ) );
  DFFHQX1 \ram_reg[58][1]  ( .D(n1511), .CK(clk), .Q(\ram[58][1] ) );
  DFFHQX1 \ram_reg[58][0]  ( .D(n1510), .CK(clk), .Q(\ram[58][0] ) );
  DFFHQX1 \ram_reg[54][15]  ( .D(n1461), .CK(clk), .Q(\ram[54][15] ) );
  DFFHQX1 \ram_reg[54][14]  ( .D(n1460), .CK(clk), .Q(\ram[54][14] ) );
  DFFHQX1 \ram_reg[54][13]  ( .D(n1459), .CK(clk), .Q(\ram[54][13] ) );
  DFFHQX1 \ram_reg[54][12]  ( .D(n1458), .CK(clk), .Q(\ram[54][12] ) );
  DFFHQX1 \ram_reg[54][11]  ( .D(n1457), .CK(clk), .Q(\ram[54][11] ) );
  DFFHQX1 \ram_reg[54][10]  ( .D(n1456), .CK(clk), .Q(\ram[54][10] ) );
  DFFHQX1 \ram_reg[54][9]  ( .D(n1455), .CK(clk), .Q(\ram[54][9] ) );
  DFFHQX1 \ram_reg[54][8]  ( .D(n1454), .CK(clk), .Q(\ram[54][8] ) );
  DFFHQX1 \ram_reg[54][7]  ( .D(n1453), .CK(clk), .Q(\ram[54][7] ) );
  DFFHQX1 \ram_reg[54][6]  ( .D(n1452), .CK(clk), .Q(\ram[54][6] ) );
  DFFHQX1 \ram_reg[54][5]  ( .D(n1451), .CK(clk), .Q(\ram[54][5] ) );
  DFFHQX1 \ram_reg[54][4]  ( .D(n1450), .CK(clk), .Q(\ram[54][4] ) );
  DFFHQX1 \ram_reg[54][3]  ( .D(n1449), .CK(clk), .Q(\ram[54][3] ) );
  DFFHQX1 \ram_reg[54][2]  ( .D(n1448), .CK(clk), .Q(\ram[54][2] ) );
  DFFHQX1 \ram_reg[54][1]  ( .D(n1447), .CK(clk), .Q(\ram[54][1] ) );
  DFFHQX1 \ram_reg[54][0]  ( .D(n1446), .CK(clk), .Q(\ram[54][0] ) );
  DFFHQX1 \ram_reg[50][15]  ( .D(n1397), .CK(clk), .Q(\ram[50][15] ) );
  DFFHQX1 \ram_reg[50][14]  ( .D(n1396), .CK(clk), .Q(\ram[50][14] ) );
  DFFHQX1 \ram_reg[50][13]  ( .D(n1395), .CK(clk), .Q(\ram[50][13] ) );
  DFFHQX1 \ram_reg[50][12]  ( .D(n1394), .CK(clk), .Q(\ram[50][12] ) );
  DFFHQX1 \ram_reg[50][11]  ( .D(n1393), .CK(clk), .Q(\ram[50][11] ) );
  DFFHQX1 \ram_reg[50][10]  ( .D(n1392), .CK(clk), .Q(\ram[50][10] ) );
  DFFHQX1 \ram_reg[50][9]  ( .D(n1391), .CK(clk), .Q(\ram[50][9] ) );
  DFFHQX1 \ram_reg[50][8]  ( .D(n1390), .CK(clk), .Q(\ram[50][8] ) );
  DFFHQX1 \ram_reg[50][7]  ( .D(n1389), .CK(clk), .Q(\ram[50][7] ) );
  DFFHQX1 \ram_reg[50][6]  ( .D(n1388), .CK(clk), .Q(\ram[50][6] ) );
  DFFHQX1 \ram_reg[50][5]  ( .D(n1387), .CK(clk), .Q(\ram[50][5] ) );
  DFFHQX1 \ram_reg[50][4]  ( .D(n1386), .CK(clk), .Q(\ram[50][4] ) );
  DFFHQX1 \ram_reg[50][3]  ( .D(n1385), .CK(clk), .Q(\ram[50][3] ) );
  DFFHQX1 \ram_reg[50][2]  ( .D(n1384), .CK(clk), .Q(\ram[50][2] ) );
  DFFHQX1 \ram_reg[50][1]  ( .D(n1383), .CK(clk), .Q(\ram[50][1] ) );
  DFFHQX1 \ram_reg[50][0]  ( .D(n1382), .CK(clk), .Q(\ram[50][0] ) );
  DFFHQX1 \ram_reg[46][15]  ( .D(n1333), .CK(clk), .Q(\ram[46][15] ) );
  DFFHQX1 \ram_reg[46][14]  ( .D(n1332), .CK(clk), .Q(\ram[46][14] ) );
  DFFHQX1 \ram_reg[46][13]  ( .D(n1331), .CK(clk), .Q(\ram[46][13] ) );
  DFFHQX1 \ram_reg[46][12]  ( .D(n1330), .CK(clk), .Q(\ram[46][12] ) );
  DFFHQX1 \ram_reg[46][11]  ( .D(n1329), .CK(clk), .Q(\ram[46][11] ) );
  DFFHQX1 \ram_reg[46][10]  ( .D(n1328), .CK(clk), .Q(\ram[46][10] ) );
  DFFHQX1 \ram_reg[46][9]  ( .D(n1327), .CK(clk), .Q(\ram[46][9] ) );
  DFFHQX1 \ram_reg[46][8]  ( .D(n1326), .CK(clk), .Q(\ram[46][8] ) );
  DFFHQX1 \ram_reg[46][7]  ( .D(n1325), .CK(clk), .Q(\ram[46][7] ) );
  DFFHQX1 \ram_reg[46][6]  ( .D(n1324), .CK(clk), .Q(\ram[46][6] ) );
  DFFHQX1 \ram_reg[46][5]  ( .D(n1323), .CK(clk), .Q(\ram[46][5] ) );
  DFFHQX1 \ram_reg[46][4]  ( .D(n1322), .CK(clk), .Q(\ram[46][4] ) );
  DFFHQX1 \ram_reg[46][3]  ( .D(n1321), .CK(clk), .Q(\ram[46][3] ) );
  DFFHQX1 \ram_reg[46][2]  ( .D(n1320), .CK(clk), .Q(\ram[46][2] ) );
  DFFHQX1 \ram_reg[46][1]  ( .D(n1319), .CK(clk), .Q(\ram[46][1] ) );
  DFFHQX1 \ram_reg[46][0]  ( .D(n1318), .CK(clk), .Q(\ram[46][0] ) );
  DFFHQX1 \ram_reg[42][15]  ( .D(n1269), .CK(clk), .Q(\ram[42][15] ) );
  DFFHQX1 \ram_reg[42][14]  ( .D(n1268), .CK(clk), .Q(\ram[42][14] ) );
  DFFHQX1 \ram_reg[42][13]  ( .D(n1267), .CK(clk), .Q(\ram[42][13] ) );
  DFFHQX1 \ram_reg[42][12]  ( .D(n1266), .CK(clk), .Q(\ram[42][12] ) );
  DFFHQX1 \ram_reg[42][11]  ( .D(n1265), .CK(clk), .Q(\ram[42][11] ) );
  DFFHQX1 \ram_reg[42][10]  ( .D(n1264), .CK(clk), .Q(\ram[42][10] ) );
  DFFHQX1 \ram_reg[42][9]  ( .D(n1263), .CK(clk), .Q(\ram[42][9] ) );
  DFFHQX1 \ram_reg[42][8]  ( .D(n1262), .CK(clk), .Q(\ram[42][8] ) );
  DFFHQX1 \ram_reg[42][7]  ( .D(n1261), .CK(clk), .Q(\ram[42][7] ) );
  DFFHQX1 \ram_reg[42][6]  ( .D(n1260), .CK(clk), .Q(\ram[42][6] ) );
  DFFHQX1 \ram_reg[42][5]  ( .D(n1259), .CK(clk), .Q(\ram[42][5] ) );
  DFFHQX1 \ram_reg[42][4]  ( .D(n1258), .CK(clk), .Q(\ram[42][4] ) );
  DFFHQX1 \ram_reg[42][3]  ( .D(n1257), .CK(clk), .Q(\ram[42][3] ) );
  DFFHQX1 \ram_reg[42][2]  ( .D(n1256), .CK(clk), .Q(\ram[42][2] ) );
  DFFHQX1 \ram_reg[42][1]  ( .D(n1255), .CK(clk), .Q(\ram[42][1] ) );
  DFFHQX1 \ram_reg[42][0]  ( .D(n1254), .CK(clk), .Q(\ram[42][0] ) );
  DFFHQX1 \ram_reg[38][15]  ( .D(n1205), .CK(clk), .Q(\ram[38][15] ) );
  DFFHQX1 \ram_reg[38][14]  ( .D(n1204), .CK(clk), .Q(\ram[38][14] ) );
  DFFHQX1 \ram_reg[38][13]  ( .D(n1203), .CK(clk), .Q(\ram[38][13] ) );
  DFFHQX1 \ram_reg[38][12]  ( .D(n1202), .CK(clk), .Q(\ram[38][12] ) );
  DFFHQX1 \ram_reg[38][11]  ( .D(n1201), .CK(clk), .Q(\ram[38][11] ) );
  DFFHQX1 \ram_reg[38][10]  ( .D(n1200), .CK(clk), .Q(\ram[38][10] ) );
  DFFHQX1 \ram_reg[38][9]  ( .D(n1199), .CK(clk), .Q(\ram[38][9] ) );
  DFFHQX1 \ram_reg[38][8]  ( .D(n1198), .CK(clk), .Q(\ram[38][8] ) );
  DFFHQX1 \ram_reg[38][7]  ( .D(n1197), .CK(clk), .Q(\ram[38][7] ) );
  DFFHQX1 \ram_reg[38][6]  ( .D(n1196), .CK(clk), .Q(\ram[38][6] ) );
  DFFHQX1 \ram_reg[38][5]  ( .D(n1195), .CK(clk), .Q(\ram[38][5] ) );
  DFFHQX1 \ram_reg[38][4]  ( .D(n1194), .CK(clk), .Q(\ram[38][4] ) );
  DFFHQX1 \ram_reg[38][3]  ( .D(n1193), .CK(clk), .Q(\ram[38][3] ) );
  DFFHQX1 \ram_reg[38][2]  ( .D(n1192), .CK(clk), .Q(\ram[38][2] ) );
  DFFHQX1 \ram_reg[38][1]  ( .D(n1191), .CK(clk), .Q(\ram[38][1] ) );
  DFFHQX1 \ram_reg[38][0]  ( .D(n1190), .CK(clk), .Q(\ram[38][0] ) );
  DFFHQX1 \ram_reg[34][15]  ( .D(n1141), .CK(clk), .Q(\ram[34][15] ) );
  DFFHQX1 \ram_reg[34][14]  ( .D(n1140), .CK(clk), .Q(\ram[34][14] ) );
  DFFHQX1 \ram_reg[34][13]  ( .D(n1139), .CK(clk), .Q(\ram[34][13] ) );
  DFFHQX1 \ram_reg[34][12]  ( .D(n1138), .CK(clk), .Q(\ram[34][12] ) );
  DFFHQX1 \ram_reg[34][11]  ( .D(n1137), .CK(clk), .Q(\ram[34][11] ) );
  DFFHQX1 \ram_reg[34][10]  ( .D(n1136), .CK(clk), .Q(\ram[34][10] ) );
  DFFHQX1 \ram_reg[34][9]  ( .D(n1135), .CK(clk), .Q(\ram[34][9] ) );
  DFFHQX1 \ram_reg[34][8]  ( .D(n1134), .CK(clk), .Q(\ram[34][8] ) );
  DFFHQX1 \ram_reg[34][7]  ( .D(n1133), .CK(clk), .Q(\ram[34][7] ) );
  DFFHQX1 \ram_reg[34][6]  ( .D(n1132), .CK(clk), .Q(\ram[34][6] ) );
  DFFHQX1 \ram_reg[34][5]  ( .D(n1131), .CK(clk), .Q(\ram[34][5] ) );
  DFFHQX1 \ram_reg[34][4]  ( .D(n1130), .CK(clk), .Q(\ram[34][4] ) );
  DFFHQX1 \ram_reg[34][3]  ( .D(n1129), .CK(clk), .Q(\ram[34][3] ) );
  DFFHQX1 \ram_reg[34][2]  ( .D(n1128), .CK(clk), .Q(\ram[34][2] ) );
  DFFHQX1 \ram_reg[34][1]  ( .D(n1127), .CK(clk), .Q(\ram[34][1] ) );
  DFFHQX1 \ram_reg[34][0]  ( .D(n1126), .CK(clk), .Q(\ram[34][0] ) );
  DFFHQX1 \ram_reg[30][15]  ( .D(n1077), .CK(clk), .Q(\ram[30][15] ) );
  DFFHQX1 \ram_reg[30][14]  ( .D(n1076), .CK(clk), .Q(\ram[30][14] ) );
  DFFHQX1 \ram_reg[30][13]  ( .D(n1075), .CK(clk), .Q(\ram[30][13] ) );
  DFFHQX1 \ram_reg[30][12]  ( .D(n1074), .CK(clk), .Q(\ram[30][12] ) );
  DFFHQX1 \ram_reg[30][11]  ( .D(n1073), .CK(clk), .Q(\ram[30][11] ) );
  DFFHQX1 \ram_reg[30][10]  ( .D(n1072), .CK(clk), .Q(\ram[30][10] ) );
  DFFHQX1 \ram_reg[30][9]  ( .D(n1071), .CK(clk), .Q(\ram[30][9] ) );
  DFFHQX1 \ram_reg[30][8]  ( .D(n1070), .CK(clk), .Q(\ram[30][8] ) );
  DFFHQX1 \ram_reg[30][7]  ( .D(n1069), .CK(clk), .Q(\ram[30][7] ) );
  DFFHQX1 \ram_reg[30][6]  ( .D(n1068), .CK(clk), .Q(\ram[30][6] ) );
  DFFHQX1 \ram_reg[30][5]  ( .D(n1067), .CK(clk), .Q(\ram[30][5] ) );
  DFFHQX1 \ram_reg[30][4]  ( .D(n1066), .CK(clk), .Q(\ram[30][4] ) );
  DFFHQX1 \ram_reg[30][3]  ( .D(n1065), .CK(clk), .Q(\ram[30][3] ) );
  DFFHQX1 \ram_reg[30][2]  ( .D(n1064), .CK(clk), .Q(\ram[30][2] ) );
  DFFHQX1 \ram_reg[30][1]  ( .D(n1063), .CK(clk), .Q(\ram[30][1] ) );
  DFFHQX1 \ram_reg[30][0]  ( .D(n1062), .CK(clk), .Q(\ram[30][0] ) );
  DFFHQX1 \ram_reg[26][15]  ( .D(n1013), .CK(clk), .Q(\ram[26][15] ) );
  DFFHQX1 \ram_reg[26][14]  ( .D(n1012), .CK(clk), .Q(\ram[26][14] ) );
  DFFHQX1 \ram_reg[26][13]  ( .D(n1011), .CK(clk), .Q(\ram[26][13] ) );
  DFFHQX1 \ram_reg[26][12]  ( .D(n1010), .CK(clk), .Q(\ram[26][12] ) );
  DFFHQX1 \ram_reg[26][11]  ( .D(n1009), .CK(clk), .Q(\ram[26][11] ) );
  DFFHQX1 \ram_reg[26][10]  ( .D(n1008), .CK(clk), .Q(\ram[26][10] ) );
  DFFHQX1 \ram_reg[26][9]  ( .D(n1007), .CK(clk), .Q(\ram[26][9] ) );
  DFFHQX1 \ram_reg[26][8]  ( .D(n1006), .CK(clk), .Q(\ram[26][8] ) );
  DFFHQX1 \ram_reg[26][7]  ( .D(n1005), .CK(clk), .Q(\ram[26][7] ) );
  DFFHQX1 \ram_reg[26][6]  ( .D(n1004), .CK(clk), .Q(\ram[26][6] ) );
  DFFHQX1 \ram_reg[26][5]  ( .D(n1003), .CK(clk), .Q(\ram[26][5] ) );
  DFFHQX1 \ram_reg[26][4]  ( .D(n1002), .CK(clk), .Q(\ram[26][4] ) );
  DFFHQX1 \ram_reg[26][3]  ( .D(n1001), .CK(clk), .Q(\ram[26][3] ) );
  DFFHQX1 \ram_reg[26][2]  ( .D(n1000), .CK(clk), .Q(\ram[26][2] ) );
  DFFHQX1 \ram_reg[26][1]  ( .D(n999), .CK(clk), .Q(\ram[26][1] ) );
  DFFHQX1 \ram_reg[26][0]  ( .D(n998), .CK(clk), .Q(\ram[26][0] ) );
  DFFHQX1 \ram_reg[22][15]  ( .D(n949), .CK(clk), .Q(\ram[22][15] ) );
  DFFHQX1 \ram_reg[22][14]  ( .D(n948), .CK(clk), .Q(\ram[22][14] ) );
  DFFHQX1 \ram_reg[22][13]  ( .D(n947), .CK(clk), .Q(\ram[22][13] ) );
  DFFHQX1 \ram_reg[22][12]  ( .D(n946), .CK(clk), .Q(\ram[22][12] ) );
  DFFHQX1 \ram_reg[22][11]  ( .D(n945), .CK(clk), .Q(\ram[22][11] ) );
  DFFHQX1 \ram_reg[22][10]  ( .D(n944), .CK(clk), .Q(\ram[22][10] ) );
  DFFHQX1 \ram_reg[22][9]  ( .D(n943), .CK(clk), .Q(\ram[22][9] ) );
  DFFHQX1 \ram_reg[22][8]  ( .D(n942), .CK(clk), .Q(\ram[22][8] ) );
  DFFHQX1 \ram_reg[22][7]  ( .D(n941), .CK(clk), .Q(\ram[22][7] ) );
  DFFHQX1 \ram_reg[22][6]  ( .D(n940), .CK(clk), .Q(\ram[22][6] ) );
  DFFHQX1 \ram_reg[22][5]  ( .D(n939), .CK(clk), .Q(\ram[22][5] ) );
  DFFHQX1 \ram_reg[22][4]  ( .D(n938), .CK(clk), .Q(\ram[22][4] ) );
  DFFHQX1 \ram_reg[22][3]  ( .D(n937), .CK(clk), .Q(\ram[22][3] ) );
  DFFHQX1 \ram_reg[22][2]  ( .D(n936), .CK(clk), .Q(\ram[22][2] ) );
  DFFHQX1 \ram_reg[22][1]  ( .D(n935), .CK(clk), .Q(\ram[22][1] ) );
  DFFHQX1 \ram_reg[22][0]  ( .D(n934), .CK(clk), .Q(\ram[22][0] ) );
  DFFHQX1 \ram_reg[18][15]  ( .D(n885), .CK(clk), .Q(\ram[18][15] ) );
  DFFHQX1 \ram_reg[18][14]  ( .D(n884), .CK(clk), .Q(\ram[18][14] ) );
  DFFHQX1 \ram_reg[18][13]  ( .D(n883), .CK(clk), .Q(\ram[18][13] ) );
  DFFHQX1 \ram_reg[18][12]  ( .D(n882), .CK(clk), .Q(\ram[18][12] ) );
  DFFHQX1 \ram_reg[18][11]  ( .D(n881), .CK(clk), .Q(\ram[18][11] ) );
  DFFHQX1 \ram_reg[18][10]  ( .D(n880), .CK(clk), .Q(\ram[18][10] ) );
  DFFHQX1 \ram_reg[18][9]  ( .D(n879), .CK(clk), .Q(\ram[18][9] ) );
  DFFHQX1 \ram_reg[18][8]  ( .D(n878), .CK(clk), .Q(\ram[18][8] ) );
  DFFHQX1 \ram_reg[18][7]  ( .D(n877), .CK(clk), .Q(\ram[18][7] ) );
  DFFHQX1 \ram_reg[18][6]  ( .D(n876), .CK(clk), .Q(\ram[18][6] ) );
  DFFHQX1 \ram_reg[18][5]  ( .D(n875), .CK(clk), .Q(\ram[18][5] ) );
  DFFHQX1 \ram_reg[18][4]  ( .D(n874), .CK(clk), .Q(\ram[18][4] ) );
  DFFHQX1 \ram_reg[18][3]  ( .D(n873), .CK(clk), .Q(\ram[18][3] ) );
  DFFHQX1 \ram_reg[18][2]  ( .D(n872), .CK(clk), .Q(\ram[18][2] ) );
  DFFHQX1 \ram_reg[18][1]  ( .D(n871), .CK(clk), .Q(\ram[18][1] ) );
  DFFHQX1 \ram_reg[18][0]  ( .D(n870), .CK(clk), .Q(\ram[18][0] ) );
  DFFHQX1 \ram_reg[14][15]  ( .D(n821), .CK(clk), .Q(\ram[14][15] ) );
  DFFHQX1 \ram_reg[14][14]  ( .D(n820), .CK(clk), .Q(\ram[14][14] ) );
  DFFHQX1 \ram_reg[14][13]  ( .D(n819), .CK(clk), .Q(\ram[14][13] ) );
  DFFHQX1 \ram_reg[14][12]  ( .D(n818), .CK(clk), .Q(\ram[14][12] ) );
  DFFHQX1 \ram_reg[14][11]  ( .D(n817), .CK(clk), .Q(\ram[14][11] ) );
  DFFHQX1 \ram_reg[14][10]  ( .D(n816), .CK(clk), .Q(\ram[14][10] ) );
  DFFHQX1 \ram_reg[14][9]  ( .D(n815), .CK(clk), .Q(\ram[14][9] ) );
  DFFHQX1 \ram_reg[14][8]  ( .D(n814), .CK(clk), .Q(\ram[14][8] ) );
  DFFHQX1 \ram_reg[14][7]  ( .D(n813), .CK(clk), .Q(\ram[14][7] ) );
  DFFHQX1 \ram_reg[14][6]  ( .D(n812), .CK(clk), .Q(\ram[14][6] ) );
  DFFHQX1 \ram_reg[14][5]  ( .D(n811), .CK(clk), .Q(\ram[14][5] ) );
  DFFHQX1 \ram_reg[14][4]  ( .D(n810), .CK(clk), .Q(\ram[14][4] ) );
  DFFHQX1 \ram_reg[14][3]  ( .D(n809), .CK(clk), .Q(\ram[14][3] ) );
  DFFHQX1 \ram_reg[14][2]  ( .D(n808), .CK(clk), .Q(\ram[14][2] ) );
  DFFHQX1 \ram_reg[14][1]  ( .D(n807), .CK(clk), .Q(\ram[14][1] ) );
  DFFHQX1 \ram_reg[14][0]  ( .D(n806), .CK(clk), .Q(\ram[14][0] ) );
  DFFHQX1 \ram_reg[10][15]  ( .D(n757), .CK(clk), .Q(\ram[10][15] ) );
  DFFHQX1 \ram_reg[10][14]  ( .D(n756), .CK(clk), .Q(\ram[10][14] ) );
  DFFHQX1 \ram_reg[10][13]  ( .D(n755), .CK(clk), .Q(\ram[10][13] ) );
  DFFHQX1 \ram_reg[10][12]  ( .D(n754), .CK(clk), .Q(\ram[10][12] ) );
  DFFHQX1 \ram_reg[10][11]  ( .D(n753), .CK(clk), .Q(\ram[10][11] ) );
  DFFHQX1 \ram_reg[10][10]  ( .D(n752), .CK(clk), .Q(\ram[10][10] ) );
  DFFHQX1 \ram_reg[10][9]  ( .D(n751), .CK(clk), .Q(\ram[10][9] ) );
  DFFHQX1 \ram_reg[10][8]  ( .D(n750), .CK(clk), .Q(\ram[10][8] ) );
  DFFHQX1 \ram_reg[10][7]  ( .D(n749), .CK(clk), .Q(\ram[10][7] ) );
  DFFHQX1 \ram_reg[10][6]  ( .D(n748), .CK(clk), .Q(\ram[10][6] ) );
  DFFHQX1 \ram_reg[10][5]  ( .D(n747), .CK(clk), .Q(\ram[10][5] ) );
  DFFHQX1 \ram_reg[10][4]  ( .D(n746), .CK(clk), .Q(\ram[10][4] ) );
  DFFHQX1 \ram_reg[10][3]  ( .D(n745), .CK(clk), .Q(\ram[10][3] ) );
  DFFHQX1 \ram_reg[10][2]  ( .D(n744), .CK(clk), .Q(\ram[10][2] ) );
  DFFHQX1 \ram_reg[10][1]  ( .D(n743), .CK(clk), .Q(\ram[10][1] ) );
  DFFHQX1 \ram_reg[10][0]  ( .D(n742), .CK(clk), .Q(\ram[10][0] ) );
  DFFHQX1 \ram_reg[6][15]  ( .D(n693), .CK(clk), .Q(\ram[6][15] ) );
  DFFHQX1 \ram_reg[6][14]  ( .D(n692), .CK(clk), .Q(\ram[6][14] ) );
  DFFHQX1 \ram_reg[6][13]  ( .D(n691), .CK(clk), .Q(\ram[6][13] ) );
  DFFHQX1 \ram_reg[6][12]  ( .D(n690), .CK(clk), .Q(\ram[6][12] ) );
  DFFHQX1 \ram_reg[6][11]  ( .D(n689), .CK(clk), .Q(\ram[6][11] ) );
  DFFHQX1 \ram_reg[6][10]  ( .D(n688), .CK(clk), .Q(\ram[6][10] ) );
  DFFHQX1 \ram_reg[6][9]  ( .D(n687), .CK(clk), .Q(\ram[6][9] ) );
  DFFHQX1 \ram_reg[6][8]  ( .D(n686), .CK(clk), .Q(\ram[6][8] ) );
  DFFHQX1 \ram_reg[6][7]  ( .D(n685), .CK(clk), .Q(\ram[6][7] ) );
  DFFHQX1 \ram_reg[6][6]  ( .D(n684), .CK(clk), .Q(\ram[6][6] ) );
  DFFHQX1 \ram_reg[6][5]  ( .D(n683), .CK(clk), .Q(\ram[6][5] ) );
  DFFHQX1 \ram_reg[6][4]  ( .D(n682), .CK(clk), .Q(\ram[6][4] ) );
  DFFHQX1 \ram_reg[6][3]  ( .D(n681), .CK(clk), .Q(\ram[6][3] ) );
  DFFHQX1 \ram_reg[6][2]  ( .D(n680), .CK(clk), .Q(\ram[6][2] ) );
  DFFHQX1 \ram_reg[6][1]  ( .D(n679), .CK(clk), .Q(\ram[6][1] ) );
  DFFHQX1 \ram_reg[6][0]  ( .D(n678), .CK(clk), .Q(\ram[6][0] ) );
  DFFHQX1 \ram_reg[2][15]  ( .D(n629), .CK(clk), .Q(\ram[2][15] ) );
  DFFHQX1 \ram_reg[2][14]  ( .D(n628), .CK(clk), .Q(\ram[2][14] ) );
  DFFHQX1 \ram_reg[2][13]  ( .D(n627), .CK(clk), .Q(\ram[2][13] ) );
  DFFHQX1 \ram_reg[2][12]  ( .D(n626), .CK(clk), .Q(\ram[2][12] ) );
  DFFHQX1 \ram_reg[2][11]  ( .D(n625), .CK(clk), .Q(\ram[2][11] ) );
  DFFHQX1 \ram_reg[2][10]  ( .D(n624), .CK(clk), .Q(\ram[2][10] ) );
  DFFHQX1 \ram_reg[2][9]  ( .D(n623), .CK(clk), .Q(\ram[2][9] ) );
  DFFHQX1 \ram_reg[2][8]  ( .D(n622), .CK(clk), .Q(\ram[2][8] ) );
  DFFHQX1 \ram_reg[2][7]  ( .D(n621), .CK(clk), .Q(\ram[2][7] ) );
  DFFHQX1 \ram_reg[2][6]  ( .D(n620), .CK(clk), .Q(\ram[2][6] ) );
  DFFHQX1 \ram_reg[2][5]  ( .D(n619), .CK(clk), .Q(\ram[2][5] ) );
  DFFHQX1 \ram_reg[2][4]  ( .D(n618), .CK(clk), .Q(\ram[2][4] ) );
  DFFHQX1 \ram_reg[2][3]  ( .D(n617), .CK(clk), .Q(\ram[2][3] ) );
  DFFHQX1 \ram_reg[2][2]  ( .D(n616), .CK(clk), .Q(\ram[2][2] ) );
  DFFHQX1 \ram_reg[2][1]  ( .D(n615), .CK(clk), .Q(\ram[2][1] ) );
  DFFHQX1 \ram_reg[2][0]  ( .D(n614), .CK(clk), .Q(\ram[2][0] ) );
  AND2X2 U2 ( .A(mem_write_data[4]), .B(n6992), .Y(n1) );
  AND2X2 U3 ( .A(mem_write_data[5]), .B(n6992), .Y(n2) );
  AND2X2 U4 ( .A(mem_write_data[6]), .B(n6992), .Y(n3) );
  AND2X2 U5 ( .A(mem_write_data[7]), .B(n6992), .Y(n4) );
  AND2X2 U6 ( .A(mem_write_data[8]), .B(n6992), .Y(n5) );
  AND2X2 U7 ( .A(mem_write_data[9]), .B(n6992), .Y(n6) );
  AND2X2 U8 ( .A(mem_write_data[10]), .B(n6992), .Y(n12) );
  AND2X2 U9 ( .A(mem_write_data[11]), .B(n6992), .Y(n13) );
  AND2X2 U10 ( .A(mem_write_data[12]), .B(n6992), .Y(n14) );
  AND2X2 U11 ( .A(mem_write_data[13]), .B(n6992), .Y(n15) );
  AND2X2 U12 ( .A(mem_write_data[14]), .B(n6992), .Y(n16) );
  AND2X2 U13 ( .A(mem_write_data[15]), .B(n6992), .Y(n17) );
  NAND2X4 U14 ( .A(n486), .B(n521), .Y(n18) );
  NAND2X4 U15 ( .A(n488), .B(n521), .Y(n19) );
  NAND2X4 U16 ( .A(n490), .B(n521), .Y(n20) );
  NAND2X4 U17 ( .A(n484), .B(n521), .Y(n21) );
  NAND2X4 U18 ( .A(n567), .B(n466), .Y(n22) );
  NAND2X4 U19 ( .A(n567), .B(n519), .Y(n23) );
  NAND2X4 U20 ( .A(n537), .B(n484), .Y(n24) );
  NAND2X4 U21 ( .A(n537), .B(n486), .Y(n25) );
  NAND2X4 U22 ( .A(n537), .B(n488), .Y(n26) );
  NAND2X4 U23 ( .A(n537), .B(n490), .Y(n28) );
  NAND2X4 U24 ( .A(n537), .B(n482), .Y(n29) );
  NAND2X4 U25 ( .A(n537), .B(n468), .Y(n31) );
  NAND2X4 U26 ( .A(n537), .B(n470), .Y(n32) );
  NAND2X4 U27 ( .A(n537), .B(n472), .Y(n34) );
  NAND2X4 U28 ( .A(n537), .B(n477), .Y(n35) );
  NAND2X4 U29 ( .A(n537), .B(n478), .Y(n37) );
  NAND2X4 U30 ( .A(n537), .B(n492), .Y(n38) );
  NAND2X4 U31 ( .A(n482), .B(n521), .Y(n40) );
  NAND2X4 U32 ( .A(n468), .B(n521), .Y(n41) );
  NAND2X4 U33 ( .A(n470), .B(n521), .Y(n43) );
  NAND2X4 U34 ( .A(n472), .B(n521), .Y(n44) );
  NAND2X4 U35 ( .A(n477), .B(n521), .Y(n46) );
  NAND2X4 U36 ( .A(n478), .B(n521), .Y(n47) );
  NAND2X4 U37 ( .A(n492), .B(n521), .Y(n49) );
  NAND2X4 U38 ( .A(n480), .B(n521), .Y(n50) );
  NAND2X4 U39 ( .A(n475), .B(n521), .Y(n52) );
  NAND2X4 U40 ( .A(n517), .B(n521), .Y(n53) );
  NAND2X4 U41 ( .A(n519), .B(n521), .Y(n55) );
  NAND2X4 U42 ( .A(n523), .B(n484), .Y(n56) );
  NAND2X4 U43 ( .A(n523), .B(n486), .Y(n58) );
  NAND2X4 U44 ( .A(n523), .B(n488), .Y(n59) );
  NAND2X4 U45 ( .A(n523), .B(n490), .Y(n61) );
  NAND2X4 U46 ( .A(n523), .B(n482), .Y(n62) );
  NAND2X4 U47 ( .A(n523), .B(n468), .Y(n64) );
  NAND2X4 U48 ( .A(n523), .B(n470), .Y(n65) );
  NAND2X4 U49 ( .A(n523), .B(n472), .Y(n67) );
  NAND2X4 U50 ( .A(n523), .B(n477), .Y(n68) );
  NAND2X4 U51 ( .A(n523), .B(n478), .Y(n70) );
  NAND2X4 U52 ( .A(n523), .B(n492), .Y(n73) );
  NAND2X4 U53 ( .A(n523), .B(n480), .Y(n75) );
  NAND2X4 U54 ( .A(n523), .B(n475), .Y(n76) );
  NAND2X4 U55 ( .A(n525), .B(n484), .Y(n78) );
  NAND2X4 U56 ( .A(n525), .B(n486), .Y(n80) );
  NAND2X4 U57 ( .A(n525), .B(n488), .Y(n82) );
  NAND2X4 U58 ( .A(n525), .B(n490), .Y(n84) );
  NAND2X4 U59 ( .A(n525), .B(n482), .Y(n86) );
  NAND2X4 U60 ( .A(n525), .B(n468), .Y(n88) );
  NAND2X4 U61 ( .A(n525), .B(n470), .Y(n90) );
  NAND2X4 U62 ( .A(n525), .B(n472), .Y(n92) );
  NAND2X4 U63 ( .A(n525), .B(n477), .Y(n94) );
  NAND2X4 U64 ( .A(n525), .B(n478), .Y(n96) );
  NAND2X4 U65 ( .A(n525), .B(n480), .Y(n98) );
  NAND2X4 U66 ( .A(n525), .B(n475), .Y(n100) );
  NAND2X4 U67 ( .A(n525), .B(n517), .Y(n102) );
  NAND2X4 U68 ( .A(n525), .B(n519), .Y(n104) );
  NAND2X4 U69 ( .A(n558), .B(n484), .Y(n107) );
  NAND2X4 U70 ( .A(n558), .B(n486), .Y(n109) );
  NAND2X4 U71 ( .A(n558), .B(n488), .Y(n110) );
  NAND2X4 U72 ( .A(n558), .B(n490), .Y(n112) );
  NAND2X4 U73 ( .A(n558), .B(n482), .Y(n114) );
  NAND2X4 U74 ( .A(n558), .B(n468), .Y(n116) );
  NAND2X4 U75 ( .A(n558), .B(n470), .Y(n118) );
  NAND2X4 U76 ( .A(n558), .B(n472), .Y(n120) );
  NAND2X4 U77 ( .A(n558), .B(n477), .Y(n122) );
  NAND2X4 U78 ( .A(n558), .B(n478), .Y(n124) );
  NAND2X4 U79 ( .A(n558), .B(n492), .Y(n126) );
  NAND2X4 U80 ( .A(n558), .B(n480), .Y(n128) );
  NAND2X4 U81 ( .A(n558), .B(n475), .Y(n130) );
  NAND2X4 U82 ( .A(n558), .B(n517), .Y(n132) );
  NAND2X4 U83 ( .A(n558), .B(n519), .Y(n134) );
  NAND2X4 U84 ( .A(n527), .B(n484), .Y(n136) );
  NAND2X4 U85 ( .A(n527), .B(n486), .Y(n138) );
  NAND2X4 U86 ( .A(n527), .B(n488), .Y(n141) );
  NAND2X4 U87 ( .A(n527), .B(n490), .Y(n143) );
  NAND2X4 U88 ( .A(n527), .B(n482), .Y(n144) );
  NAND2X4 U89 ( .A(n527), .B(n468), .Y(n146) );
  NAND2X4 U90 ( .A(n527), .B(n470), .Y(n148) );
  NAND2X4 U91 ( .A(n527), .B(n472), .Y(n150) );
  NAND2X4 U92 ( .A(n527), .B(n477), .Y(n152) );
  NAND2X4 U93 ( .A(n527), .B(n478), .Y(n154) );
  NAND2X4 U94 ( .A(n527), .B(n492), .Y(n156) );
  NAND2X4 U95 ( .A(n527), .B(n480), .Y(n158) );
  NAND2X4 U96 ( .A(n527), .B(n475), .Y(n160) );
  NAND2X4 U97 ( .A(n527), .B(n517), .Y(n162) );
  NAND2X4 U98 ( .A(n527), .B(n466), .Y(n164) );
  NAND2X4 U99 ( .A(n527), .B(n519), .Y(n166) );
  NAND2X4 U100 ( .A(n529), .B(n484), .Y(n168) );
  NAND2X4 U101 ( .A(n529), .B(n486), .Y(n170) );
  NAND2X4 U102 ( .A(n529), .B(n488), .Y(n172) );
  NAND2X4 U103 ( .A(n529), .B(n490), .Y(n175) );
  NAND2X4 U104 ( .A(n529), .B(n482), .Y(n177) );
  NAND2X4 U105 ( .A(n529), .B(n468), .Y(n178) );
  NAND2X4 U106 ( .A(n529), .B(n470), .Y(n180) );
  NAND2X4 U107 ( .A(n529), .B(n472), .Y(n182) );
  NAND2X4 U108 ( .A(n529), .B(n477), .Y(n184) );
  NAND2X4 U109 ( .A(n529), .B(n478), .Y(n186) );
  NAND2X4 U110 ( .A(n529), .B(n492), .Y(n188) );
  NAND2X4 U111 ( .A(n529), .B(n480), .Y(n190) );
  NAND2X4 U112 ( .A(n529), .B(n475), .Y(n192) );
  NAND2X4 U113 ( .A(n529), .B(n517), .Y(n194) );
  NAND2X4 U114 ( .A(n529), .B(n466), .Y(n196) );
  NAND2X4 U115 ( .A(n529), .B(n519), .Y(n198) );
  NAND2X4 U116 ( .A(n539), .B(n484), .Y(n200) );
  NAND2X4 U117 ( .A(n539), .B(n486), .Y(n202) );
  NAND2X4 U118 ( .A(n539), .B(n488), .Y(n204) );
  NAND2X4 U119 ( .A(n539), .B(n490), .Y(n206) );
  NAND2X4 U120 ( .A(n539), .B(n482), .Y(n209) );
  NAND2X4 U121 ( .A(n539), .B(n468), .Y(n211) );
  NAND2X4 U122 ( .A(n539), .B(n470), .Y(n212) );
  NAND2X4 U123 ( .A(n539), .B(n472), .Y(n214) );
  NAND2X4 U124 ( .A(n539), .B(n477), .Y(n216) );
  NAND2X4 U125 ( .A(n539), .B(n478), .Y(n218) );
  NAND2X4 U126 ( .A(n539), .B(n480), .Y(n220) );
  NAND2X4 U127 ( .A(n539), .B(n475), .Y(n222) );
  NAND2X4 U128 ( .A(n539), .B(n517), .Y(n224) );
  NAND2X4 U129 ( .A(n539), .B(n466), .Y(n226) );
  NAND2X4 U130 ( .A(n539), .B(n519), .Y(n228) );
  NAND2X4 U131 ( .A(n560), .B(n484), .Y(n230) );
  NAND2X4 U132 ( .A(n560), .B(n486), .Y(n232) );
  NAND2X4 U133 ( .A(n560), .B(n488), .Y(n234) );
  NAND2X4 U134 ( .A(n560), .B(n490), .Y(n236) );
  NAND2X4 U135 ( .A(n560), .B(n482), .Y(n238) );
  NAND2X4 U136 ( .A(n560), .B(n468), .Y(n240) );
  NAND2X4 U137 ( .A(n560), .B(n470), .Y(n242) );
  NAND2X4 U138 ( .A(n560), .B(n472), .Y(n244) );
  NAND2X4 U139 ( .A(n560), .B(n477), .Y(n245) );
  NAND2X4 U140 ( .A(n560), .B(n478), .Y(n247) );
  NAND2X4 U141 ( .A(n560), .B(n492), .Y(n249) );
  NAND2X4 U142 ( .A(n560), .B(n480), .Y(n251) );
  NAND2X4 U143 ( .A(n560), .B(n475), .Y(n253) );
  NAND2X4 U144 ( .A(n560), .B(n517), .Y(n255) );
  NAND2X4 U145 ( .A(n560), .B(n466), .Y(n257) );
  NAND2X4 U146 ( .A(n560), .B(n519), .Y(n259) );
  NAND2X4 U147 ( .A(n531), .B(n484), .Y(n261) );
  NAND2X4 U148 ( .A(n531), .B(n486), .Y(n263) );
  NAND2X4 U149 ( .A(n531), .B(n488), .Y(n265) );
  NAND2X4 U150 ( .A(n531), .B(n490), .Y(n267) );
  NAND2X4 U151 ( .A(n531), .B(n482), .Y(n269) );
  NAND2X4 U152 ( .A(n531), .B(n477), .Y(n271) );
  NAND2X4 U153 ( .A(n531), .B(n478), .Y(n273) );
  NAND2X4 U154 ( .A(n531), .B(n492), .Y(n275) );
  NAND2X4 U155 ( .A(n531), .B(n480), .Y(n277) );
  NAND2X4 U156 ( .A(n531), .B(n475), .Y(n278) );
  NAND2X4 U157 ( .A(n531), .B(n517), .Y(n280) );
  NAND2X4 U158 ( .A(n531), .B(n466), .Y(n282) );
  NAND2X4 U159 ( .A(n531), .B(n519), .Y(n284) );
  NAND2X4 U160 ( .A(n562), .B(n484), .Y(n286) );
  NAND2X4 U161 ( .A(n562), .B(n486), .Y(n288) );
  NAND2X4 U162 ( .A(n562), .B(n488), .Y(n290) );
  NAND2X4 U163 ( .A(n562), .B(n490), .Y(n292) );
  NAND2X4 U164 ( .A(n562), .B(n482), .Y(n294) );
  NAND2X4 U165 ( .A(n562), .B(n477), .Y(n296) );
  NAND2X4 U166 ( .A(n562), .B(n478), .Y(n298) );
  NAND2X4 U167 ( .A(n562), .B(n492), .Y(n300) );
  NAND2X4 U168 ( .A(n562), .B(n480), .Y(n302) );
  NAND2X4 U169 ( .A(n562), .B(n475), .Y(n304) );
  NAND2X4 U170 ( .A(n562), .B(n517), .Y(n306) );
  NAND2X4 U171 ( .A(n562), .B(n466), .Y(n308) );
  NAND2X4 U172 ( .A(n562), .B(n519), .Y(n310) );
  NAND2X4 U173 ( .A(n533), .B(n484), .Y(n311) );
  NAND2X4 U174 ( .A(n533), .B(n486), .Y(n313) );
  NAND2X4 U175 ( .A(n533), .B(n488), .Y(n315) );
  NAND2X4 U176 ( .A(n533), .B(n490), .Y(n317) );
  NAND2X4 U177 ( .A(n533), .B(n482), .Y(n319) );
  NAND2X4 U178 ( .A(n533), .B(n477), .Y(n321) );
  NAND2X4 U179 ( .A(n533), .B(n478), .Y(n323) );
  NAND2X4 U180 ( .A(n533), .B(n480), .Y(n325) );
  NAND2X4 U181 ( .A(n533), .B(n475), .Y(n327) );
  NAND2X4 U182 ( .A(n533), .B(n517), .Y(n329) );
  NAND2X4 U183 ( .A(n533), .B(n466), .Y(n331) );
  NAND2X4 U184 ( .A(n533), .B(n519), .Y(n333) );
  NAND2X4 U185 ( .A(n564), .B(n484), .Y(n335) );
  NAND2X4 U186 ( .A(n564), .B(n486), .Y(n337) );
  NAND2X4 U187 ( .A(n564), .B(n488), .Y(n339) );
  NAND2X4 U188 ( .A(n564), .B(n490), .Y(n342) );
  NAND2X4 U189 ( .A(n564), .B(n482), .Y(n344) );
  NAND2X4 U190 ( .A(n564), .B(n477), .Y(n345) );
  NAND2X4 U191 ( .A(n564), .B(n478), .Y(n347) );
  NAND2X4 U192 ( .A(n564), .B(n492), .Y(n349) );
  NAND2X4 U193 ( .A(n564), .B(n480), .Y(n351) );
  NAND2X4 U194 ( .A(n564), .B(n475), .Y(n353) );
  NAND2X4 U195 ( .A(n564), .B(n517), .Y(n355) );
  NAND2X4 U196 ( .A(n564), .B(n466), .Y(n357) );
  NAND2X4 U197 ( .A(n564), .B(n519), .Y(n359) );
  NAND2X4 U198 ( .A(n535), .B(n484), .Y(n361) );
  NAND2X4 U199 ( .A(n535), .B(n486), .Y(n363) );
  NAND2X4 U200 ( .A(n535), .B(n488), .Y(n365) );
  NAND2X4 U201 ( .A(n535), .B(n490), .Y(n367) );
  NAND2X4 U202 ( .A(n535), .B(n482), .Y(n369) );
  NAND2X4 U203 ( .A(n535), .B(n468), .Y(n371) );
  NAND2X4 U204 ( .A(n535), .B(n470), .Y(n373) );
  NAND2X4 U205 ( .A(n535), .B(n472), .Y(n375) );
  NAND2X4 U206 ( .A(n535), .B(n477), .Y(n377) );
  NAND2X4 U207 ( .A(n535), .B(n478), .Y(n378) );
  NAND2X4 U208 ( .A(n535), .B(n492), .Y(n380) );
  NAND2X4 U209 ( .A(n535), .B(n480), .Y(n382) );
  NAND2X4 U210 ( .A(n535), .B(n475), .Y(n384) );
  NAND2X4 U211 ( .A(n535), .B(n517), .Y(n386) );
  NAND2X4 U212 ( .A(n535), .B(n466), .Y(n388) );
  NAND2X4 U213 ( .A(n535), .B(n519), .Y(n390) );
  NAND2X4 U214 ( .A(n567), .B(n484), .Y(n392) );
  NAND2X4 U215 ( .A(n567), .B(n486), .Y(n394) );
  NAND2X4 U216 ( .A(n567), .B(n488), .Y(n396) );
  NAND2X4 U217 ( .A(n567), .B(n490), .Y(n398) );
  NAND2X4 U218 ( .A(n567), .B(n482), .Y(n400) );
  NAND2X4 U219 ( .A(n567), .B(n468), .Y(n402) );
  NAND2X4 U220 ( .A(n567), .B(n470), .Y(n404) );
  NAND2X4 U221 ( .A(n567), .B(n472), .Y(n406) );
  NAND2X4 U222 ( .A(n567), .B(n477), .Y(n408) );
  NAND2X4 U223 ( .A(n567), .B(n478), .Y(n410) );
  NAND2X4 U224 ( .A(n567), .B(n492), .Y(n411) );
  NAND2X4 U225 ( .A(n567), .B(n480), .Y(n413) );
  NAND2X4 U226 ( .A(n567), .B(n475), .Y(n415) );
  NAND2X4 U227 ( .A(n567), .B(n517), .Y(n417) );
  NAND2X4 U228 ( .A(n537), .B(n480), .Y(n419) );
  NAND2X4 U229 ( .A(n537), .B(n475), .Y(n421) );
  NAND2X4 U230 ( .A(n537), .B(n517), .Y(n423) );
  NAND2X4 U231 ( .A(n537), .B(n466), .Y(n425) );
  NAND2X4 U232 ( .A(n537), .B(n519), .Y(n427) );
  NAND2X4 U233 ( .A(n569), .B(n484), .Y(n429) );
  NAND2X4 U234 ( .A(n569), .B(n486), .Y(n431) );
  NAND2X4 U235 ( .A(n569), .B(n488), .Y(n433) );
  NAND2X4 U236 ( .A(n569), .B(n490), .Y(n435) );
  NAND2X4 U237 ( .A(n569), .B(n482), .Y(n437) );
  NAND2X4 U238 ( .A(n569), .B(n468), .Y(n439) );
  NAND2X4 U239 ( .A(n569), .B(n470), .Y(n441) );
  NAND2X4 U240 ( .A(n569), .B(n472), .Y(n443) );
  NAND2X4 U241 ( .A(n569), .B(n477), .Y(n444) );
  NAND2X4 U242 ( .A(n569), .B(n478), .Y(n446) );
  NAND2X4 U243 ( .A(n569), .B(n492), .Y(n448) );
  NAND2X4 U244 ( .A(n569), .B(n480), .Y(n450) );
  NAND2X4 U245 ( .A(n569), .B(n475), .Y(n452) );
  NAND2X4 U246 ( .A(n569), .B(n517), .Y(n454) );
  NAND2X4 U247 ( .A(n569), .B(n466), .Y(n456) );
  NAND2X4 U248 ( .A(n569), .B(n519), .Y(n458) );
  NAND2X4 U249 ( .A(n525), .B(n492), .Y(n460) );
  NAND2X4 U250 ( .A(n539), .B(n492), .Y(n462) );
  NAND2X4 U251 ( .A(n533), .B(n492), .Y(n464) );
  AND2X4 U252 ( .A(n575), .B(n551), .Y(n466) );
  AND2X4 U253 ( .A(n557), .B(n548), .Y(n468) );
  AND2X4 U254 ( .A(n557), .B(n551), .Y(n470) );
  AND2X4 U255 ( .A(n557), .B(n554), .Y(n472) );
  AND2X4 U256 ( .A(n575), .B(n545), .Y(n475) );
  AND2X4 U257 ( .A(n566), .B(n545), .Y(n477) );
  AND2X4 U258 ( .A(n566), .B(n548), .Y(n478) );
  AND2X4 U259 ( .A(n566), .B(n554), .Y(n480) );
  AND2X4 U260 ( .A(n557), .B(n545), .Y(n482) );
  AND2X4 U261 ( .A(n544), .B(n545), .Y(n484) );
  AND2X4 U262 ( .A(n548), .B(n544), .Y(n486) );
  AND2X4 U263 ( .A(n551), .B(n544), .Y(n488) );
  AND2X4 U264 ( .A(n554), .B(n544), .Y(n490) );
  AND2X4 U265 ( .A(n566), .B(n551), .Y(n492) );
  NAND2X4 U266 ( .A(n466), .B(n521), .Y(n494) );
  NAND2X4 U267 ( .A(n525), .B(n466), .Y(n496) );
  NAND2X4 U268 ( .A(n558), .B(n466), .Y(n498) );
  NAND2X4 U269 ( .A(n531), .B(n468), .Y(n500) );
  NAND2X4 U270 ( .A(n531), .B(n470), .Y(n502) );
  NAND2X4 U271 ( .A(n531), .B(n472), .Y(n504) );
  NAND2X4 U272 ( .A(n562), .B(n468), .Y(n506) );
  NAND2X4 U273 ( .A(n562), .B(n470), .Y(n508) );
  NAND2X4 U274 ( .A(n562), .B(n472), .Y(n510) );
  NAND2X4 U275 ( .A(n564), .B(n468), .Y(n511) );
  NAND2X4 U276 ( .A(n564), .B(n470), .Y(n513) );
  NAND2X4 U277 ( .A(n564), .B(n472), .Y(n515) );
  AND2X4 U278 ( .A(n575), .B(n548), .Y(n517) );
  AND2X4 U279 ( .A(n575), .B(n554), .Y(n519) );
  AND2X4 U280 ( .A(n71), .B(n72), .Y(n521) );
  AND2X4 U281 ( .A(n106), .B(n71), .Y(n523) );
  AND2X4 U282 ( .A(n140), .B(n71), .Y(n525) );
  AND2X4 U283 ( .A(n208), .B(n72), .Y(n527) );
  AND2X4 U284 ( .A(n208), .B(n106), .Y(n529) );
  AND2X4 U285 ( .A(n341), .B(n72), .Y(n531) );
  AND2X4 U286 ( .A(n341), .B(n140), .Y(n533) );
  AND2X4 U287 ( .A(n474), .B(n72), .Y(n535) );
  AND2X4 U288 ( .A(n474), .B(n140), .Y(n537) );
  AND2X4 U289 ( .A(n208), .B(n140), .Y(n539) );
  NAND2X4 U290 ( .A(n523), .B(n517), .Y(n541) );
  NAND2X4 U291 ( .A(n523), .B(n466), .Y(n543) );
  NAND2X4 U292 ( .A(n523), .B(n519), .Y(n546) );
  NAND2X4 U293 ( .A(n533), .B(n468), .Y(n549) );
  NAND2X4 U294 ( .A(n533), .B(n470), .Y(n552) );
  NAND2X4 U295 ( .A(n533), .B(n472), .Y(n555) );
  AND2X4 U296 ( .A(n174), .B(n71), .Y(n558) );
  AND2X4 U297 ( .A(n208), .B(n174), .Y(n560) );
  AND2X4 U298 ( .A(n341), .B(n106), .Y(n562) );
  AND2X4 U299 ( .A(n341), .B(n174), .Y(n564) );
  AND2X4 U300 ( .A(n474), .B(n106), .Y(n567) );
  AND2X4 U301 ( .A(n474), .B(n174), .Y(n569) );
  OAI2BB2XL U302 ( .B0(n6962), .B1(n18), .A0N(\ram[1][0] ), .A1N(n6609), .Y(
        n598) );
  OAI2BB2XL U303 ( .B0(n6939), .B1(n18), .A0N(\ram[1][1] ), .A1N(n6609), .Y(
        n599) );
  OAI2BB2XL U304 ( .B0(n6916), .B1(n18), .A0N(\ram[1][2] ), .A1N(n6609), .Y(
        n600) );
  OAI2BB2XL U305 ( .B0(n6893), .B1(n18), .A0N(\ram[1][3] ), .A1N(n6609), .Y(
        n601) );
  OAI2BB2XL U306 ( .B0(n6879), .B1(n18), .A0N(\ram[1][4] ), .A1N(n6609), .Y(
        n602) );
  OAI2BB2XL U307 ( .B0(n6856), .B1(n18), .A0N(\ram[1][5] ), .A1N(n6609), .Y(
        n603) );
  OAI2BB2XL U308 ( .B0(n6833), .B1(n18), .A0N(\ram[1][6] ), .A1N(n6609), .Y(
        n604) );
  OAI2BB2XL U309 ( .B0(n6810), .B1(n18), .A0N(\ram[1][7] ), .A1N(n6609), .Y(
        n605) );
  OAI2BB2XL U310 ( .B0(n6787), .B1(n18), .A0N(\ram[1][8] ), .A1N(n6609), .Y(
        n606) );
  OAI2BB2XL U311 ( .B0(n6764), .B1(n18), .A0N(\ram[1][9] ), .A1N(n6609), .Y(
        n607) );
  OAI2BB2XL U312 ( .B0(n6741), .B1(n18), .A0N(\ram[1][10] ), .A1N(n6609), .Y(
        n608) );
  OAI2BB2XL U313 ( .B0(n6718), .B1(n18), .A0N(\ram[1][11] ), .A1N(n6609), .Y(
        n609) );
  OAI2BB2XL U314 ( .B0(n6695), .B1(n18), .A0N(\ram[1][12] ), .A1N(n6609), .Y(
        n610) );
  OAI2BB2XL U315 ( .B0(n6672), .B1(n18), .A0N(\ram[1][13] ), .A1N(n6609), .Y(
        n611) );
  OAI2BB2XL U316 ( .B0(n6649), .B1(n18), .A0N(\ram[1][14] ), .A1N(n6609), .Y(
        n612) );
  OAI2BB2XL U317 ( .B0(n6626), .B1(n18), .A0N(\ram[1][15] ), .A1N(n6609), .Y(
        n613) );
  OAI2BB2XL U318 ( .B0(n6961), .B1(n19), .A0N(\ram[2][0] ), .A1N(n6608), .Y(
        n614) );
  OAI2BB2XL U319 ( .B0(n6938), .B1(n19), .A0N(\ram[2][1] ), .A1N(n6608), .Y(
        n615) );
  OAI2BB2XL U320 ( .B0(n6915), .B1(n19), .A0N(\ram[2][2] ), .A1N(n6608), .Y(
        n616) );
  OAI2BB2XL U321 ( .B0(n6892), .B1(n19), .A0N(\ram[2][3] ), .A1N(n6608), .Y(
        n617) );
  OAI2BB2XL U322 ( .B0(n6878), .B1(n19), .A0N(\ram[2][4] ), .A1N(n6608), .Y(
        n618) );
  OAI2BB2XL U323 ( .B0(n6855), .B1(n19), .A0N(\ram[2][5] ), .A1N(n6608), .Y(
        n619) );
  OAI2BB2XL U324 ( .B0(n6832), .B1(n19), .A0N(\ram[2][6] ), .A1N(n6608), .Y(
        n620) );
  OAI2BB2XL U325 ( .B0(n6809), .B1(n19), .A0N(\ram[2][7] ), .A1N(n6608), .Y(
        n621) );
  OAI2BB2XL U326 ( .B0(n6786), .B1(n19), .A0N(\ram[2][8] ), .A1N(n6608), .Y(
        n622) );
  OAI2BB2XL U327 ( .B0(n6763), .B1(n19), .A0N(\ram[2][9] ), .A1N(n6608), .Y(
        n623) );
  OAI2BB2XL U328 ( .B0(n6740), .B1(n19), .A0N(\ram[2][10] ), .A1N(n6608), .Y(
        n624) );
  OAI2BB2XL U329 ( .B0(n6717), .B1(n19), .A0N(\ram[2][11] ), .A1N(n6608), .Y(
        n625) );
  OAI2BB2XL U330 ( .B0(n6694), .B1(n19), .A0N(\ram[2][12] ), .A1N(n6608), .Y(
        n626) );
  OAI2BB2XL U331 ( .B0(n6671), .B1(n19), .A0N(\ram[2][13] ), .A1N(n6608), .Y(
        n627) );
  OAI2BB2XL U332 ( .B0(n6648), .B1(n19), .A0N(\ram[2][14] ), .A1N(n6608), .Y(
        n628) );
  OAI2BB2XL U333 ( .B0(n6625), .B1(n19), .A0N(\ram[2][15] ), .A1N(n6608), .Y(
        n629) );
  OAI2BB2XL U334 ( .B0(n6961), .B1(n20), .A0N(\ram[3][0] ), .A1N(n6607), .Y(
        n630) );
  OAI2BB2XL U335 ( .B0(n6938), .B1(n20), .A0N(\ram[3][1] ), .A1N(n6607), .Y(
        n631) );
  OAI2BB2XL U336 ( .B0(n6915), .B1(n20), .A0N(\ram[3][2] ), .A1N(n6607), .Y(
        n632) );
  OAI2BB2XL U337 ( .B0(n6892), .B1(n20), .A0N(\ram[3][3] ), .A1N(n6607), .Y(
        n633) );
  OAI2BB2XL U338 ( .B0(n6879), .B1(n20), .A0N(\ram[3][4] ), .A1N(n6607), .Y(
        n634) );
  OAI2BB2XL U339 ( .B0(n6856), .B1(n20), .A0N(\ram[3][5] ), .A1N(n6607), .Y(
        n635) );
  OAI2BB2XL U340 ( .B0(n6833), .B1(n20), .A0N(\ram[3][6] ), .A1N(n6607), .Y(
        n636) );
  OAI2BB2XL U341 ( .B0(n6810), .B1(n20), .A0N(\ram[3][7] ), .A1N(n6607), .Y(
        n637) );
  OAI2BB2XL U342 ( .B0(n6787), .B1(n20), .A0N(\ram[3][8] ), .A1N(n6607), .Y(
        n638) );
  OAI2BB2XL U343 ( .B0(n6764), .B1(n20), .A0N(\ram[3][9] ), .A1N(n6607), .Y(
        n639) );
  OAI2BB2XL U344 ( .B0(n6741), .B1(n20), .A0N(\ram[3][10] ), .A1N(n6607), .Y(
        n640) );
  OAI2BB2XL U345 ( .B0(n6718), .B1(n20), .A0N(\ram[3][11] ), .A1N(n6607), .Y(
        n641) );
  OAI2BB2XL U346 ( .B0(n6695), .B1(n20), .A0N(\ram[3][12] ), .A1N(n6607), .Y(
        n642) );
  OAI2BB2XL U347 ( .B0(n6672), .B1(n20), .A0N(\ram[3][13] ), .A1N(n6607), .Y(
        n643) );
  OAI2BB2XL U348 ( .B0(n6649), .B1(n20), .A0N(\ram[3][14] ), .A1N(n6607), .Y(
        n644) );
  OAI2BB2XL U349 ( .B0(n6626), .B1(n20), .A0N(\ram[3][15] ), .A1N(n6607), .Y(
        n645) );
  OAI2BB2XL U350 ( .B0(n6972), .B1(n40), .A0N(\ram[4][0] ), .A1N(n6606), .Y(
        n646) );
  OAI2BB2XL U351 ( .B0(n6949), .B1(n40), .A0N(\ram[4][1] ), .A1N(n6606), .Y(
        n647) );
  OAI2BB2XL U352 ( .B0(n6926), .B1(n40), .A0N(\ram[4][2] ), .A1N(n6606), .Y(
        n648) );
  OAI2BB2XL U353 ( .B0(n6903), .B1(n40), .A0N(\ram[4][3] ), .A1N(n6606), .Y(
        n649) );
  OAI2BB2XL U354 ( .B0(n6882), .B1(n40), .A0N(\ram[4][4] ), .A1N(n6606), .Y(
        n650) );
  OAI2BB2XL U355 ( .B0(n6859), .B1(n40), .A0N(\ram[4][5] ), .A1N(n6606), .Y(
        n651) );
  OAI2BB2XL U356 ( .B0(n6836), .B1(n40), .A0N(\ram[4][6] ), .A1N(n6606), .Y(
        n652) );
  OAI2BB2XL U357 ( .B0(n6813), .B1(n40), .A0N(\ram[4][7] ), .A1N(n6606), .Y(
        n653) );
  OAI2BB2XL U358 ( .B0(n6790), .B1(n40), .A0N(\ram[4][8] ), .A1N(n6606), .Y(
        n654) );
  OAI2BB2XL U359 ( .B0(n6767), .B1(n40), .A0N(\ram[4][9] ), .A1N(n6606), .Y(
        n655) );
  OAI2BB2XL U360 ( .B0(n6744), .B1(n40), .A0N(\ram[4][10] ), .A1N(n6606), .Y(
        n656) );
  OAI2BB2XL U361 ( .B0(n6721), .B1(n40), .A0N(\ram[4][11] ), .A1N(n6606), .Y(
        n657) );
  OAI2BB2XL U362 ( .B0(n6698), .B1(n40), .A0N(\ram[4][12] ), .A1N(n6606), .Y(
        n658) );
  OAI2BB2XL U363 ( .B0(n6675), .B1(n40), .A0N(\ram[4][13] ), .A1N(n6606), .Y(
        n659) );
  OAI2BB2XL U364 ( .B0(n6652), .B1(n40), .A0N(\ram[4][14] ), .A1N(n6606), .Y(
        n660) );
  OAI2BB2XL U365 ( .B0(n6629), .B1(n40), .A0N(\ram[4][15] ), .A1N(n6606), .Y(
        n661) );
  OAI2BB2XL U366 ( .B0(n6971), .B1(n46), .A0N(\ram[8][0] ), .A1N(n6602), .Y(
        n710) );
  OAI2BB2XL U367 ( .B0(n6948), .B1(n46), .A0N(\ram[8][1] ), .A1N(n6602), .Y(
        n711) );
  OAI2BB2XL U368 ( .B0(n6925), .B1(n46), .A0N(\ram[8][2] ), .A1N(n6602), .Y(
        n712) );
  OAI2BB2XL U369 ( .B0(n6902), .B1(n46), .A0N(\ram[8][3] ), .A1N(n6602), .Y(
        n713) );
  OAI2BB2XL U370 ( .B0(n6882), .B1(n46), .A0N(\ram[8][4] ), .A1N(n6602), .Y(
        n714) );
  OAI2BB2XL U371 ( .B0(n6859), .B1(n46), .A0N(\ram[8][5] ), .A1N(n6602), .Y(
        n715) );
  OAI2BB2XL U372 ( .B0(n6836), .B1(n46), .A0N(\ram[8][6] ), .A1N(n6602), .Y(
        n716) );
  OAI2BB2XL U373 ( .B0(n6813), .B1(n46), .A0N(\ram[8][7] ), .A1N(n6602), .Y(
        n717) );
  OAI2BB2XL U374 ( .B0(n6790), .B1(n46), .A0N(\ram[8][8] ), .A1N(n6602), .Y(
        n718) );
  OAI2BB2XL U375 ( .B0(n6767), .B1(n46), .A0N(\ram[8][9] ), .A1N(n6602), .Y(
        n719) );
  OAI2BB2XL U376 ( .B0(n6744), .B1(n46), .A0N(\ram[8][10] ), .A1N(n6602), .Y(
        n720) );
  OAI2BB2XL U377 ( .B0(n6721), .B1(n46), .A0N(\ram[8][11] ), .A1N(n6602), .Y(
        n721) );
  OAI2BB2XL U378 ( .B0(n6698), .B1(n46), .A0N(\ram[8][12] ), .A1N(n6602), .Y(
        n722) );
  OAI2BB2XL U379 ( .B0(n6675), .B1(n46), .A0N(\ram[8][13] ), .A1N(n6602), .Y(
        n723) );
  OAI2BB2XL U380 ( .B0(n6652), .B1(n46), .A0N(\ram[8][14] ), .A1N(n6602), .Y(
        n724) );
  OAI2BB2XL U381 ( .B0(n6629), .B1(n46), .A0N(\ram[8][15] ), .A1N(n6602), .Y(
        n725) );
  OAI2BB2XL U382 ( .B0(n6970), .B1(n52), .A0N(\ram[12][0] ), .A1N(n6598), .Y(
        n774) );
  OAI2BB2XL U383 ( .B0(n6947), .B1(n52), .A0N(\ram[12][1] ), .A1N(n6598), .Y(
        n775) );
  OAI2BB2XL U384 ( .B0(n6924), .B1(n52), .A0N(\ram[12][2] ), .A1N(n6598), .Y(
        n776) );
  OAI2BB2XL U385 ( .B0(n6901), .B1(n52), .A0N(\ram[12][3] ), .A1N(n6598), .Y(
        n777) );
  OAI2BB2XL U386 ( .B0(n6882), .B1(n52), .A0N(\ram[12][4] ), .A1N(n6598), .Y(
        n778) );
  OAI2BB2XL U387 ( .B0(n6859), .B1(n52), .A0N(\ram[12][5] ), .A1N(n6598), .Y(
        n779) );
  OAI2BB2XL U388 ( .B0(n6836), .B1(n52), .A0N(\ram[12][6] ), .A1N(n6598), .Y(
        n780) );
  OAI2BB2XL U389 ( .B0(n6813), .B1(n52), .A0N(\ram[12][7] ), .A1N(n6598), .Y(
        n781) );
  OAI2BB2XL U390 ( .B0(n6790), .B1(n52), .A0N(\ram[12][8] ), .A1N(n6598), .Y(
        n782) );
  OAI2BB2XL U391 ( .B0(n6767), .B1(n52), .A0N(\ram[12][9] ), .A1N(n6598), .Y(
        n783) );
  OAI2BB2XL U392 ( .B0(n6744), .B1(n52), .A0N(\ram[12][10] ), .A1N(n6598), .Y(
        n784) );
  OAI2BB2XL U393 ( .B0(n6721), .B1(n52), .A0N(\ram[12][11] ), .A1N(n6598), .Y(
        n785) );
  OAI2BB2XL U394 ( .B0(n6698), .B1(n52), .A0N(\ram[12][12] ), .A1N(n6598), .Y(
        n786) );
  OAI2BB2XL U395 ( .B0(n6675), .B1(n52), .A0N(\ram[12][13] ), .A1N(n6598), .Y(
        n787) );
  OAI2BB2XL U396 ( .B0(n6652), .B1(n52), .A0N(\ram[12][14] ), .A1N(n6598), .Y(
        n788) );
  OAI2BB2XL U397 ( .B0(n6629), .B1(n52), .A0N(\ram[12][15] ), .A1N(n6598), .Y(
        n789) );
  OAI2BB2XL U398 ( .B0(n6974), .B1(n136), .A0N(\ram[64][0] ), .A1N(n6546), .Y(
        n1606) );
  OAI2BB2XL U399 ( .B0(n6951), .B1(n136), .A0N(\ram[64][1] ), .A1N(n6546), .Y(
        n1607) );
  OAI2BB2XL U400 ( .B0(n6928), .B1(n136), .A0N(\ram[64][2] ), .A1N(n6546), .Y(
        n1608) );
  OAI2BB2XL U401 ( .B0(n6905), .B1(n136), .A0N(\ram[64][3] ), .A1N(n6546), .Y(
        n1609) );
  OAI2BB2XL U402 ( .B0(n6877), .B1(n136), .A0N(\ram[64][4] ), .A1N(n6546), .Y(
        n1610) );
  OAI2BB2XL U403 ( .B0(n6854), .B1(n136), .A0N(\ram[64][5] ), .A1N(n6546), .Y(
        n1611) );
  OAI2BB2XL U404 ( .B0(n6831), .B1(n136), .A0N(\ram[64][6] ), .A1N(n6546), .Y(
        n1612) );
  OAI2BB2XL U405 ( .B0(n6808), .B1(n136), .A0N(\ram[64][7] ), .A1N(n6546), .Y(
        n1613) );
  OAI2BB2XL U406 ( .B0(n6785), .B1(n136), .A0N(\ram[64][8] ), .A1N(n6546), .Y(
        n1614) );
  OAI2BB2XL U407 ( .B0(n6762), .B1(n136), .A0N(\ram[64][9] ), .A1N(n6546), .Y(
        n1615) );
  OAI2BB2XL U408 ( .B0(n6739), .B1(n136), .A0N(\ram[64][10] ), .A1N(n6546), 
        .Y(n1616) );
  OAI2BB2XL U409 ( .B0(n6716), .B1(n136), .A0N(\ram[64][11] ), .A1N(n6546), 
        .Y(n1617) );
  OAI2BB2XL U410 ( .B0(n6693), .B1(n136), .A0N(\ram[64][12] ), .A1N(n6546), 
        .Y(n1618) );
  OAI2BB2XL U411 ( .B0(n6670), .B1(n136), .A0N(\ram[64][13] ), .A1N(n6546), 
        .Y(n1619) );
  OAI2BB2XL U412 ( .B0(n6647), .B1(n136), .A0N(\ram[64][14] ), .A1N(n6546), 
        .Y(n1620) );
  OAI2BB2XL U413 ( .B0(n6624), .B1(n136), .A0N(\ram[64][15] ), .A1N(n6546), 
        .Y(n1621) );
  OAI2BB2XL U414 ( .B0(n6974), .B1(n138), .A0N(\ram[65][0] ), .A1N(n6545), .Y(
        n1622) );
  OAI2BB2XL U415 ( .B0(n6951), .B1(n138), .A0N(\ram[65][1] ), .A1N(n6545), .Y(
        n1623) );
  OAI2BB2XL U416 ( .B0(n6928), .B1(n138), .A0N(\ram[65][2] ), .A1N(n6545), .Y(
        n1624) );
  OAI2BB2XL U417 ( .B0(n6905), .B1(n138), .A0N(\ram[65][3] ), .A1N(n6545), .Y(
        n1625) );
  OAI2BB2XL U418 ( .B0(n6877), .B1(n138), .A0N(\ram[65][4] ), .A1N(n6545), .Y(
        n1626) );
  OAI2BB2XL U419 ( .B0(n6854), .B1(n138), .A0N(\ram[65][5] ), .A1N(n6545), .Y(
        n1627) );
  OAI2BB2XL U420 ( .B0(n6831), .B1(n138), .A0N(\ram[65][6] ), .A1N(n6545), .Y(
        n1628) );
  OAI2BB2XL U421 ( .B0(n6808), .B1(n138), .A0N(\ram[65][7] ), .A1N(n6545), .Y(
        n1629) );
  OAI2BB2XL U422 ( .B0(n6785), .B1(n138), .A0N(\ram[65][8] ), .A1N(n6545), .Y(
        n1630) );
  OAI2BB2XL U423 ( .B0(n6762), .B1(n138), .A0N(\ram[65][9] ), .A1N(n6545), .Y(
        n1631) );
  OAI2BB2XL U424 ( .B0(n6739), .B1(n138), .A0N(\ram[65][10] ), .A1N(n6545), 
        .Y(n1632) );
  OAI2BB2XL U425 ( .B0(n6716), .B1(n138), .A0N(\ram[65][11] ), .A1N(n6545), 
        .Y(n1633) );
  OAI2BB2XL U426 ( .B0(n6693), .B1(n138), .A0N(\ram[65][12] ), .A1N(n6545), 
        .Y(n1634) );
  OAI2BB2XL U427 ( .B0(n6670), .B1(n138), .A0N(\ram[65][13] ), .A1N(n6545), 
        .Y(n1635) );
  OAI2BB2XL U428 ( .B0(n6647), .B1(n138), .A0N(\ram[65][14] ), .A1N(n6545), 
        .Y(n1636) );
  OAI2BB2XL U429 ( .B0(n6624), .B1(n138), .A0N(\ram[65][15] ), .A1N(n6545), 
        .Y(n1637) );
  OAI2BB2XL U430 ( .B0(n6974), .B1(n141), .A0N(\ram[66][0] ), .A1N(n6544), .Y(
        n1638) );
  OAI2BB2XL U431 ( .B0(n6951), .B1(n141), .A0N(\ram[66][1] ), .A1N(n6544), .Y(
        n1639) );
  OAI2BB2XL U432 ( .B0(n6928), .B1(n141), .A0N(\ram[66][2] ), .A1N(n6544), .Y(
        n1640) );
  OAI2BB2XL U433 ( .B0(n6905), .B1(n141), .A0N(\ram[66][3] ), .A1N(n6544), .Y(
        n1641) );
  OAI2BB2XL U434 ( .B0(n6877), .B1(n141), .A0N(\ram[66][4] ), .A1N(n6544), .Y(
        n1642) );
  OAI2BB2XL U435 ( .B0(n6854), .B1(n141), .A0N(\ram[66][5] ), .A1N(n6544), .Y(
        n1643) );
  OAI2BB2XL U436 ( .B0(n6831), .B1(n141), .A0N(\ram[66][6] ), .A1N(n6544), .Y(
        n1644) );
  OAI2BB2XL U437 ( .B0(n6808), .B1(n141), .A0N(\ram[66][7] ), .A1N(n6544), .Y(
        n1645) );
  OAI2BB2XL U438 ( .B0(n6785), .B1(n141), .A0N(\ram[66][8] ), .A1N(n6544), .Y(
        n1646) );
  OAI2BB2XL U439 ( .B0(n6762), .B1(n141), .A0N(\ram[66][9] ), .A1N(n6544), .Y(
        n1647) );
  OAI2BB2XL U440 ( .B0(n6739), .B1(n141), .A0N(\ram[66][10] ), .A1N(n6544), 
        .Y(n1648) );
  OAI2BB2XL U441 ( .B0(n6716), .B1(n141), .A0N(\ram[66][11] ), .A1N(n6544), 
        .Y(n1649) );
  OAI2BB2XL U442 ( .B0(n6693), .B1(n141), .A0N(\ram[66][12] ), .A1N(n6544), 
        .Y(n1650) );
  OAI2BB2XL U443 ( .B0(n6670), .B1(n141), .A0N(\ram[66][13] ), .A1N(n6544), 
        .Y(n1651) );
  OAI2BB2XL U444 ( .B0(n6647), .B1(n141), .A0N(\ram[66][14] ), .A1N(n6544), 
        .Y(n1652) );
  OAI2BB2XL U445 ( .B0(n6624), .B1(n141), .A0N(\ram[66][15] ), .A1N(n6544), 
        .Y(n1653) );
  OAI2BB2XL U446 ( .B0(n6974), .B1(n143), .A0N(\ram[67][0] ), .A1N(n6543), .Y(
        n1654) );
  OAI2BB2XL U447 ( .B0(n6951), .B1(n143), .A0N(\ram[67][1] ), .A1N(n6543), .Y(
        n1655) );
  OAI2BB2XL U448 ( .B0(n6928), .B1(n143), .A0N(\ram[67][2] ), .A1N(n6543), .Y(
        n1656) );
  OAI2BB2XL U449 ( .B0(n6905), .B1(n143), .A0N(\ram[67][3] ), .A1N(n6543), .Y(
        n1657) );
  OAI2BB2XL U450 ( .B0(n6877), .B1(n143), .A0N(\ram[67][4] ), .A1N(n6543), .Y(
        n1658) );
  OAI2BB2XL U451 ( .B0(n6854), .B1(n143), .A0N(\ram[67][5] ), .A1N(n6543), .Y(
        n1659) );
  OAI2BB2XL U452 ( .B0(n6831), .B1(n143), .A0N(\ram[67][6] ), .A1N(n6543), .Y(
        n1660) );
  OAI2BB2XL U453 ( .B0(n6808), .B1(n143), .A0N(\ram[67][7] ), .A1N(n6543), .Y(
        n1661) );
  OAI2BB2XL U454 ( .B0(n6785), .B1(n143), .A0N(\ram[67][8] ), .A1N(n6543), .Y(
        n1662) );
  OAI2BB2XL U455 ( .B0(n6762), .B1(n143), .A0N(\ram[67][9] ), .A1N(n6543), .Y(
        n1663) );
  OAI2BB2XL U456 ( .B0(n6739), .B1(n143), .A0N(\ram[67][10] ), .A1N(n6543), 
        .Y(n1664) );
  OAI2BB2XL U457 ( .B0(n6716), .B1(n143), .A0N(\ram[67][11] ), .A1N(n6543), 
        .Y(n1665) );
  OAI2BB2XL U458 ( .B0(n6693), .B1(n143), .A0N(\ram[67][12] ), .A1N(n6543), 
        .Y(n1666) );
  OAI2BB2XL U459 ( .B0(n6670), .B1(n143), .A0N(\ram[67][13] ), .A1N(n6543), 
        .Y(n1667) );
  OAI2BB2XL U460 ( .B0(n6647), .B1(n143), .A0N(\ram[67][14] ), .A1N(n6543), 
        .Y(n1668) );
  OAI2BB2XL U461 ( .B0(n6624), .B1(n143), .A0N(\ram[67][15] ), .A1N(n6543), 
        .Y(n1669) );
  OAI2BB2XL U462 ( .B0(n6974), .B1(n144), .A0N(\ram[68][0] ), .A1N(n6542), .Y(
        n1670) );
  OAI2BB2XL U463 ( .B0(n6951), .B1(n144), .A0N(\ram[68][1] ), .A1N(n6542), .Y(
        n1671) );
  OAI2BB2XL U464 ( .B0(n6928), .B1(n144), .A0N(\ram[68][2] ), .A1N(n6542), .Y(
        n1672) );
  OAI2BB2XL U465 ( .B0(n6905), .B1(n144), .A0N(\ram[68][3] ), .A1N(n6542), .Y(
        n1673) );
  OAI2BB2XL U466 ( .B0(n6877), .B1(n144), .A0N(\ram[68][4] ), .A1N(n6542), .Y(
        n1674) );
  OAI2BB2XL U467 ( .B0(n6854), .B1(n144), .A0N(\ram[68][5] ), .A1N(n6542), .Y(
        n1675) );
  OAI2BB2XL U468 ( .B0(n6831), .B1(n144), .A0N(\ram[68][6] ), .A1N(n6542), .Y(
        n1676) );
  OAI2BB2XL U469 ( .B0(n6808), .B1(n144), .A0N(\ram[68][7] ), .A1N(n6542), .Y(
        n1677) );
  OAI2BB2XL U470 ( .B0(n6785), .B1(n144), .A0N(\ram[68][8] ), .A1N(n6542), .Y(
        n1678) );
  OAI2BB2XL U471 ( .B0(n6762), .B1(n144), .A0N(\ram[68][9] ), .A1N(n6542), .Y(
        n1679) );
  OAI2BB2XL U472 ( .B0(n6739), .B1(n144), .A0N(\ram[68][10] ), .A1N(n6542), 
        .Y(n1680) );
  OAI2BB2XL U473 ( .B0(n6716), .B1(n144), .A0N(\ram[68][11] ), .A1N(n6542), 
        .Y(n1681) );
  OAI2BB2XL U474 ( .B0(n6693), .B1(n144), .A0N(\ram[68][12] ), .A1N(n6542), 
        .Y(n1682) );
  OAI2BB2XL U475 ( .B0(n6670), .B1(n144), .A0N(\ram[68][13] ), .A1N(n6542), 
        .Y(n1683) );
  OAI2BB2XL U476 ( .B0(n6647), .B1(n144), .A0N(\ram[68][14] ), .A1N(n6542), 
        .Y(n1684) );
  OAI2BB2XL U477 ( .B0(n6624), .B1(n144), .A0N(\ram[68][15] ), .A1N(n6542), 
        .Y(n1685) );
  OAI2BB2XL U478 ( .B0(n6974), .B1(n146), .A0N(\ram[69][0] ), .A1N(n6541), .Y(
        n1686) );
  OAI2BB2XL U479 ( .B0(n6951), .B1(n146), .A0N(\ram[69][1] ), .A1N(n6541), .Y(
        n1687) );
  OAI2BB2XL U480 ( .B0(n6928), .B1(n146), .A0N(\ram[69][2] ), .A1N(n6541), .Y(
        n1688) );
  OAI2BB2XL U481 ( .B0(n6905), .B1(n146), .A0N(\ram[69][3] ), .A1N(n6541), .Y(
        n1689) );
  OAI2BB2XL U482 ( .B0(n6877), .B1(n146), .A0N(\ram[69][4] ), .A1N(n6541), .Y(
        n1690) );
  OAI2BB2XL U483 ( .B0(n6854), .B1(n146), .A0N(\ram[69][5] ), .A1N(n6541), .Y(
        n1691) );
  OAI2BB2XL U484 ( .B0(n6831), .B1(n146), .A0N(\ram[69][6] ), .A1N(n6541), .Y(
        n1692) );
  OAI2BB2XL U485 ( .B0(n6808), .B1(n146), .A0N(\ram[69][7] ), .A1N(n6541), .Y(
        n1693) );
  OAI2BB2XL U486 ( .B0(n6785), .B1(n146), .A0N(\ram[69][8] ), .A1N(n6541), .Y(
        n1694) );
  OAI2BB2XL U487 ( .B0(n6762), .B1(n146), .A0N(\ram[69][9] ), .A1N(n6541), .Y(
        n1695) );
  OAI2BB2XL U488 ( .B0(n6739), .B1(n146), .A0N(\ram[69][10] ), .A1N(n6541), 
        .Y(n1696) );
  OAI2BB2XL U489 ( .B0(n6716), .B1(n146), .A0N(\ram[69][11] ), .A1N(n6541), 
        .Y(n1697) );
  OAI2BB2XL U490 ( .B0(n6693), .B1(n146), .A0N(\ram[69][12] ), .A1N(n6541), 
        .Y(n1698) );
  OAI2BB2XL U491 ( .B0(n6670), .B1(n146), .A0N(\ram[69][13] ), .A1N(n6541), 
        .Y(n1699) );
  OAI2BB2XL U492 ( .B0(n6647), .B1(n146), .A0N(\ram[69][14] ), .A1N(n6541), 
        .Y(n1700) );
  OAI2BB2XL U493 ( .B0(n6624), .B1(n146), .A0N(\ram[69][15] ), .A1N(n6541), 
        .Y(n1701) );
  OAI2BB2XL U494 ( .B0(n6974), .B1(n148), .A0N(\ram[70][0] ), .A1N(n6540), .Y(
        n1702) );
  OAI2BB2XL U495 ( .B0(n6951), .B1(n148), .A0N(\ram[70][1] ), .A1N(n6540), .Y(
        n1703) );
  OAI2BB2XL U496 ( .B0(n6928), .B1(n148), .A0N(\ram[70][2] ), .A1N(n6540), .Y(
        n1704) );
  OAI2BB2XL U497 ( .B0(n6905), .B1(n148), .A0N(\ram[70][3] ), .A1N(n6540), .Y(
        n1705) );
  OAI2BB2XL U498 ( .B0(n6877), .B1(n148), .A0N(\ram[70][4] ), .A1N(n6540), .Y(
        n1706) );
  OAI2BB2XL U499 ( .B0(n6854), .B1(n148), .A0N(\ram[70][5] ), .A1N(n6540), .Y(
        n1707) );
  OAI2BB2XL U500 ( .B0(n6831), .B1(n148), .A0N(\ram[70][6] ), .A1N(n6540), .Y(
        n1708) );
  OAI2BB2XL U501 ( .B0(n6808), .B1(n148), .A0N(\ram[70][7] ), .A1N(n6540), .Y(
        n1709) );
  OAI2BB2XL U502 ( .B0(n6785), .B1(n148), .A0N(\ram[70][8] ), .A1N(n6540), .Y(
        n1710) );
  OAI2BB2XL U503 ( .B0(n6762), .B1(n148), .A0N(\ram[70][9] ), .A1N(n6540), .Y(
        n1711) );
  OAI2BB2XL U504 ( .B0(n6739), .B1(n148), .A0N(\ram[70][10] ), .A1N(n6540), 
        .Y(n1712) );
  OAI2BB2XL U505 ( .B0(n6716), .B1(n148), .A0N(\ram[70][11] ), .A1N(n6540), 
        .Y(n1713) );
  OAI2BB2XL U506 ( .B0(n6693), .B1(n148), .A0N(\ram[70][12] ), .A1N(n6540), 
        .Y(n1714) );
  OAI2BB2XL U507 ( .B0(n6670), .B1(n148), .A0N(\ram[70][13] ), .A1N(n6540), 
        .Y(n1715) );
  OAI2BB2XL U508 ( .B0(n6647), .B1(n148), .A0N(\ram[70][14] ), .A1N(n6540), 
        .Y(n1716) );
  OAI2BB2XL U509 ( .B0(n6624), .B1(n148), .A0N(\ram[70][15] ), .A1N(n6540), 
        .Y(n1717) );
  OAI2BB2XL U510 ( .B0(n6974), .B1(n150), .A0N(\ram[71][0] ), .A1N(n6539), .Y(
        n1718) );
  OAI2BB2XL U511 ( .B0(n6951), .B1(n150), .A0N(\ram[71][1] ), .A1N(n6539), .Y(
        n1719) );
  OAI2BB2XL U512 ( .B0(n6928), .B1(n150), .A0N(\ram[71][2] ), .A1N(n6539), .Y(
        n1720) );
  OAI2BB2XL U513 ( .B0(n6905), .B1(n150), .A0N(\ram[71][3] ), .A1N(n6539), .Y(
        n1721) );
  OAI2BB2XL U514 ( .B0(n6877), .B1(n150), .A0N(\ram[71][4] ), .A1N(n6539), .Y(
        n1722) );
  OAI2BB2XL U515 ( .B0(n6854), .B1(n150), .A0N(\ram[71][5] ), .A1N(n6539), .Y(
        n1723) );
  OAI2BB2XL U516 ( .B0(n6831), .B1(n150), .A0N(\ram[71][6] ), .A1N(n6539), .Y(
        n1724) );
  OAI2BB2XL U517 ( .B0(n6808), .B1(n150), .A0N(\ram[71][7] ), .A1N(n6539), .Y(
        n1725) );
  OAI2BB2XL U518 ( .B0(n6785), .B1(n150), .A0N(\ram[71][8] ), .A1N(n6539), .Y(
        n1726) );
  OAI2BB2XL U519 ( .B0(n6762), .B1(n150), .A0N(\ram[71][9] ), .A1N(n6539), .Y(
        n1727) );
  OAI2BB2XL U520 ( .B0(n6739), .B1(n150), .A0N(\ram[71][10] ), .A1N(n6539), 
        .Y(n1728) );
  OAI2BB2XL U521 ( .B0(n6716), .B1(n150), .A0N(\ram[71][11] ), .A1N(n6539), 
        .Y(n1729) );
  OAI2BB2XL U522 ( .B0(n6693), .B1(n150), .A0N(\ram[71][12] ), .A1N(n6539), 
        .Y(n1730) );
  OAI2BB2XL U523 ( .B0(n6670), .B1(n150), .A0N(\ram[71][13] ), .A1N(n6539), 
        .Y(n1731) );
  OAI2BB2XL U524 ( .B0(n6647), .B1(n150), .A0N(\ram[71][14] ), .A1N(n6539), 
        .Y(n1732) );
  OAI2BB2XL U525 ( .B0(n6624), .B1(n150), .A0N(\ram[71][15] ), .A1N(n6539), 
        .Y(n1733) );
  OAI2BB2XL U526 ( .B0(n6974), .B1(n152), .A0N(\ram[72][0] ), .A1N(n6538), .Y(
        n1734) );
  OAI2BB2XL U527 ( .B0(n6951), .B1(n152), .A0N(\ram[72][1] ), .A1N(n6538), .Y(
        n1735) );
  OAI2BB2XL U528 ( .B0(n6928), .B1(n152), .A0N(\ram[72][2] ), .A1N(n6538), .Y(
        n1736) );
  OAI2BB2XL U529 ( .B0(n6905), .B1(n152), .A0N(\ram[72][3] ), .A1N(n6538), .Y(
        n1737) );
  OAI2BB2XL U530 ( .B0(n6877), .B1(n152), .A0N(\ram[72][4] ), .A1N(n6538), .Y(
        n1738) );
  OAI2BB2XL U531 ( .B0(n6854), .B1(n152), .A0N(\ram[72][5] ), .A1N(n6538), .Y(
        n1739) );
  OAI2BB2XL U532 ( .B0(n6831), .B1(n152), .A0N(\ram[72][6] ), .A1N(n6538), .Y(
        n1740) );
  OAI2BB2XL U533 ( .B0(n6808), .B1(n152), .A0N(\ram[72][7] ), .A1N(n6538), .Y(
        n1741) );
  OAI2BB2XL U534 ( .B0(n6785), .B1(n152), .A0N(\ram[72][8] ), .A1N(n6538), .Y(
        n1742) );
  OAI2BB2XL U535 ( .B0(n6762), .B1(n152), .A0N(\ram[72][9] ), .A1N(n6538), .Y(
        n1743) );
  OAI2BB2XL U536 ( .B0(n6739), .B1(n152), .A0N(\ram[72][10] ), .A1N(n6538), 
        .Y(n1744) );
  OAI2BB2XL U537 ( .B0(n6716), .B1(n152), .A0N(\ram[72][11] ), .A1N(n6538), 
        .Y(n1745) );
  OAI2BB2XL U538 ( .B0(n6693), .B1(n152), .A0N(\ram[72][12] ), .A1N(n6538), 
        .Y(n1746) );
  OAI2BB2XL U539 ( .B0(n6670), .B1(n152), .A0N(\ram[72][13] ), .A1N(n6538), 
        .Y(n1747) );
  OAI2BB2XL U540 ( .B0(n6647), .B1(n152), .A0N(\ram[72][14] ), .A1N(n6538), 
        .Y(n1748) );
  OAI2BB2XL U541 ( .B0(n6624), .B1(n152), .A0N(\ram[72][15] ), .A1N(n6538), 
        .Y(n1749) );
  OAI2BB2XL U542 ( .B0(n6974), .B1(n154), .A0N(\ram[73][0] ), .A1N(n6537), .Y(
        n1750) );
  OAI2BB2XL U543 ( .B0(n6951), .B1(n154), .A0N(\ram[73][1] ), .A1N(n6537), .Y(
        n1751) );
  OAI2BB2XL U544 ( .B0(n6928), .B1(n154), .A0N(\ram[73][2] ), .A1N(n6537), .Y(
        n1752) );
  OAI2BB2XL U545 ( .B0(n6905), .B1(n154), .A0N(\ram[73][3] ), .A1N(n6537), .Y(
        n1753) );
  OAI2BB2XL U546 ( .B0(n6877), .B1(n154), .A0N(\ram[73][4] ), .A1N(n6537), .Y(
        n1754) );
  OAI2BB2XL U547 ( .B0(n6854), .B1(n154), .A0N(\ram[73][5] ), .A1N(n6537), .Y(
        n1755) );
  OAI2BB2XL U548 ( .B0(n6831), .B1(n154), .A0N(\ram[73][6] ), .A1N(n6537), .Y(
        n1756) );
  OAI2BB2XL U549 ( .B0(n6808), .B1(n154), .A0N(\ram[73][7] ), .A1N(n6537), .Y(
        n1757) );
  OAI2BB2XL U550 ( .B0(n6785), .B1(n154), .A0N(\ram[73][8] ), .A1N(n6537), .Y(
        n1758) );
  OAI2BB2XL U551 ( .B0(n6762), .B1(n154), .A0N(\ram[73][9] ), .A1N(n6537), .Y(
        n1759) );
  OAI2BB2XL U552 ( .B0(n6739), .B1(n154), .A0N(\ram[73][10] ), .A1N(n6537), 
        .Y(n1760) );
  OAI2BB2XL U553 ( .B0(n6716), .B1(n154), .A0N(\ram[73][11] ), .A1N(n6537), 
        .Y(n1761) );
  OAI2BB2XL U554 ( .B0(n6693), .B1(n154), .A0N(\ram[73][12] ), .A1N(n6537), 
        .Y(n1762) );
  OAI2BB2XL U555 ( .B0(n6670), .B1(n154), .A0N(\ram[73][13] ), .A1N(n6537), 
        .Y(n1763) );
  OAI2BB2XL U556 ( .B0(n6647), .B1(n154), .A0N(\ram[73][14] ), .A1N(n6537), 
        .Y(n1764) );
  OAI2BB2XL U557 ( .B0(n6624), .B1(n154), .A0N(\ram[73][15] ), .A1N(n6537), 
        .Y(n1765) );
  OAI2BB2XL U558 ( .B0(n6974), .B1(n156), .A0N(\ram[74][0] ), .A1N(n6536), .Y(
        n1766) );
  OAI2BB2XL U559 ( .B0(n6951), .B1(n156), .A0N(\ram[74][1] ), .A1N(n6536), .Y(
        n1767) );
  OAI2BB2XL U560 ( .B0(n6928), .B1(n156), .A0N(\ram[74][2] ), .A1N(n6536), .Y(
        n1768) );
  OAI2BB2XL U561 ( .B0(n6905), .B1(n156), .A0N(\ram[74][3] ), .A1N(n6536), .Y(
        n1769) );
  OAI2BB2XL U562 ( .B0(n6877), .B1(n156), .A0N(\ram[74][4] ), .A1N(n6536), .Y(
        n1770) );
  OAI2BB2XL U563 ( .B0(n6854), .B1(n156), .A0N(\ram[74][5] ), .A1N(n6536), .Y(
        n1771) );
  OAI2BB2XL U564 ( .B0(n6831), .B1(n156), .A0N(\ram[74][6] ), .A1N(n6536), .Y(
        n1772) );
  OAI2BB2XL U565 ( .B0(n6808), .B1(n156), .A0N(\ram[74][7] ), .A1N(n6536), .Y(
        n1773) );
  OAI2BB2XL U566 ( .B0(n6785), .B1(n156), .A0N(\ram[74][8] ), .A1N(n6536), .Y(
        n1774) );
  OAI2BB2XL U567 ( .B0(n6762), .B1(n156), .A0N(\ram[74][9] ), .A1N(n6536), .Y(
        n1775) );
  OAI2BB2XL U568 ( .B0(n6739), .B1(n156), .A0N(\ram[74][10] ), .A1N(n6536), 
        .Y(n1776) );
  OAI2BB2XL U569 ( .B0(n6716), .B1(n156), .A0N(\ram[74][11] ), .A1N(n6536), 
        .Y(n1777) );
  OAI2BB2XL U570 ( .B0(n6693), .B1(n156), .A0N(\ram[74][12] ), .A1N(n6536), 
        .Y(n1778) );
  OAI2BB2XL U571 ( .B0(n6670), .B1(n156), .A0N(\ram[74][13] ), .A1N(n6536), 
        .Y(n1779) );
  OAI2BB2XL U572 ( .B0(n6647), .B1(n156), .A0N(\ram[74][14] ), .A1N(n6536), 
        .Y(n1780) );
  OAI2BB2XL U573 ( .B0(n6624), .B1(n156), .A0N(\ram[74][15] ), .A1N(n6536), 
        .Y(n1781) );
  OAI2BB2XL U574 ( .B0(n6974), .B1(n158), .A0N(\ram[75][0] ), .A1N(n6535), .Y(
        n1782) );
  OAI2BB2XL U575 ( .B0(n6951), .B1(n158), .A0N(\ram[75][1] ), .A1N(n6535), .Y(
        n1783) );
  OAI2BB2XL U576 ( .B0(n6928), .B1(n158), .A0N(\ram[75][2] ), .A1N(n6535), .Y(
        n1784) );
  OAI2BB2XL U577 ( .B0(n6905), .B1(n158), .A0N(\ram[75][3] ), .A1N(n6535), .Y(
        n1785) );
  OAI2BB2XL U578 ( .B0(n6877), .B1(n158), .A0N(\ram[75][4] ), .A1N(n6535), .Y(
        n1786) );
  OAI2BB2XL U579 ( .B0(n6854), .B1(n158), .A0N(\ram[75][5] ), .A1N(n6535), .Y(
        n1787) );
  OAI2BB2XL U580 ( .B0(n6831), .B1(n158), .A0N(\ram[75][6] ), .A1N(n6535), .Y(
        n1788) );
  OAI2BB2XL U581 ( .B0(n6808), .B1(n158), .A0N(\ram[75][7] ), .A1N(n6535), .Y(
        n1789) );
  OAI2BB2XL U582 ( .B0(n6785), .B1(n158), .A0N(\ram[75][8] ), .A1N(n6535), .Y(
        n1790) );
  OAI2BB2XL U583 ( .B0(n6762), .B1(n158), .A0N(\ram[75][9] ), .A1N(n6535), .Y(
        n1791) );
  OAI2BB2XL U584 ( .B0(n6739), .B1(n158), .A0N(\ram[75][10] ), .A1N(n6535), 
        .Y(n1792) );
  OAI2BB2XL U585 ( .B0(n6716), .B1(n158), .A0N(\ram[75][11] ), .A1N(n6535), 
        .Y(n1793) );
  OAI2BB2XL U586 ( .B0(n6693), .B1(n158), .A0N(\ram[75][12] ), .A1N(n6535), 
        .Y(n1794) );
  OAI2BB2XL U587 ( .B0(n6670), .B1(n158), .A0N(\ram[75][13] ), .A1N(n6535), 
        .Y(n1795) );
  OAI2BB2XL U588 ( .B0(n6647), .B1(n158), .A0N(\ram[75][14] ), .A1N(n6535), 
        .Y(n1796) );
  OAI2BB2XL U589 ( .B0(n6624), .B1(n158), .A0N(\ram[75][15] ), .A1N(n6535), 
        .Y(n1797) );
  OAI2BB2XL U590 ( .B0(n6973), .B1(n160), .A0N(\ram[76][0] ), .A1N(n6534), .Y(
        n1798) );
  OAI2BB2XL U591 ( .B0(n6950), .B1(n160), .A0N(\ram[76][1] ), .A1N(n6534), .Y(
        n1799) );
  OAI2BB2XL U592 ( .B0(n6927), .B1(n160), .A0N(\ram[76][2] ), .A1N(n6534), .Y(
        n1800) );
  OAI2BB2XL U593 ( .B0(n6904), .B1(n160), .A0N(\ram[76][3] ), .A1N(n6534), .Y(
        n1801) );
  OAI2BB2XL U594 ( .B0(n6876), .B1(n160), .A0N(\ram[76][4] ), .A1N(n6534), .Y(
        n1802) );
  OAI2BB2XL U595 ( .B0(n6853), .B1(n160), .A0N(\ram[76][5] ), .A1N(n6534), .Y(
        n1803) );
  OAI2BB2XL U596 ( .B0(n6830), .B1(n160), .A0N(\ram[76][6] ), .A1N(n6534), .Y(
        n1804) );
  OAI2BB2XL U597 ( .B0(n6807), .B1(n160), .A0N(\ram[76][7] ), .A1N(n6534), .Y(
        n1805) );
  OAI2BB2XL U598 ( .B0(n6784), .B1(n160), .A0N(\ram[76][8] ), .A1N(n6534), .Y(
        n1806) );
  OAI2BB2XL U599 ( .B0(n6761), .B1(n160), .A0N(\ram[76][9] ), .A1N(n6534), .Y(
        n1807) );
  OAI2BB2XL U600 ( .B0(n6738), .B1(n160), .A0N(\ram[76][10] ), .A1N(n6534), 
        .Y(n1808) );
  OAI2BB2XL U601 ( .B0(n6715), .B1(n160), .A0N(\ram[76][11] ), .A1N(n6534), 
        .Y(n1809) );
  OAI2BB2XL U602 ( .B0(n6692), .B1(n160), .A0N(\ram[76][12] ), .A1N(n6534), 
        .Y(n1810) );
  OAI2BB2XL U603 ( .B0(n6669), .B1(n160), .A0N(\ram[76][13] ), .A1N(n6534), 
        .Y(n1811) );
  OAI2BB2XL U604 ( .B0(n6646), .B1(n160), .A0N(\ram[76][14] ), .A1N(n6534), 
        .Y(n1812) );
  OAI2BB2XL U605 ( .B0(n6623), .B1(n160), .A0N(\ram[76][15] ), .A1N(n6534), 
        .Y(n1813) );
  OAI2BB2XL U606 ( .B0(n6973), .B1(n162), .A0N(\ram[77][0] ), .A1N(n6533), .Y(
        n1814) );
  OAI2BB2XL U607 ( .B0(n6950), .B1(n162), .A0N(\ram[77][1] ), .A1N(n6533), .Y(
        n1815) );
  OAI2BB2XL U608 ( .B0(n6927), .B1(n162), .A0N(\ram[77][2] ), .A1N(n6533), .Y(
        n1816) );
  OAI2BB2XL U609 ( .B0(n6904), .B1(n162), .A0N(\ram[77][3] ), .A1N(n6533), .Y(
        n1817) );
  OAI2BB2XL U610 ( .B0(n6876), .B1(n162), .A0N(\ram[77][4] ), .A1N(n6533), .Y(
        n1818) );
  OAI2BB2XL U611 ( .B0(n6853), .B1(n162), .A0N(\ram[77][5] ), .A1N(n6533), .Y(
        n1819) );
  OAI2BB2XL U612 ( .B0(n6830), .B1(n162), .A0N(\ram[77][6] ), .A1N(n6533), .Y(
        n1820) );
  OAI2BB2XL U613 ( .B0(n6807), .B1(n162), .A0N(\ram[77][7] ), .A1N(n6533), .Y(
        n1821) );
  OAI2BB2XL U614 ( .B0(n6784), .B1(n162), .A0N(\ram[77][8] ), .A1N(n6533), .Y(
        n1822) );
  OAI2BB2XL U615 ( .B0(n6761), .B1(n162), .A0N(\ram[77][9] ), .A1N(n6533), .Y(
        n1823) );
  OAI2BB2XL U616 ( .B0(n6738), .B1(n162), .A0N(\ram[77][10] ), .A1N(n6533), 
        .Y(n1824) );
  OAI2BB2XL U617 ( .B0(n6715), .B1(n162), .A0N(\ram[77][11] ), .A1N(n6533), 
        .Y(n1825) );
  OAI2BB2XL U618 ( .B0(n6692), .B1(n162), .A0N(\ram[77][12] ), .A1N(n6533), 
        .Y(n1826) );
  OAI2BB2XL U619 ( .B0(n6669), .B1(n162), .A0N(\ram[77][13] ), .A1N(n6533), 
        .Y(n1827) );
  OAI2BB2XL U620 ( .B0(n6646), .B1(n162), .A0N(\ram[77][14] ), .A1N(n6533), 
        .Y(n1828) );
  OAI2BB2XL U621 ( .B0(n6623), .B1(n162), .A0N(\ram[77][15] ), .A1N(n6533), 
        .Y(n1829) );
  OAI2BB2XL U622 ( .B0(n6973), .B1(n164), .A0N(\ram[78][0] ), .A1N(n6532), .Y(
        n1830) );
  OAI2BB2XL U623 ( .B0(n6950), .B1(n164), .A0N(\ram[78][1] ), .A1N(n6532), .Y(
        n1831) );
  OAI2BB2XL U624 ( .B0(n6927), .B1(n164), .A0N(\ram[78][2] ), .A1N(n6532), .Y(
        n1832) );
  OAI2BB2XL U625 ( .B0(n6904), .B1(n164), .A0N(\ram[78][3] ), .A1N(n6532), .Y(
        n1833) );
  OAI2BB2XL U626 ( .B0(n6876), .B1(n164), .A0N(\ram[78][4] ), .A1N(n6532), .Y(
        n1834) );
  OAI2BB2XL U627 ( .B0(n6853), .B1(n164), .A0N(\ram[78][5] ), .A1N(n6532), .Y(
        n1835) );
  OAI2BB2XL U628 ( .B0(n6830), .B1(n164), .A0N(\ram[78][6] ), .A1N(n6532), .Y(
        n1836) );
  OAI2BB2XL U629 ( .B0(n6807), .B1(n164), .A0N(\ram[78][7] ), .A1N(n6532), .Y(
        n1837) );
  OAI2BB2XL U630 ( .B0(n6784), .B1(n164), .A0N(\ram[78][8] ), .A1N(n6532), .Y(
        n1838) );
  OAI2BB2XL U631 ( .B0(n6761), .B1(n164), .A0N(\ram[78][9] ), .A1N(n6532), .Y(
        n1839) );
  OAI2BB2XL U632 ( .B0(n6738), .B1(n164), .A0N(\ram[78][10] ), .A1N(n6532), 
        .Y(n1840) );
  OAI2BB2XL U633 ( .B0(n6715), .B1(n164), .A0N(\ram[78][11] ), .A1N(n6532), 
        .Y(n1841) );
  OAI2BB2XL U634 ( .B0(n6692), .B1(n164), .A0N(\ram[78][12] ), .A1N(n6532), 
        .Y(n1842) );
  OAI2BB2XL U635 ( .B0(n6669), .B1(n164), .A0N(\ram[78][13] ), .A1N(n6532), 
        .Y(n1843) );
  OAI2BB2XL U636 ( .B0(n6646), .B1(n164), .A0N(\ram[78][14] ), .A1N(n6532), 
        .Y(n1844) );
  OAI2BB2XL U637 ( .B0(n6623), .B1(n164), .A0N(\ram[78][15] ), .A1N(n6532), 
        .Y(n1845) );
  OAI2BB2XL U638 ( .B0(n6973), .B1(n166), .A0N(\ram[79][0] ), .A1N(n6531), .Y(
        n1846) );
  OAI2BB2XL U639 ( .B0(n6950), .B1(n166), .A0N(\ram[79][1] ), .A1N(n6531), .Y(
        n1847) );
  OAI2BB2XL U640 ( .B0(n6927), .B1(n166), .A0N(\ram[79][2] ), .A1N(n6531), .Y(
        n1848) );
  OAI2BB2XL U641 ( .B0(n6904), .B1(n166), .A0N(\ram[79][3] ), .A1N(n6531), .Y(
        n1849) );
  OAI2BB2XL U642 ( .B0(n6876), .B1(n166), .A0N(\ram[79][4] ), .A1N(n6531), .Y(
        n1850) );
  OAI2BB2XL U643 ( .B0(n6853), .B1(n166), .A0N(\ram[79][5] ), .A1N(n6531), .Y(
        n1851) );
  OAI2BB2XL U644 ( .B0(n6830), .B1(n166), .A0N(\ram[79][6] ), .A1N(n6531), .Y(
        n1852) );
  OAI2BB2XL U645 ( .B0(n6807), .B1(n166), .A0N(\ram[79][7] ), .A1N(n6531), .Y(
        n1853) );
  OAI2BB2XL U646 ( .B0(n6784), .B1(n166), .A0N(\ram[79][8] ), .A1N(n6531), .Y(
        n1854) );
  OAI2BB2XL U647 ( .B0(n6761), .B1(n166), .A0N(\ram[79][9] ), .A1N(n6531), .Y(
        n1855) );
  OAI2BB2XL U648 ( .B0(n6738), .B1(n166), .A0N(\ram[79][10] ), .A1N(n6531), 
        .Y(n1856) );
  OAI2BB2XL U649 ( .B0(n6715), .B1(n166), .A0N(\ram[79][11] ), .A1N(n6531), 
        .Y(n1857) );
  OAI2BB2XL U650 ( .B0(n6692), .B1(n166), .A0N(\ram[79][12] ), .A1N(n6531), 
        .Y(n1858) );
  OAI2BB2XL U651 ( .B0(n6669), .B1(n166), .A0N(\ram[79][13] ), .A1N(n6531), 
        .Y(n1859) );
  OAI2BB2XL U652 ( .B0(n6646), .B1(n166), .A0N(\ram[79][14] ), .A1N(n6531), 
        .Y(n1860) );
  OAI2BB2XL U653 ( .B0(n6623), .B1(n166), .A0N(\ram[79][15] ), .A1N(n6531), 
        .Y(n1861) );
  OAI2BB2XL U654 ( .B0(n6969), .B1(n261), .A0N(\ram[128][0] ), .A1N(n6482), 
        .Y(n2630) );
  OAI2BB2XL U655 ( .B0(n6946), .B1(n261), .A0N(\ram[128][1] ), .A1N(n6482), 
        .Y(n2631) );
  OAI2BB2XL U656 ( .B0(n6923), .B1(n261), .A0N(\ram[128][2] ), .A1N(n6482), 
        .Y(n2632) );
  OAI2BB2XL U657 ( .B0(n6900), .B1(n261), .A0N(\ram[128][3] ), .A1N(n6482), 
        .Y(n2633) );
  OAI2BB2XL U658 ( .B0(n6872), .B1(n261), .A0N(\ram[128][4] ), .A1N(n6482), 
        .Y(n2634) );
  OAI2BB2XL U659 ( .B0(n6849), .B1(n261), .A0N(\ram[128][5] ), .A1N(n6482), 
        .Y(n2635) );
  OAI2BB2XL U660 ( .B0(n6826), .B1(n261), .A0N(\ram[128][6] ), .A1N(n6482), 
        .Y(n2636) );
  OAI2BB2XL U661 ( .B0(n6803), .B1(n261), .A0N(\ram[128][7] ), .A1N(n6482), 
        .Y(n2637) );
  OAI2BB2XL U662 ( .B0(n6780), .B1(n261), .A0N(\ram[128][8] ), .A1N(n6482), 
        .Y(n2638) );
  OAI2BB2XL U663 ( .B0(n6757), .B1(n261), .A0N(\ram[128][9] ), .A1N(n6482), 
        .Y(n2639) );
  OAI2BB2XL U664 ( .B0(n6734), .B1(n261), .A0N(\ram[128][10] ), .A1N(n6482), 
        .Y(n2640) );
  OAI2BB2XL U665 ( .B0(n6711), .B1(n261), .A0N(\ram[128][11] ), .A1N(n6482), 
        .Y(n2641) );
  OAI2BB2XL U666 ( .B0(n6688), .B1(n261), .A0N(\ram[128][12] ), .A1N(n6482), 
        .Y(n2642) );
  OAI2BB2XL U667 ( .B0(n6665), .B1(n261), .A0N(\ram[128][13] ), .A1N(n6482), 
        .Y(n2643) );
  OAI2BB2XL U668 ( .B0(n6642), .B1(n261), .A0N(\ram[128][14] ), .A1N(n6482), 
        .Y(n2644) );
  OAI2BB2XL U669 ( .B0(n6619), .B1(n261), .A0N(\ram[128][15] ), .A1N(n6482), 
        .Y(n2645) );
  OAI2BB2XL U670 ( .B0(n6969), .B1(n263), .A0N(\ram[129][0] ), .A1N(n6481), 
        .Y(n2646) );
  OAI2BB2XL U671 ( .B0(n6946), .B1(n263), .A0N(\ram[129][1] ), .A1N(n6481), 
        .Y(n2647) );
  OAI2BB2XL U672 ( .B0(n6923), .B1(n263), .A0N(\ram[129][2] ), .A1N(n6481), 
        .Y(n2648) );
  OAI2BB2XL U673 ( .B0(n6900), .B1(n263), .A0N(\ram[129][3] ), .A1N(n6481), 
        .Y(n2649) );
  OAI2BB2XL U674 ( .B0(n6872), .B1(n263), .A0N(\ram[129][4] ), .A1N(n6481), 
        .Y(n2650) );
  OAI2BB2XL U675 ( .B0(n6849), .B1(n263), .A0N(\ram[129][5] ), .A1N(n6481), 
        .Y(n2651) );
  OAI2BB2XL U676 ( .B0(n6826), .B1(n263), .A0N(\ram[129][6] ), .A1N(n6481), 
        .Y(n2652) );
  OAI2BB2XL U677 ( .B0(n6803), .B1(n263), .A0N(\ram[129][7] ), .A1N(n6481), 
        .Y(n2653) );
  OAI2BB2XL U678 ( .B0(n6780), .B1(n263), .A0N(\ram[129][8] ), .A1N(n6481), 
        .Y(n2654) );
  OAI2BB2XL U679 ( .B0(n6757), .B1(n263), .A0N(\ram[129][9] ), .A1N(n6481), 
        .Y(n2655) );
  OAI2BB2XL U680 ( .B0(n6734), .B1(n263), .A0N(\ram[129][10] ), .A1N(n6481), 
        .Y(n2656) );
  OAI2BB2XL U681 ( .B0(n6711), .B1(n263), .A0N(\ram[129][11] ), .A1N(n6481), 
        .Y(n2657) );
  OAI2BB2XL U682 ( .B0(n6688), .B1(n263), .A0N(\ram[129][12] ), .A1N(n6481), 
        .Y(n2658) );
  OAI2BB2XL U683 ( .B0(n6665), .B1(n263), .A0N(\ram[129][13] ), .A1N(n6481), 
        .Y(n2659) );
  OAI2BB2XL U684 ( .B0(n6642), .B1(n263), .A0N(\ram[129][14] ), .A1N(n6481), 
        .Y(n2660) );
  OAI2BB2XL U685 ( .B0(n6619), .B1(n263), .A0N(\ram[129][15] ), .A1N(n6481), 
        .Y(n2661) );
  OAI2BB2XL U686 ( .B0(n6969), .B1(n265), .A0N(\ram[130][0] ), .A1N(n6480), 
        .Y(n2662) );
  OAI2BB2XL U687 ( .B0(n6946), .B1(n265), .A0N(\ram[130][1] ), .A1N(n6480), 
        .Y(n2663) );
  OAI2BB2XL U688 ( .B0(n6923), .B1(n265), .A0N(\ram[130][2] ), .A1N(n6480), 
        .Y(n2664) );
  OAI2BB2XL U689 ( .B0(n6900), .B1(n265), .A0N(\ram[130][3] ), .A1N(n6480), 
        .Y(n2665) );
  OAI2BB2XL U690 ( .B0(n6872), .B1(n265), .A0N(\ram[130][4] ), .A1N(n6480), 
        .Y(n2666) );
  OAI2BB2XL U691 ( .B0(n6849), .B1(n265), .A0N(\ram[130][5] ), .A1N(n6480), 
        .Y(n2667) );
  OAI2BB2XL U692 ( .B0(n6826), .B1(n265), .A0N(\ram[130][6] ), .A1N(n6480), 
        .Y(n2668) );
  OAI2BB2XL U693 ( .B0(n6803), .B1(n265), .A0N(\ram[130][7] ), .A1N(n6480), 
        .Y(n2669) );
  OAI2BB2XL U694 ( .B0(n6780), .B1(n265), .A0N(\ram[130][8] ), .A1N(n6480), 
        .Y(n2670) );
  OAI2BB2XL U695 ( .B0(n6757), .B1(n265), .A0N(\ram[130][9] ), .A1N(n6480), 
        .Y(n2671) );
  OAI2BB2XL U696 ( .B0(n6734), .B1(n265), .A0N(\ram[130][10] ), .A1N(n6480), 
        .Y(n2672) );
  OAI2BB2XL U697 ( .B0(n6711), .B1(n265), .A0N(\ram[130][11] ), .A1N(n6480), 
        .Y(n2673) );
  OAI2BB2XL U698 ( .B0(n6688), .B1(n265), .A0N(\ram[130][12] ), .A1N(n6480), 
        .Y(n2674) );
  OAI2BB2XL U699 ( .B0(n6665), .B1(n265), .A0N(\ram[130][13] ), .A1N(n6480), 
        .Y(n2675) );
  OAI2BB2XL U700 ( .B0(n6642), .B1(n265), .A0N(\ram[130][14] ), .A1N(n6480), 
        .Y(n2676) );
  OAI2BB2XL U701 ( .B0(n6619), .B1(n265), .A0N(\ram[130][15] ), .A1N(n6480), 
        .Y(n2677) );
  OAI2BB2XL U702 ( .B0(n6969), .B1(n267), .A0N(\ram[131][0] ), .A1N(n6479), 
        .Y(n2678) );
  OAI2BB2XL U703 ( .B0(n6946), .B1(n267), .A0N(\ram[131][1] ), .A1N(n6479), 
        .Y(n2679) );
  OAI2BB2XL U704 ( .B0(n6923), .B1(n267), .A0N(\ram[131][2] ), .A1N(n6479), 
        .Y(n2680) );
  OAI2BB2XL U705 ( .B0(n6900), .B1(n267), .A0N(\ram[131][3] ), .A1N(n6479), 
        .Y(n2681) );
  OAI2BB2XL U706 ( .B0(n6872), .B1(n267), .A0N(\ram[131][4] ), .A1N(n6479), 
        .Y(n2682) );
  OAI2BB2XL U707 ( .B0(n6849), .B1(n267), .A0N(\ram[131][5] ), .A1N(n6479), 
        .Y(n2683) );
  OAI2BB2XL U708 ( .B0(n6826), .B1(n267), .A0N(\ram[131][6] ), .A1N(n6479), 
        .Y(n2684) );
  OAI2BB2XL U709 ( .B0(n6803), .B1(n267), .A0N(\ram[131][7] ), .A1N(n6479), 
        .Y(n2685) );
  OAI2BB2XL U710 ( .B0(n6780), .B1(n267), .A0N(\ram[131][8] ), .A1N(n6479), 
        .Y(n2686) );
  OAI2BB2XL U711 ( .B0(n6757), .B1(n267), .A0N(\ram[131][9] ), .A1N(n6479), 
        .Y(n2687) );
  OAI2BB2XL U712 ( .B0(n6734), .B1(n267), .A0N(\ram[131][10] ), .A1N(n6479), 
        .Y(n2688) );
  OAI2BB2XL U713 ( .B0(n6711), .B1(n267), .A0N(\ram[131][11] ), .A1N(n6479), 
        .Y(n2689) );
  OAI2BB2XL U714 ( .B0(n6688), .B1(n267), .A0N(\ram[131][12] ), .A1N(n6479), 
        .Y(n2690) );
  OAI2BB2XL U715 ( .B0(n6665), .B1(n267), .A0N(\ram[131][13] ), .A1N(n6479), 
        .Y(n2691) );
  OAI2BB2XL U716 ( .B0(n6642), .B1(n267), .A0N(\ram[131][14] ), .A1N(n6479), 
        .Y(n2692) );
  OAI2BB2XL U717 ( .B0(n6619), .B1(n267), .A0N(\ram[131][15] ), .A1N(n6479), 
        .Y(n2693) );
  OAI2BB2XL U718 ( .B0(n6969), .B1(n269), .A0N(\ram[132][0] ), .A1N(n6478), 
        .Y(n2694) );
  OAI2BB2XL U719 ( .B0(n6946), .B1(n269), .A0N(\ram[132][1] ), .A1N(n6478), 
        .Y(n2695) );
  OAI2BB2XL U720 ( .B0(n6923), .B1(n269), .A0N(\ram[132][2] ), .A1N(n6478), 
        .Y(n2696) );
  OAI2BB2XL U721 ( .B0(n6900), .B1(n269), .A0N(\ram[132][3] ), .A1N(n6478), 
        .Y(n2697) );
  OAI2BB2XL U722 ( .B0(n6872), .B1(n269), .A0N(\ram[132][4] ), .A1N(n6478), 
        .Y(n2698) );
  OAI2BB2XL U723 ( .B0(n6849), .B1(n269), .A0N(\ram[132][5] ), .A1N(n6478), 
        .Y(n2699) );
  OAI2BB2XL U724 ( .B0(n6826), .B1(n269), .A0N(\ram[132][6] ), .A1N(n6478), 
        .Y(n2700) );
  OAI2BB2XL U725 ( .B0(n6803), .B1(n269), .A0N(\ram[132][7] ), .A1N(n6478), 
        .Y(n2701) );
  OAI2BB2XL U726 ( .B0(n6780), .B1(n269), .A0N(\ram[132][8] ), .A1N(n6478), 
        .Y(n2702) );
  OAI2BB2XL U727 ( .B0(n6757), .B1(n269), .A0N(\ram[132][9] ), .A1N(n6478), 
        .Y(n2703) );
  OAI2BB2XL U728 ( .B0(n6734), .B1(n269), .A0N(\ram[132][10] ), .A1N(n6478), 
        .Y(n2704) );
  OAI2BB2XL U729 ( .B0(n6711), .B1(n269), .A0N(\ram[132][11] ), .A1N(n6478), 
        .Y(n2705) );
  OAI2BB2XL U730 ( .B0(n6688), .B1(n269), .A0N(\ram[132][12] ), .A1N(n6478), 
        .Y(n2706) );
  OAI2BB2XL U731 ( .B0(n6665), .B1(n269), .A0N(\ram[132][13] ), .A1N(n6478), 
        .Y(n2707) );
  OAI2BB2XL U732 ( .B0(n6642), .B1(n269), .A0N(\ram[132][14] ), .A1N(n6478), 
        .Y(n2708) );
  OAI2BB2XL U733 ( .B0(n6619), .B1(n269), .A0N(\ram[132][15] ), .A1N(n6478), 
        .Y(n2709) );
  OAI2BB2XL U734 ( .B0(n6969), .B1(n500), .A0N(\ram[133][0] ), .A1N(n6477), 
        .Y(n2710) );
  OAI2BB2XL U735 ( .B0(n6946), .B1(n500), .A0N(\ram[133][1] ), .A1N(n6477), 
        .Y(n2711) );
  OAI2BB2XL U736 ( .B0(n6923), .B1(n500), .A0N(\ram[133][2] ), .A1N(n6477), 
        .Y(n2712) );
  OAI2BB2XL U737 ( .B0(n6900), .B1(n500), .A0N(\ram[133][3] ), .A1N(n6477), 
        .Y(n2713) );
  OAI2BB2XL U738 ( .B0(n6872), .B1(n500), .A0N(\ram[133][4] ), .A1N(n6477), 
        .Y(n2714) );
  OAI2BB2XL U739 ( .B0(n6849), .B1(n500), .A0N(\ram[133][5] ), .A1N(n6477), 
        .Y(n2715) );
  OAI2BB2XL U740 ( .B0(n6826), .B1(n500), .A0N(\ram[133][6] ), .A1N(n6477), 
        .Y(n2716) );
  OAI2BB2XL U741 ( .B0(n6803), .B1(n500), .A0N(\ram[133][7] ), .A1N(n6477), 
        .Y(n2717) );
  OAI2BB2XL U742 ( .B0(n6780), .B1(n500), .A0N(\ram[133][8] ), .A1N(n6477), 
        .Y(n2718) );
  OAI2BB2XL U743 ( .B0(n6757), .B1(n500), .A0N(\ram[133][9] ), .A1N(n6477), 
        .Y(n2719) );
  OAI2BB2XL U744 ( .B0(n6734), .B1(n500), .A0N(\ram[133][10] ), .A1N(n6477), 
        .Y(n2720) );
  OAI2BB2XL U745 ( .B0(n6711), .B1(n500), .A0N(\ram[133][11] ), .A1N(n6477), 
        .Y(n2721) );
  OAI2BB2XL U746 ( .B0(n6688), .B1(n500), .A0N(\ram[133][12] ), .A1N(n6477), 
        .Y(n2722) );
  OAI2BB2XL U747 ( .B0(n6665), .B1(n500), .A0N(\ram[133][13] ), .A1N(n6477), 
        .Y(n2723) );
  OAI2BB2XL U748 ( .B0(n6642), .B1(n500), .A0N(\ram[133][14] ), .A1N(n6477), 
        .Y(n2724) );
  OAI2BB2XL U749 ( .B0(n6619), .B1(n500), .A0N(\ram[133][15] ), .A1N(n6477), 
        .Y(n2725) );
  OAI2BB2XL U750 ( .B0(n6969), .B1(n502), .A0N(\ram[134][0] ), .A1N(n6476), 
        .Y(n2726) );
  OAI2BB2XL U751 ( .B0(n6946), .B1(n502), .A0N(\ram[134][1] ), .A1N(n6476), 
        .Y(n2727) );
  OAI2BB2XL U752 ( .B0(n6923), .B1(n502), .A0N(\ram[134][2] ), .A1N(n6476), 
        .Y(n2728) );
  OAI2BB2XL U753 ( .B0(n6900), .B1(n502), .A0N(\ram[134][3] ), .A1N(n6476), 
        .Y(n2729) );
  OAI2BB2XL U754 ( .B0(n6872), .B1(n502), .A0N(\ram[134][4] ), .A1N(n6476), 
        .Y(n2730) );
  OAI2BB2XL U755 ( .B0(n6849), .B1(n502), .A0N(\ram[134][5] ), .A1N(n6476), 
        .Y(n2731) );
  OAI2BB2XL U756 ( .B0(n6826), .B1(n502), .A0N(\ram[134][6] ), .A1N(n6476), 
        .Y(n2732) );
  OAI2BB2XL U757 ( .B0(n6803), .B1(n502), .A0N(\ram[134][7] ), .A1N(n6476), 
        .Y(n2733) );
  OAI2BB2XL U758 ( .B0(n6780), .B1(n502), .A0N(\ram[134][8] ), .A1N(n6476), 
        .Y(n2734) );
  OAI2BB2XL U759 ( .B0(n6757), .B1(n502), .A0N(\ram[134][9] ), .A1N(n6476), 
        .Y(n2735) );
  OAI2BB2XL U760 ( .B0(n6734), .B1(n502), .A0N(\ram[134][10] ), .A1N(n6476), 
        .Y(n2736) );
  OAI2BB2XL U761 ( .B0(n6711), .B1(n502), .A0N(\ram[134][11] ), .A1N(n6476), 
        .Y(n2737) );
  OAI2BB2XL U762 ( .B0(n6688), .B1(n502), .A0N(\ram[134][12] ), .A1N(n6476), 
        .Y(n2738) );
  OAI2BB2XL U763 ( .B0(n6665), .B1(n502), .A0N(\ram[134][13] ), .A1N(n6476), 
        .Y(n2739) );
  OAI2BB2XL U764 ( .B0(n6642), .B1(n502), .A0N(\ram[134][14] ), .A1N(n6476), 
        .Y(n2740) );
  OAI2BB2XL U765 ( .B0(n6619), .B1(n502), .A0N(\ram[134][15] ), .A1N(n6476), 
        .Y(n2741) );
  OAI2BB2XL U766 ( .B0(n6969), .B1(n504), .A0N(\ram[135][0] ), .A1N(n6475), 
        .Y(n2742) );
  OAI2BB2XL U767 ( .B0(n6946), .B1(n504), .A0N(\ram[135][1] ), .A1N(n6475), 
        .Y(n2743) );
  OAI2BB2XL U768 ( .B0(n6923), .B1(n504), .A0N(\ram[135][2] ), .A1N(n6475), 
        .Y(n2744) );
  OAI2BB2XL U769 ( .B0(n6900), .B1(n504), .A0N(\ram[135][3] ), .A1N(n6475), 
        .Y(n2745) );
  OAI2BB2XL U770 ( .B0(n6872), .B1(n504), .A0N(\ram[135][4] ), .A1N(n6475), 
        .Y(n2746) );
  OAI2BB2XL U771 ( .B0(n6849), .B1(n504), .A0N(\ram[135][5] ), .A1N(n6475), 
        .Y(n2747) );
  OAI2BB2XL U772 ( .B0(n6826), .B1(n504), .A0N(\ram[135][6] ), .A1N(n6475), 
        .Y(n2748) );
  OAI2BB2XL U773 ( .B0(n6803), .B1(n504), .A0N(\ram[135][7] ), .A1N(n6475), 
        .Y(n2749) );
  OAI2BB2XL U774 ( .B0(n6780), .B1(n504), .A0N(\ram[135][8] ), .A1N(n6475), 
        .Y(n2750) );
  OAI2BB2XL U775 ( .B0(n6757), .B1(n504), .A0N(\ram[135][9] ), .A1N(n6475), 
        .Y(n2751) );
  OAI2BB2XL U776 ( .B0(n6734), .B1(n504), .A0N(\ram[135][10] ), .A1N(n6475), 
        .Y(n2752) );
  OAI2BB2XL U777 ( .B0(n6711), .B1(n504), .A0N(\ram[135][11] ), .A1N(n6475), 
        .Y(n2753) );
  OAI2BB2XL U778 ( .B0(n6688), .B1(n504), .A0N(\ram[135][12] ), .A1N(n6475), 
        .Y(n2754) );
  OAI2BB2XL U779 ( .B0(n6665), .B1(n504), .A0N(\ram[135][13] ), .A1N(n6475), 
        .Y(n2755) );
  OAI2BB2XL U780 ( .B0(n6642), .B1(n504), .A0N(\ram[135][14] ), .A1N(n6475), 
        .Y(n2756) );
  OAI2BB2XL U781 ( .B0(n6619), .B1(n504), .A0N(\ram[135][15] ), .A1N(n6475), 
        .Y(n2757) );
  OAI2BB2XL U782 ( .B0(n6968), .B1(n271), .A0N(\ram[136][0] ), .A1N(n6474), 
        .Y(n2758) );
  OAI2BB2XL U783 ( .B0(n6945), .B1(n271), .A0N(\ram[136][1] ), .A1N(n6474), 
        .Y(n2759) );
  OAI2BB2XL U784 ( .B0(n6922), .B1(n271), .A0N(\ram[136][2] ), .A1N(n6474), 
        .Y(n2760) );
  OAI2BB2XL U785 ( .B0(n6899), .B1(n271), .A0N(\ram[136][3] ), .A1N(n6474), 
        .Y(n2761) );
  OAI2BB2XL U786 ( .B0(n6871), .B1(n271), .A0N(\ram[136][4] ), .A1N(n6474), 
        .Y(n2762) );
  OAI2BB2XL U787 ( .B0(n6848), .B1(n271), .A0N(\ram[136][5] ), .A1N(n6474), 
        .Y(n2763) );
  OAI2BB2XL U788 ( .B0(n6825), .B1(n271), .A0N(\ram[136][6] ), .A1N(n6474), 
        .Y(n2764) );
  OAI2BB2XL U789 ( .B0(n6802), .B1(n271), .A0N(\ram[136][7] ), .A1N(n6474), 
        .Y(n2765) );
  OAI2BB2XL U790 ( .B0(n6779), .B1(n271), .A0N(\ram[136][8] ), .A1N(n6474), 
        .Y(n2766) );
  OAI2BB2XL U791 ( .B0(n6756), .B1(n271), .A0N(\ram[136][9] ), .A1N(n6474), 
        .Y(n2767) );
  OAI2BB2XL U792 ( .B0(n6733), .B1(n271), .A0N(\ram[136][10] ), .A1N(n6474), 
        .Y(n2768) );
  OAI2BB2XL U793 ( .B0(n6710), .B1(n271), .A0N(\ram[136][11] ), .A1N(n6474), 
        .Y(n2769) );
  OAI2BB2XL U794 ( .B0(n6687), .B1(n271), .A0N(\ram[136][12] ), .A1N(n6474), 
        .Y(n2770) );
  OAI2BB2XL U795 ( .B0(n6664), .B1(n271), .A0N(\ram[136][13] ), .A1N(n6474), 
        .Y(n2771) );
  OAI2BB2XL U796 ( .B0(n6641), .B1(n271), .A0N(\ram[136][14] ), .A1N(n6474), 
        .Y(n2772) );
  OAI2BB2XL U797 ( .B0(n6618), .B1(n271), .A0N(\ram[136][15] ), .A1N(n6474), 
        .Y(n2773) );
  OAI2BB2XL U798 ( .B0(n6968), .B1(n273), .A0N(\ram[137][0] ), .A1N(n6473), 
        .Y(n2774) );
  OAI2BB2XL U799 ( .B0(n6945), .B1(n273), .A0N(\ram[137][1] ), .A1N(n6473), 
        .Y(n2775) );
  OAI2BB2XL U800 ( .B0(n6922), .B1(n273), .A0N(\ram[137][2] ), .A1N(n6473), 
        .Y(n2776) );
  OAI2BB2XL U801 ( .B0(n6899), .B1(n273), .A0N(\ram[137][3] ), .A1N(n6473), 
        .Y(n2777) );
  OAI2BB2XL U802 ( .B0(n6871), .B1(n273), .A0N(\ram[137][4] ), .A1N(n6473), 
        .Y(n2778) );
  OAI2BB2XL U803 ( .B0(n6848), .B1(n273), .A0N(\ram[137][5] ), .A1N(n6473), 
        .Y(n2779) );
  OAI2BB2XL U804 ( .B0(n6825), .B1(n273), .A0N(\ram[137][6] ), .A1N(n6473), 
        .Y(n2780) );
  OAI2BB2XL U805 ( .B0(n6802), .B1(n273), .A0N(\ram[137][7] ), .A1N(n6473), 
        .Y(n2781) );
  OAI2BB2XL U806 ( .B0(n6779), .B1(n273), .A0N(\ram[137][8] ), .A1N(n6473), 
        .Y(n2782) );
  OAI2BB2XL U807 ( .B0(n6756), .B1(n273), .A0N(\ram[137][9] ), .A1N(n6473), 
        .Y(n2783) );
  OAI2BB2XL U808 ( .B0(n6733), .B1(n273), .A0N(\ram[137][10] ), .A1N(n6473), 
        .Y(n2784) );
  OAI2BB2XL U809 ( .B0(n6710), .B1(n273), .A0N(\ram[137][11] ), .A1N(n6473), 
        .Y(n2785) );
  OAI2BB2XL U810 ( .B0(n6687), .B1(n273), .A0N(\ram[137][12] ), .A1N(n6473), 
        .Y(n2786) );
  OAI2BB2XL U811 ( .B0(n6664), .B1(n273), .A0N(\ram[137][13] ), .A1N(n6473), 
        .Y(n2787) );
  OAI2BB2XL U812 ( .B0(n6641), .B1(n273), .A0N(\ram[137][14] ), .A1N(n6473), 
        .Y(n2788) );
  OAI2BB2XL U813 ( .B0(n6618), .B1(n273), .A0N(\ram[137][15] ), .A1N(n6473), 
        .Y(n2789) );
  OAI2BB2XL U814 ( .B0(n6968), .B1(n275), .A0N(\ram[138][0] ), .A1N(n6472), 
        .Y(n2790) );
  OAI2BB2XL U815 ( .B0(n6945), .B1(n275), .A0N(\ram[138][1] ), .A1N(n6472), 
        .Y(n2791) );
  OAI2BB2XL U816 ( .B0(n6922), .B1(n275), .A0N(\ram[138][2] ), .A1N(n6472), 
        .Y(n2792) );
  OAI2BB2XL U817 ( .B0(n6899), .B1(n275), .A0N(\ram[138][3] ), .A1N(n6472), 
        .Y(n2793) );
  OAI2BB2XL U818 ( .B0(n6871), .B1(n275), .A0N(\ram[138][4] ), .A1N(n6472), 
        .Y(n2794) );
  OAI2BB2XL U819 ( .B0(n6848), .B1(n275), .A0N(\ram[138][5] ), .A1N(n6472), 
        .Y(n2795) );
  OAI2BB2XL U820 ( .B0(n6825), .B1(n275), .A0N(\ram[138][6] ), .A1N(n6472), 
        .Y(n2796) );
  OAI2BB2XL U821 ( .B0(n6802), .B1(n275), .A0N(\ram[138][7] ), .A1N(n6472), 
        .Y(n2797) );
  OAI2BB2XL U822 ( .B0(n6779), .B1(n275), .A0N(\ram[138][8] ), .A1N(n6472), 
        .Y(n2798) );
  OAI2BB2XL U823 ( .B0(n6756), .B1(n275), .A0N(\ram[138][9] ), .A1N(n6472), 
        .Y(n2799) );
  OAI2BB2XL U824 ( .B0(n6733), .B1(n275), .A0N(\ram[138][10] ), .A1N(n6472), 
        .Y(n2800) );
  OAI2BB2XL U825 ( .B0(n6710), .B1(n275), .A0N(\ram[138][11] ), .A1N(n6472), 
        .Y(n2801) );
  OAI2BB2XL U826 ( .B0(n6687), .B1(n275), .A0N(\ram[138][12] ), .A1N(n6472), 
        .Y(n2802) );
  OAI2BB2XL U827 ( .B0(n6664), .B1(n275), .A0N(\ram[138][13] ), .A1N(n6472), 
        .Y(n2803) );
  OAI2BB2XL U828 ( .B0(n6641), .B1(n275), .A0N(\ram[138][14] ), .A1N(n6472), 
        .Y(n2804) );
  OAI2BB2XL U829 ( .B0(n6618), .B1(n275), .A0N(\ram[138][15] ), .A1N(n6472), 
        .Y(n2805) );
  OAI2BB2XL U830 ( .B0(n6968), .B1(n277), .A0N(\ram[139][0] ), .A1N(n6471), 
        .Y(n2806) );
  OAI2BB2XL U831 ( .B0(n6945), .B1(n277), .A0N(\ram[139][1] ), .A1N(n6471), 
        .Y(n2807) );
  OAI2BB2XL U832 ( .B0(n6922), .B1(n277), .A0N(\ram[139][2] ), .A1N(n6471), 
        .Y(n2808) );
  OAI2BB2XL U833 ( .B0(n6899), .B1(n277), .A0N(\ram[139][3] ), .A1N(n6471), 
        .Y(n2809) );
  OAI2BB2XL U834 ( .B0(n6871), .B1(n277), .A0N(\ram[139][4] ), .A1N(n6471), 
        .Y(n2810) );
  OAI2BB2XL U835 ( .B0(n6848), .B1(n277), .A0N(\ram[139][5] ), .A1N(n6471), 
        .Y(n2811) );
  OAI2BB2XL U836 ( .B0(n6825), .B1(n277), .A0N(\ram[139][6] ), .A1N(n6471), 
        .Y(n2812) );
  OAI2BB2XL U837 ( .B0(n6802), .B1(n277), .A0N(\ram[139][7] ), .A1N(n6471), 
        .Y(n2813) );
  OAI2BB2XL U838 ( .B0(n6779), .B1(n277), .A0N(\ram[139][8] ), .A1N(n6471), 
        .Y(n2814) );
  OAI2BB2XL U839 ( .B0(n6756), .B1(n277), .A0N(\ram[139][9] ), .A1N(n6471), 
        .Y(n2815) );
  OAI2BB2XL U840 ( .B0(n6733), .B1(n277), .A0N(\ram[139][10] ), .A1N(n6471), 
        .Y(n2816) );
  OAI2BB2XL U841 ( .B0(n6710), .B1(n277), .A0N(\ram[139][11] ), .A1N(n6471), 
        .Y(n2817) );
  OAI2BB2XL U842 ( .B0(n6687), .B1(n277), .A0N(\ram[139][12] ), .A1N(n6471), 
        .Y(n2818) );
  OAI2BB2XL U843 ( .B0(n6664), .B1(n277), .A0N(\ram[139][13] ), .A1N(n6471), 
        .Y(n2819) );
  OAI2BB2XL U844 ( .B0(n6641), .B1(n277), .A0N(\ram[139][14] ), .A1N(n6471), 
        .Y(n2820) );
  OAI2BB2XL U845 ( .B0(n6618), .B1(n277), .A0N(\ram[139][15] ), .A1N(n6471), 
        .Y(n2821) );
  OAI2BB2XL U846 ( .B0(n6968), .B1(n278), .A0N(\ram[140][0] ), .A1N(n6470), 
        .Y(n2822) );
  OAI2BB2XL U847 ( .B0(n6945), .B1(n278), .A0N(\ram[140][1] ), .A1N(n6470), 
        .Y(n2823) );
  OAI2BB2XL U848 ( .B0(n6922), .B1(n278), .A0N(\ram[140][2] ), .A1N(n6470), 
        .Y(n2824) );
  OAI2BB2XL U849 ( .B0(n6899), .B1(n278), .A0N(\ram[140][3] ), .A1N(n6470), 
        .Y(n2825) );
  OAI2BB2XL U850 ( .B0(n6871), .B1(n278), .A0N(\ram[140][4] ), .A1N(n6470), 
        .Y(n2826) );
  OAI2BB2XL U851 ( .B0(n6848), .B1(n278), .A0N(\ram[140][5] ), .A1N(n6470), 
        .Y(n2827) );
  OAI2BB2XL U852 ( .B0(n6825), .B1(n278), .A0N(\ram[140][6] ), .A1N(n6470), 
        .Y(n2828) );
  OAI2BB2XL U853 ( .B0(n6802), .B1(n278), .A0N(\ram[140][7] ), .A1N(n6470), 
        .Y(n2829) );
  OAI2BB2XL U854 ( .B0(n6779), .B1(n278), .A0N(\ram[140][8] ), .A1N(n6470), 
        .Y(n2830) );
  OAI2BB2XL U855 ( .B0(n6756), .B1(n278), .A0N(\ram[140][9] ), .A1N(n6470), 
        .Y(n2831) );
  OAI2BB2XL U856 ( .B0(n6733), .B1(n278), .A0N(\ram[140][10] ), .A1N(n6470), 
        .Y(n2832) );
  OAI2BB2XL U857 ( .B0(n6710), .B1(n278), .A0N(\ram[140][11] ), .A1N(n6470), 
        .Y(n2833) );
  OAI2BB2XL U858 ( .B0(n6687), .B1(n278), .A0N(\ram[140][12] ), .A1N(n6470), 
        .Y(n2834) );
  OAI2BB2XL U859 ( .B0(n6664), .B1(n278), .A0N(\ram[140][13] ), .A1N(n6470), 
        .Y(n2835) );
  OAI2BB2XL U860 ( .B0(n6641), .B1(n278), .A0N(\ram[140][14] ), .A1N(n6470), 
        .Y(n2836) );
  OAI2BB2XL U861 ( .B0(n6618), .B1(n278), .A0N(\ram[140][15] ), .A1N(n6470), 
        .Y(n2837) );
  OAI2BB2XL U862 ( .B0(n6968), .B1(n280), .A0N(\ram[141][0] ), .A1N(n6469), 
        .Y(n2838) );
  OAI2BB2XL U863 ( .B0(n6945), .B1(n280), .A0N(\ram[141][1] ), .A1N(n6469), 
        .Y(n2839) );
  OAI2BB2XL U864 ( .B0(n6922), .B1(n280), .A0N(\ram[141][2] ), .A1N(n6469), 
        .Y(n2840) );
  OAI2BB2XL U865 ( .B0(n6899), .B1(n280), .A0N(\ram[141][3] ), .A1N(n6469), 
        .Y(n2841) );
  OAI2BB2XL U866 ( .B0(n6871), .B1(n280), .A0N(\ram[141][4] ), .A1N(n6469), 
        .Y(n2842) );
  OAI2BB2XL U867 ( .B0(n6848), .B1(n280), .A0N(\ram[141][5] ), .A1N(n6469), 
        .Y(n2843) );
  OAI2BB2XL U868 ( .B0(n6825), .B1(n280), .A0N(\ram[141][6] ), .A1N(n6469), 
        .Y(n2844) );
  OAI2BB2XL U869 ( .B0(n6802), .B1(n280), .A0N(\ram[141][7] ), .A1N(n6469), 
        .Y(n2845) );
  OAI2BB2XL U870 ( .B0(n6779), .B1(n280), .A0N(\ram[141][8] ), .A1N(n6469), 
        .Y(n2846) );
  OAI2BB2XL U871 ( .B0(n6756), .B1(n280), .A0N(\ram[141][9] ), .A1N(n6469), 
        .Y(n2847) );
  OAI2BB2XL U872 ( .B0(n6733), .B1(n280), .A0N(\ram[141][10] ), .A1N(n6469), 
        .Y(n2848) );
  OAI2BB2XL U873 ( .B0(n6710), .B1(n280), .A0N(\ram[141][11] ), .A1N(n6469), 
        .Y(n2849) );
  OAI2BB2XL U874 ( .B0(n6687), .B1(n280), .A0N(\ram[141][12] ), .A1N(n6469), 
        .Y(n2850) );
  OAI2BB2XL U875 ( .B0(n6664), .B1(n280), .A0N(\ram[141][13] ), .A1N(n6469), 
        .Y(n2851) );
  OAI2BB2XL U876 ( .B0(n6641), .B1(n280), .A0N(\ram[141][14] ), .A1N(n6469), 
        .Y(n2852) );
  OAI2BB2XL U877 ( .B0(n6618), .B1(n280), .A0N(\ram[141][15] ), .A1N(n6469), 
        .Y(n2853) );
  OAI2BB2XL U878 ( .B0(n6968), .B1(n282), .A0N(\ram[142][0] ), .A1N(n6468), 
        .Y(n2854) );
  OAI2BB2XL U879 ( .B0(n6945), .B1(n282), .A0N(\ram[142][1] ), .A1N(n6468), 
        .Y(n2855) );
  OAI2BB2XL U880 ( .B0(n6922), .B1(n282), .A0N(\ram[142][2] ), .A1N(n6468), 
        .Y(n2856) );
  OAI2BB2XL U881 ( .B0(n6899), .B1(n282), .A0N(\ram[142][3] ), .A1N(n6468), 
        .Y(n2857) );
  OAI2BB2XL U882 ( .B0(n6871), .B1(n282), .A0N(\ram[142][4] ), .A1N(n6468), 
        .Y(n2858) );
  OAI2BB2XL U883 ( .B0(n6848), .B1(n282), .A0N(\ram[142][5] ), .A1N(n6468), 
        .Y(n2859) );
  OAI2BB2XL U884 ( .B0(n6825), .B1(n282), .A0N(\ram[142][6] ), .A1N(n6468), 
        .Y(n2860) );
  OAI2BB2XL U885 ( .B0(n6802), .B1(n282), .A0N(\ram[142][7] ), .A1N(n6468), 
        .Y(n2861) );
  OAI2BB2XL U886 ( .B0(n6779), .B1(n282), .A0N(\ram[142][8] ), .A1N(n6468), 
        .Y(n2862) );
  OAI2BB2XL U887 ( .B0(n6756), .B1(n282), .A0N(\ram[142][9] ), .A1N(n6468), 
        .Y(n2863) );
  OAI2BB2XL U888 ( .B0(n6733), .B1(n282), .A0N(\ram[142][10] ), .A1N(n6468), 
        .Y(n2864) );
  OAI2BB2XL U889 ( .B0(n6710), .B1(n282), .A0N(\ram[142][11] ), .A1N(n6468), 
        .Y(n2865) );
  OAI2BB2XL U890 ( .B0(n6687), .B1(n282), .A0N(\ram[142][12] ), .A1N(n6468), 
        .Y(n2866) );
  OAI2BB2XL U891 ( .B0(n6664), .B1(n282), .A0N(\ram[142][13] ), .A1N(n6468), 
        .Y(n2867) );
  OAI2BB2XL U892 ( .B0(n6641), .B1(n282), .A0N(\ram[142][14] ), .A1N(n6468), 
        .Y(n2868) );
  OAI2BB2XL U893 ( .B0(n6618), .B1(n282), .A0N(\ram[142][15] ), .A1N(n6468), 
        .Y(n2869) );
  OAI2BB2XL U894 ( .B0(n6968), .B1(n284), .A0N(\ram[143][0] ), .A1N(n6467), 
        .Y(n2870) );
  OAI2BB2XL U895 ( .B0(n6945), .B1(n284), .A0N(\ram[143][1] ), .A1N(n6467), 
        .Y(n2871) );
  OAI2BB2XL U896 ( .B0(n6922), .B1(n284), .A0N(\ram[143][2] ), .A1N(n6467), 
        .Y(n2872) );
  OAI2BB2XL U897 ( .B0(n6899), .B1(n284), .A0N(\ram[143][3] ), .A1N(n6467), 
        .Y(n2873) );
  OAI2BB2XL U898 ( .B0(n6871), .B1(n284), .A0N(\ram[143][4] ), .A1N(n6467), 
        .Y(n2874) );
  OAI2BB2XL U899 ( .B0(n6848), .B1(n284), .A0N(\ram[143][5] ), .A1N(n6467), 
        .Y(n2875) );
  OAI2BB2XL U900 ( .B0(n6825), .B1(n284), .A0N(\ram[143][6] ), .A1N(n6467), 
        .Y(n2876) );
  OAI2BB2XL U901 ( .B0(n6802), .B1(n284), .A0N(\ram[143][7] ), .A1N(n6467), 
        .Y(n2877) );
  OAI2BB2XL U902 ( .B0(n6779), .B1(n284), .A0N(\ram[143][8] ), .A1N(n6467), 
        .Y(n2878) );
  OAI2BB2XL U903 ( .B0(n6756), .B1(n284), .A0N(\ram[143][9] ), .A1N(n6467), 
        .Y(n2879) );
  OAI2BB2XL U904 ( .B0(n6733), .B1(n284), .A0N(\ram[143][10] ), .A1N(n6467), 
        .Y(n2880) );
  OAI2BB2XL U905 ( .B0(n6710), .B1(n284), .A0N(\ram[143][11] ), .A1N(n6467), 
        .Y(n2881) );
  OAI2BB2XL U906 ( .B0(n6687), .B1(n284), .A0N(\ram[143][12] ), .A1N(n6467), 
        .Y(n2882) );
  OAI2BB2XL U907 ( .B0(n6664), .B1(n284), .A0N(\ram[143][13] ), .A1N(n6467), 
        .Y(n2883) );
  OAI2BB2XL U908 ( .B0(n6641), .B1(n284), .A0N(\ram[143][14] ), .A1N(n6467), 
        .Y(n2884) );
  OAI2BB2XL U909 ( .B0(n6618), .B1(n284), .A0N(\ram[143][15] ), .A1N(n6467), 
        .Y(n2885) );
  OAI2BB2XL U910 ( .B0(n6964), .B1(n361), .A0N(\ram[192][0] ), .A1N(n6418), 
        .Y(n3654) );
  OAI2BB2XL U911 ( .B0(n6941), .B1(n361), .A0N(\ram[192][1] ), .A1N(n6418), 
        .Y(n3655) );
  OAI2BB2XL U912 ( .B0(n6918), .B1(n361), .A0N(\ram[192][2] ), .A1N(n6418), 
        .Y(n3656) );
  OAI2BB2XL U913 ( .B0(n6895), .B1(n361), .A0N(\ram[192][3] ), .A1N(n6418), 
        .Y(n3657) );
  OAI2BB2XL U914 ( .B0(n6868), .B1(n361), .A0N(\ram[192][4] ), .A1N(n6418), 
        .Y(n3658) );
  OAI2BB2XL U915 ( .B0(n6845), .B1(n361), .A0N(\ram[192][5] ), .A1N(n6418), 
        .Y(n3659) );
  OAI2BB2XL U916 ( .B0(n6822), .B1(n361), .A0N(\ram[192][6] ), .A1N(n6418), 
        .Y(n3660) );
  OAI2BB2XL U917 ( .B0(n6799), .B1(n361), .A0N(\ram[192][7] ), .A1N(n6418), 
        .Y(n3661) );
  OAI2BB2XL U918 ( .B0(n6776), .B1(n361), .A0N(\ram[192][8] ), .A1N(n6418), 
        .Y(n3662) );
  OAI2BB2XL U919 ( .B0(n6753), .B1(n361), .A0N(\ram[192][9] ), .A1N(n6418), 
        .Y(n3663) );
  OAI2BB2XL U920 ( .B0(n6730), .B1(n361), .A0N(\ram[192][10] ), .A1N(n6418), 
        .Y(n3664) );
  OAI2BB2XL U921 ( .B0(n6707), .B1(n361), .A0N(\ram[192][11] ), .A1N(n6418), 
        .Y(n3665) );
  OAI2BB2XL U922 ( .B0(n6684), .B1(n361), .A0N(\ram[192][12] ), .A1N(n6418), 
        .Y(n3666) );
  OAI2BB2XL U923 ( .B0(n6661), .B1(n361), .A0N(\ram[192][13] ), .A1N(n6418), 
        .Y(n3667) );
  OAI2BB2XL U924 ( .B0(n6638), .B1(n361), .A0N(\ram[192][14] ), .A1N(n6418), 
        .Y(n3668) );
  OAI2BB2XL U925 ( .B0(n6615), .B1(n361), .A0N(\ram[192][15] ), .A1N(n6418), 
        .Y(n3669) );
  OAI2BB2XL U926 ( .B0(n6964), .B1(n363), .A0N(\ram[193][0] ), .A1N(n6417), 
        .Y(n3670) );
  OAI2BB2XL U927 ( .B0(n6941), .B1(n363), .A0N(\ram[193][1] ), .A1N(n6417), 
        .Y(n3671) );
  OAI2BB2XL U928 ( .B0(n6918), .B1(n363), .A0N(\ram[193][2] ), .A1N(n6417), 
        .Y(n3672) );
  OAI2BB2XL U929 ( .B0(n6895), .B1(n363), .A0N(\ram[193][3] ), .A1N(n6417), 
        .Y(n3673) );
  OAI2BB2XL U930 ( .B0(n6868), .B1(n363), .A0N(\ram[193][4] ), .A1N(n6417), 
        .Y(n3674) );
  OAI2BB2XL U931 ( .B0(n6845), .B1(n363), .A0N(\ram[193][5] ), .A1N(n6417), 
        .Y(n3675) );
  OAI2BB2XL U932 ( .B0(n6822), .B1(n363), .A0N(\ram[193][6] ), .A1N(n6417), 
        .Y(n3676) );
  OAI2BB2XL U933 ( .B0(n6799), .B1(n363), .A0N(\ram[193][7] ), .A1N(n6417), 
        .Y(n3677) );
  OAI2BB2XL U934 ( .B0(n6776), .B1(n363), .A0N(\ram[193][8] ), .A1N(n6417), 
        .Y(n3678) );
  OAI2BB2XL U935 ( .B0(n6753), .B1(n363), .A0N(\ram[193][9] ), .A1N(n6417), 
        .Y(n3679) );
  OAI2BB2XL U936 ( .B0(n6730), .B1(n363), .A0N(\ram[193][10] ), .A1N(n6417), 
        .Y(n3680) );
  OAI2BB2XL U937 ( .B0(n6707), .B1(n363), .A0N(\ram[193][11] ), .A1N(n6417), 
        .Y(n3681) );
  OAI2BB2XL U938 ( .B0(n6684), .B1(n363), .A0N(\ram[193][12] ), .A1N(n6417), 
        .Y(n3682) );
  OAI2BB2XL U939 ( .B0(n6661), .B1(n363), .A0N(\ram[193][13] ), .A1N(n6417), 
        .Y(n3683) );
  OAI2BB2XL U940 ( .B0(n6638), .B1(n363), .A0N(\ram[193][14] ), .A1N(n6417), 
        .Y(n3684) );
  OAI2BB2XL U941 ( .B0(n6615), .B1(n363), .A0N(\ram[193][15] ), .A1N(n6417), 
        .Y(n3685) );
  OAI2BB2XL U942 ( .B0(n6964), .B1(n365), .A0N(\ram[194][0] ), .A1N(n6416), 
        .Y(n3686) );
  OAI2BB2XL U943 ( .B0(n6941), .B1(n365), .A0N(\ram[194][1] ), .A1N(n6416), 
        .Y(n3687) );
  OAI2BB2XL U944 ( .B0(n6918), .B1(n365), .A0N(\ram[194][2] ), .A1N(n6416), 
        .Y(n3688) );
  OAI2BB2XL U945 ( .B0(n6895), .B1(n365), .A0N(\ram[194][3] ), .A1N(n6416), 
        .Y(n3689) );
  OAI2BB2XL U946 ( .B0(n6868), .B1(n365), .A0N(\ram[194][4] ), .A1N(n6416), 
        .Y(n3690) );
  OAI2BB2XL U947 ( .B0(n6845), .B1(n365), .A0N(\ram[194][5] ), .A1N(n6416), 
        .Y(n3691) );
  OAI2BB2XL U948 ( .B0(n6822), .B1(n365), .A0N(\ram[194][6] ), .A1N(n6416), 
        .Y(n3692) );
  OAI2BB2XL U949 ( .B0(n6799), .B1(n365), .A0N(\ram[194][7] ), .A1N(n6416), 
        .Y(n3693) );
  OAI2BB2XL U950 ( .B0(n6776), .B1(n365), .A0N(\ram[194][8] ), .A1N(n6416), 
        .Y(n3694) );
  OAI2BB2XL U951 ( .B0(n6753), .B1(n365), .A0N(\ram[194][9] ), .A1N(n6416), 
        .Y(n3695) );
  OAI2BB2XL U952 ( .B0(n6730), .B1(n365), .A0N(\ram[194][10] ), .A1N(n6416), 
        .Y(n3696) );
  OAI2BB2XL U953 ( .B0(n6707), .B1(n365), .A0N(\ram[194][11] ), .A1N(n6416), 
        .Y(n3697) );
  OAI2BB2XL U954 ( .B0(n6684), .B1(n365), .A0N(\ram[194][12] ), .A1N(n6416), 
        .Y(n3698) );
  OAI2BB2XL U955 ( .B0(n6661), .B1(n365), .A0N(\ram[194][13] ), .A1N(n6416), 
        .Y(n3699) );
  OAI2BB2XL U956 ( .B0(n6638), .B1(n365), .A0N(\ram[194][14] ), .A1N(n6416), 
        .Y(n3700) );
  OAI2BB2XL U957 ( .B0(n6615), .B1(n365), .A0N(\ram[194][15] ), .A1N(n6416), 
        .Y(n3701) );
  OAI2BB2XL U958 ( .B0(n6964), .B1(n367), .A0N(\ram[195][0] ), .A1N(n6415), 
        .Y(n3702) );
  OAI2BB2XL U959 ( .B0(n6941), .B1(n367), .A0N(\ram[195][1] ), .A1N(n6415), 
        .Y(n3703) );
  OAI2BB2XL U960 ( .B0(n6918), .B1(n367), .A0N(\ram[195][2] ), .A1N(n6415), 
        .Y(n3704) );
  OAI2BB2XL U961 ( .B0(n6895), .B1(n367), .A0N(\ram[195][3] ), .A1N(n6415), 
        .Y(n3705) );
  OAI2BB2XL U962 ( .B0(n6868), .B1(n367), .A0N(\ram[195][4] ), .A1N(n6415), 
        .Y(n3706) );
  OAI2BB2XL U963 ( .B0(n6845), .B1(n367), .A0N(\ram[195][5] ), .A1N(n6415), 
        .Y(n3707) );
  OAI2BB2XL U964 ( .B0(n6822), .B1(n367), .A0N(\ram[195][6] ), .A1N(n6415), 
        .Y(n3708) );
  OAI2BB2XL U965 ( .B0(n6799), .B1(n367), .A0N(\ram[195][7] ), .A1N(n6415), 
        .Y(n3709) );
  OAI2BB2XL U966 ( .B0(n6776), .B1(n367), .A0N(\ram[195][8] ), .A1N(n6415), 
        .Y(n3710) );
  OAI2BB2XL U967 ( .B0(n6753), .B1(n367), .A0N(\ram[195][9] ), .A1N(n6415), 
        .Y(n3711) );
  OAI2BB2XL U968 ( .B0(n6730), .B1(n367), .A0N(\ram[195][10] ), .A1N(n6415), 
        .Y(n3712) );
  OAI2BB2XL U969 ( .B0(n6707), .B1(n367), .A0N(\ram[195][11] ), .A1N(n6415), 
        .Y(n3713) );
  OAI2BB2XL U970 ( .B0(n6684), .B1(n367), .A0N(\ram[195][12] ), .A1N(n6415), 
        .Y(n3714) );
  OAI2BB2XL U971 ( .B0(n6661), .B1(n367), .A0N(\ram[195][13] ), .A1N(n6415), 
        .Y(n3715) );
  OAI2BB2XL U972 ( .B0(n6638), .B1(n367), .A0N(\ram[195][14] ), .A1N(n6415), 
        .Y(n3716) );
  OAI2BB2XL U973 ( .B0(n6615), .B1(n367), .A0N(\ram[195][15] ), .A1N(n6415), 
        .Y(n3717) );
  OAI2BB2XL U974 ( .B0(n6963), .B1(n369), .A0N(\ram[196][0] ), .A1N(n6414), 
        .Y(n3718) );
  OAI2BB2XL U975 ( .B0(n6940), .B1(n369), .A0N(\ram[196][1] ), .A1N(n6414), 
        .Y(n3719) );
  OAI2BB2XL U976 ( .B0(n6917), .B1(n369), .A0N(\ram[196][2] ), .A1N(n6414), 
        .Y(n3720) );
  OAI2BB2XL U977 ( .B0(n6894), .B1(n369), .A0N(\ram[196][3] ), .A1N(n6414), 
        .Y(n3721) );
  OAI2BB2XL U978 ( .B0(n6867), .B1(n369), .A0N(\ram[196][4] ), .A1N(n6414), 
        .Y(n3722) );
  OAI2BB2XL U979 ( .B0(n6844), .B1(n369), .A0N(\ram[196][5] ), .A1N(n6414), 
        .Y(n3723) );
  OAI2BB2XL U980 ( .B0(n6821), .B1(n369), .A0N(\ram[196][6] ), .A1N(n6414), 
        .Y(n3724) );
  OAI2BB2XL U981 ( .B0(n6798), .B1(n369), .A0N(\ram[196][7] ), .A1N(n6414), 
        .Y(n3725) );
  OAI2BB2XL U982 ( .B0(n6775), .B1(n369), .A0N(\ram[196][8] ), .A1N(n6414), 
        .Y(n3726) );
  OAI2BB2XL U983 ( .B0(n6752), .B1(n369), .A0N(\ram[196][9] ), .A1N(n6414), 
        .Y(n3727) );
  OAI2BB2XL U984 ( .B0(n6729), .B1(n369), .A0N(\ram[196][10] ), .A1N(n6414), 
        .Y(n3728) );
  OAI2BB2XL U985 ( .B0(n6706), .B1(n369), .A0N(\ram[196][11] ), .A1N(n6414), 
        .Y(n3729) );
  OAI2BB2XL U986 ( .B0(n6683), .B1(n369), .A0N(\ram[196][12] ), .A1N(n6414), 
        .Y(n3730) );
  OAI2BB2XL U987 ( .B0(n6660), .B1(n369), .A0N(\ram[196][13] ), .A1N(n6414), 
        .Y(n3731) );
  OAI2BB2XL U988 ( .B0(n6637), .B1(n369), .A0N(\ram[196][14] ), .A1N(n6414), 
        .Y(n3732) );
  OAI2BB2XL U989 ( .B0(n6614), .B1(n369), .A0N(\ram[196][15] ), .A1N(n6414), 
        .Y(n3733) );
  OAI2BB2XL U990 ( .B0(n6963), .B1(n371), .A0N(\ram[197][0] ), .A1N(n6413), 
        .Y(n3734) );
  OAI2BB2XL U991 ( .B0(n6940), .B1(n371), .A0N(\ram[197][1] ), .A1N(n6413), 
        .Y(n3735) );
  OAI2BB2XL U992 ( .B0(n6917), .B1(n371), .A0N(\ram[197][2] ), .A1N(n6413), 
        .Y(n3736) );
  OAI2BB2XL U993 ( .B0(n6894), .B1(n371), .A0N(\ram[197][3] ), .A1N(n6413), 
        .Y(n3737) );
  OAI2BB2XL U994 ( .B0(n6867), .B1(n371), .A0N(\ram[197][4] ), .A1N(n6413), 
        .Y(n3738) );
  OAI2BB2XL U995 ( .B0(n6844), .B1(n371), .A0N(\ram[197][5] ), .A1N(n6413), 
        .Y(n3739) );
  OAI2BB2XL U996 ( .B0(n6821), .B1(n371), .A0N(\ram[197][6] ), .A1N(n6413), 
        .Y(n3740) );
  OAI2BB2XL U997 ( .B0(n6798), .B1(n371), .A0N(\ram[197][7] ), .A1N(n6413), 
        .Y(n3741) );
  OAI2BB2XL U998 ( .B0(n6775), .B1(n371), .A0N(\ram[197][8] ), .A1N(n6413), 
        .Y(n3742) );
  OAI2BB2XL U999 ( .B0(n6752), .B1(n371), .A0N(\ram[197][9] ), .A1N(n6413), 
        .Y(n3743) );
  OAI2BB2XL U1000 ( .B0(n6729), .B1(n371), .A0N(\ram[197][10] ), .A1N(n6413), 
        .Y(n3744) );
  OAI2BB2XL U1001 ( .B0(n6706), .B1(n371), .A0N(\ram[197][11] ), .A1N(n6413), 
        .Y(n3745) );
  OAI2BB2XL U1002 ( .B0(n6683), .B1(n371), .A0N(\ram[197][12] ), .A1N(n6413), 
        .Y(n3746) );
  OAI2BB2XL U1003 ( .B0(n6660), .B1(n371), .A0N(\ram[197][13] ), .A1N(n6413), 
        .Y(n3747) );
  OAI2BB2XL U1004 ( .B0(n6637), .B1(n371), .A0N(\ram[197][14] ), .A1N(n6413), 
        .Y(n3748) );
  OAI2BB2XL U1005 ( .B0(n6614), .B1(n371), .A0N(\ram[197][15] ), .A1N(n6413), 
        .Y(n3749) );
  OAI2BB2XL U1006 ( .B0(n6963), .B1(n373), .A0N(\ram[198][0] ), .A1N(n6412), 
        .Y(n3750) );
  OAI2BB2XL U1007 ( .B0(n6940), .B1(n373), .A0N(\ram[198][1] ), .A1N(n6412), 
        .Y(n3751) );
  OAI2BB2XL U1008 ( .B0(n6917), .B1(n373), .A0N(\ram[198][2] ), .A1N(n6412), 
        .Y(n3752) );
  OAI2BB2XL U1009 ( .B0(n6894), .B1(n373), .A0N(\ram[198][3] ), .A1N(n6412), 
        .Y(n3753) );
  OAI2BB2XL U1010 ( .B0(n6867), .B1(n373), .A0N(\ram[198][4] ), .A1N(n6412), 
        .Y(n3754) );
  OAI2BB2XL U1011 ( .B0(n6844), .B1(n373), .A0N(\ram[198][5] ), .A1N(n6412), 
        .Y(n3755) );
  OAI2BB2XL U1012 ( .B0(n6821), .B1(n373), .A0N(\ram[198][6] ), .A1N(n6412), 
        .Y(n3756) );
  OAI2BB2XL U1013 ( .B0(n6798), .B1(n373), .A0N(\ram[198][7] ), .A1N(n6412), 
        .Y(n3757) );
  OAI2BB2XL U1014 ( .B0(n6775), .B1(n373), .A0N(\ram[198][8] ), .A1N(n6412), 
        .Y(n3758) );
  OAI2BB2XL U1015 ( .B0(n6752), .B1(n373), .A0N(\ram[198][9] ), .A1N(n6412), 
        .Y(n3759) );
  OAI2BB2XL U1016 ( .B0(n6729), .B1(n373), .A0N(\ram[198][10] ), .A1N(n6412), 
        .Y(n3760) );
  OAI2BB2XL U1017 ( .B0(n6706), .B1(n373), .A0N(\ram[198][11] ), .A1N(n6412), 
        .Y(n3761) );
  OAI2BB2XL U1018 ( .B0(n6683), .B1(n373), .A0N(\ram[198][12] ), .A1N(n6412), 
        .Y(n3762) );
  OAI2BB2XL U1019 ( .B0(n6660), .B1(n373), .A0N(\ram[198][13] ), .A1N(n6412), 
        .Y(n3763) );
  OAI2BB2XL U1020 ( .B0(n6637), .B1(n373), .A0N(\ram[198][14] ), .A1N(n6412), 
        .Y(n3764) );
  OAI2BB2XL U1021 ( .B0(n6614), .B1(n373), .A0N(\ram[198][15] ), .A1N(n6412), 
        .Y(n3765) );
  OAI2BB2XL U1022 ( .B0(n6963), .B1(n375), .A0N(\ram[199][0] ), .A1N(n6411), 
        .Y(n3766) );
  OAI2BB2XL U1023 ( .B0(n6940), .B1(n375), .A0N(\ram[199][1] ), .A1N(n6411), 
        .Y(n3767) );
  OAI2BB2XL U1024 ( .B0(n6917), .B1(n375), .A0N(\ram[199][2] ), .A1N(n6411), 
        .Y(n3768) );
  OAI2BB2XL U1025 ( .B0(n6894), .B1(n375), .A0N(\ram[199][3] ), .A1N(n6411), 
        .Y(n3769) );
  OAI2BB2XL U1026 ( .B0(n6867), .B1(n375), .A0N(\ram[199][4] ), .A1N(n6411), 
        .Y(n3770) );
  OAI2BB2XL U1027 ( .B0(n6844), .B1(n375), .A0N(\ram[199][5] ), .A1N(n6411), 
        .Y(n3771) );
  OAI2BB2XL U1028 ( .B0(n6821), .B1(n375), .A0N(\ram[199][6] ), .A1N(n6411), 
        .Y(n3772) );
  OAI2BB2XL U1029 ( .B0(n6798), .B1(n375), .A0N(\ram[199][7] ), .A1N(n6411), 
        .Y(n3773) );
  OAI2BB2XL U1030 ( .B0(n6775), .B1(n375), .A0N(\ram[199][8] ), .A1N(n6411), 
        .Y(n3774) );
  OAI2BB2XL U1031 ( .B0(n6752), .B1(n375), .A0N(\ram[199][9] ), .A1N(n6411), 
        .Y(n3775) );
  OAI2BB2XL U1032 ( .B0(n6729), .B1(n375), .A0N(\ram[199][10] ), .A1N(n6411), 
        .Y(n3776) );
  OAI2BB2XL U1033 ( .B0(n6706), .B1(n375), .A0N(\ram[199][11] ), .A1N(n6411), 
        .Y(n3777) );
  OAI2BB2XL U1034 ( .B0(n6683), .B1(n375), .A0N(\ram[199][12] ), .A1N(n6411), 
        .Y(n3778) );
  OAI2BB2XL U1035 ( .B0(n6660), .B1(n375), .A0N(\ram[199][13] ), .A1N(n6411), 
        .Y(n3779) );
  OAI2BB2XL U1036 ( .B0(n6637), .B1(n375), .A0N(\ram[199][14] ), .A1N(n6411), 
        .Y(n3780) );
  OAI2BB2XL U1037 ( .B0(n6614), .B1(n375), .A0N(\ram[199][15] ), .A1N(n6411), 
        .Y(n3781) );
  OAI2BB2XL U1038 ( .B0(n6963), .B1(n377), .A0N(\ram[200][0] ), .A1N(n6410), 
        .Y(n3782) );
  OAI2BB2XL U1039 ( .B0(n6940), .B1(n377), .A0N(\ram[200][1] ), .A1N(n6410), 
        .Y(n3783) );
  OAI2BB2XL U1040 ( .B0(n6917), .B1(n377), .A0N(\ram[200][2] ), .A1N(n6410), 
        .Y(n3784) );
  OAI2BB2XL U1041 ( .B0(n6894), .B1(n377), .A0N(\ram[200][3] ), .A1N(n6410), 
        .Y(n3785) );
  OAI2BB2XL U1042 ( .B0(n6867), .B1(n377), .A0N(\ram[200][4] ), .A1N(n6410), 
        .Y(n3786) );
  OAI2BB2XL U1043 ( .B0(n6844), .B1(n377), .A0N(\ram[200][5] ), .A1N(n6410), 
        .Y(n3787) );
  OAI2BB2XL U1044 ( .B0(n6821), .B1(n377), .A0N(\ram[200][6] ), .A1N(n6410), 
        .Y(n3788) );
  OAI2BB2XL U1045 ( .B0(n6798), .B1(n377), .A0N(\ram[200][7] ), .A1N(n6410), 
        .Y(n3789) );
  OAI2BB2XL U1046 ( .B0(n6775), .B1(n377), .A0N(\ram[200][8] ), .A1N(n6410), 
        .Y(n3790) );
  OAI2BB2XL U1047 ( .B0(n6752), .B1(n377), .A0N(\ram[200][9] ), .A1N(n6410), 
        .Y(n3791) );
  OAI2BB2XL U1048 ( .B0(n6729), .B1(n377), .A0N(\ram[200][10] ), .A1N(n6410), 
        .Y(n3792) );
  OAI2BB2XL U1049 ( .B0(n6706), .B1(n377), .A0N(\ram[200][11] ), .A1N(n6410), 
        .Y(n3793) );
  OAI2BB2XL U1050 ( .B0(n6683), .B1(n377), .A0N(\ram[200][12] ), .A1N(n6410), 
        .Y(n3794) );
  OAI2BB2XL U1051 ( .B0(n6660), .B1(n377), .A0N(\ram[200][13] ), .A1N(n6410), 
        .Y(n3795) );
  OAI2BB2XL U1052 ( .B0(n6637), .B1(n377), .A0N(\ram[200][14] ), .A1N(n6410), 
        .Y(n3796) );
  OAI2BB2XL U1053 ( .B0(n6614), .B1(n377), .A0N(\ram[200][15] ), .A1N(n6410), 
        .Y(n3797) );
  OAI2BB2XL U1054 ( .B0(n6963), .B1(n378), .A0N(\ram[201][0] ), .A1N(n6409), 
        .Y(n3798) );
  OAI2BB2XL U1055 ( .B0(n6940), .B1(n378), .A0N(\ram[201][1] ), .A1N(n6409), 
        .Y(n3799) );
  OAI2BB2XL U1056 ( .B0(n6917), .B1(n378), .A0N(\ram[201][2] ), .A1N(n6409), 
        .Y(n3800) );
  OAI2BB2XL U1057 ( .B0(n6894), .B1(n378), .A0N(\ram[201][3] ), .A1N(n6409), 
        .Y(n3801) );
  OAI2BB2XL U1058 ( .B0(n6867), .B1(n378), .A0N(\ram[201][4] ), .A1N(n6409), 
        .Y(n3802) );
  OAI2BB2XL U1059 ( .B0(n6844), .B1(n378), .A0N(\ram[201][5] ), .A1N(n6409), 
        .Y(n3803) );
  OAI2BB2XL U1060 ( .B0(n6821), .B1(n378), .A0N(\ram[201][6] ), .A1N(n6409), 
        .Y(n3804) );
  OAI2BB2XL U1061 ( .B0(n6798), .B1(n378), .A0N(\ram[201][7] ), .A1N(n6409), 
        .Y(n3805) );
  OAI2BB2XL U1062 ( .B0(n6775), .B1(n378), .A0N(\ram[201][8] ), .A1N(n6409), 
        .Y(n3806) );
  OAI2BB2XL U1063 ( .B0(n6752), .B1(n378), .A0N(\ram[201][9] ), .A1N(n6409), 
        .Y(n3807) );
  OAI2BB2XL U1064 ( .B0(n6729), .B1(n378), .A0N(\ram[201][10] ), .A1N(n6409), 
        .Y(n3808) );
  OAI2BB2XL U1065 ( .B0(n6706), .B1(n378), .A0N(\ram[201][11] ), .A1N(n6409), 
        .Y(n3809) );
  OAI2BB2XL U1066 ( .B0(n6683), .B1(n378), .A0N(\ram[201][12] ), .A1N(n6409), 
        .Y(n3810) );
  OAI2BB2XL U1067 ( .B0(n6660), .B1(n378), .A0N(\ram[201][13] ), .A1N(n6409), 
        .Y(n3811) );
  OAI2BB2XL U1068 ( .B0(n6637), .B1(n378), .A0N(\ram[201][14] ), .A1N(n6409), 
        .Y(n3812) );
  OAI2BB2XL U1069 ( .B0(n6614), .B1(n378), .A0N(\ram[201][15] ), .A1N(n6409), 
        .Y(n3813) );
  OAI2BB2XL U1070 ( .B0(n6963), .B1(n380), .A0N(\ram[202][0] ), .A1N(n6408), 
        .Y(n3814) );
  OAI2BB2XL U1071 ( .B0(n6940), .B1(n380), .A0N(\ram[202][1] ), .A1N(n6408), 
        .Y(n3815) );
  OAI2BB2XL U1072 ( .B0(n6917), .B1(n380), .A0N(\ram[202][2] ), .A1N(n6408), 
        .Y(n3816) );
  OAI2BB2XL U1073 ( .B0(n6894), .B1(n380), .A0N(\ram[202][3] ), .A1N(n6408), 
        .Y(n3817) );
  OAI2BB2XL U1074 ( .B0(n6867), .B1(n380), .A0N(\ram[202][4] ), .A1N(n6408), 
        .Y(n3818) );
  OAI2BB2XL U1075 ( .B0(n6844), .B1(n380), .A0N(\ram[202][5] ), .A1N(n6408), 
        .Y(n3819) );
  OAI2BB2XL U1076 ( .B0(n6821), .B1(n380), .A0N(\ram[202][6] ), .A1N(n6408), 
        .Y(n3820) );
  OAI2BB2XL U1077 ( .B0(n6798), .B1(n380), .A0N(\ram[202][7] ), .A1N(n6408), 
        .Y(n3821) );
  OAI2BB2XL U1078 ( .B0(n6775), .B1(n380), .A0N(\ram[202][8] ), .A1N(n6408), 
        .Y(n3822) );
  OAI2BB2XL U1079 ( .B0(n6752), .B1(n380), .A0N(\ram[202][9] ), .A1N(n6408), 
        .Y(n3823) );
  OAI2BB2XL U1080 ( .B0(n6729), .B1(n380), .A0N(\ram[202][10] ), .A1N(n6408), 
        .Y(n3824) );
  OAI2BB2XL U1081 ( .B0(n6706), .B1(n380), .A0N(\ram[202][11] ), .A1N(n6408), 
        .Y(n3825) );
  OAI2BB2XL U1082 ( .B0(n6683), .B1(n380), .A0N(\ram[202][12] ), .A1N(n6408), 
        .Y(n3826) );
  OAI2BB2XL U1083 ( .B0(n6660), .B1(n380), .A0N(\ram[202][13] ), .A1N(n6408), 
        .Y(n3827) );
  OAI2BB2XL U1084 ( .B0(n6637), .B1(n380), .A0N(\ram[202][14] ), .A1N(n6408), 
        .Y(n3828) );
  OAI2BB2XL U1085 ( .B0(n6614), .B1(n380), .A0N(\ram[202][15] ), .A1N(n6408), 
        .Y(n3829) );
  OAI2BB2XL U1086 ( .B0(n6963), .B1(n382), .A0N(\ram[203][0] ), .A1N(n6407), 
        .Y(n3830) );
  OAI2BB2XL U1087 ( .B0(n6940), .B1(n382), .A0N(\ram[203][1] ), .A1N(n6407), 
        .Y(n3831) );
  OAI2BB2XL U1088 ( .B0(n6917), .B1(n382), .A0N(\ram[203][2] ), .A1N(n6407), 
        .Y(n3832) );
  OAI2BB2XL U1089 ( .B0(n6894), .B1(n382), .A0N(\ram[203][3] ), .A1N(n6407), 
        .Y(n3833) );
  OAI2BB2XL U1090 ( .B0(n6867), .B1(n382), .A0N(\ram[203][4] ), .A1N(n6407), 
        .Y(n3834) );
  OAI2BB2XL U1091 ( .B0(n6844), .B1(n382), .A0N(\ram[203][5] ), .A1N(n6407), 
        .Y(n3835) );
  OAI2BB2XL U1092 ( .B0(n6821), .B1(n382), .A0N(\ram[203][6] ), .A1N(n6407), 
        .Y(n3836) );
  OAI2BB2XL U1093 ( .B0(n6798), .B1(n382), .A0N(\ram[203][7] ), .A1N(n6407), 
        .Y(n3837) );
  OAI2BB2XL U1094 ( .B0(n6775), .B1(n382), .A0N(\ram[203][8] ), .A1N(n6407), 
        .Y(n3838) );
  OAI2BB2XL U1095 ( .B0(n6752), .B1(n382), .A0N(\ram[203][9] ), .A1N(n6407), 
        .Y(n3839) );
  OAI2BB2XL U1096 ( .B0(n6729), .B1(n382), .A0N(\ram[203][10] ), .A1N(n6407), 
        .Y(n3840) );
  OAI2BB2XL U1097 ( .B0(n6706), .B1(n382), .A0N(\ram[203][11] ), .A1N(n6407), 
        .Y(n3841) );
  OAI2BB2XL U1098 ( .B0(n6683), .B1(n382), .A0N(\ram[203][12] ), .A1N(n6407), 
        .Y(n3842) );
  OAI2BB2XL U1099 ( .B0(n6660), .B1(n382), .A0N(\ram[203][13] ), .A1N(n6407), 
        .Y(n3843) );
  OAI2BB2XL U1100 ( .B0(n6637), .B1(n382), .A0N(\ram[203][14] ), .A1N(n6407), 
        .Y(n3844) );
  OAI2BB2XL U1101 ( .B0(n6614), .B1(n382), .A0N(\ram[203][15] ), .A1N(n6407), 
        .Y(n3845) );
  OAI2BB2XL U1102 ( .B0(n6963), .B1(n384), .A0N(\ram[204][0] ), .A1N(n6406), 
        .Y(n3846) );
  OAI2BB2XL U1103 ( .B0(n6940), .B1(n384), .A0N(\ram[204][1] ), .A1N(n6406), 
        .Y(n3847) );
  OAI2BB2XL U1104 ( .B0(n6917), .B1(n384), .A0N(\ram[204][2] ), .A1N(n6406), 
        .Y(n3848) );
  OAI2BB2XL U1105 ( .B0(n6894), .B1(n384), .A0N(\ram[204][3] ), .A1N(n6406), 
        .Y(n3849) );
  OAI2BB2XL U1106 ( .B0(n6867), .B1(n384), .A0N(\ram[204][4] ), .A1N(n6406), 
        .Y(n3850) );
  OAI2BB2XL U1107 ( .B0(n6844), .B1(n384), .A0N(\ram[204][5] ), .A1N(n6406), 
        .Y(n3851) );
  OAI2BB2XL U1108 ( .B0(n6821), .B1(n384), .A0N(\ram[204][6] ), .A1N(n6406), 
        .Y(n3852) );
  OAI2BB2XL U1109 ( .B0(n6798), .B1(n384), .A0N(\ram[204][7] ), .A1N(n6406), 
        .Y(n3853) );
  OAI2BB2XL U1110 ( .B0(n6775), .B1(n384), .A0N(\ram[204][8] ), .A1N(n6406), 
        .Y(n3854) );
  OAI2BB2XL U1111 ( .B0(n6752), .B1(n384), .A0N(\ram[204][9] ), .A1N(n6406), 
        .Y(n3855) );
  OAI2BB2XL U1112 ( .B0(n6729), .B1(n384), .A0N(\ram[204][10] ), .A1N(n6406), 
        .Y(n3856) );
  OAI2BB2XL U1113 ( .B0(n6706), .B1(n384), .A0N(\ram[204][11] ), .A1N(n6406), 
        .Y(n3857) );
  OAI2BB2XL U1114 ( .B0(n6683), .B1(n384), .A0N(\ram[204][12] ), .A1N(n6406), 
        .Y(n3858) );
  OAI2BB2XL U1115 ( .B0(n6660), .B1(n384), .A0N(\ram[204][13] ), .A1N(n6406), 
        .Y(n3859) );
  OAI2BB2XL U1116 ( .B0(n6637), .B1(n384), .A0N(\ram[204][14] ), .A1N(n6406), 
        .Y(n3860) );
  OAI2BB2XL U1117 ( .B0(n6614), .B1(n384), .A0N(\ram[204][15] ), .A1N(n6406), 
        .Y(n3861) );
  OAI2BB2XL U1118 ( .B0(n6963), .B1(n386), .A0N(\ram[205][0] ), .A1N(n6405), 
        .Y(n3862) );
  OAI2BB2XL U1119 ( .B0(n6940), .B1(n386), .A0N(\ram[205][1] ), .A1N(n6405), 
        .Y(n3863) );
  OAI2BB2XL U1120 ( .B0(n6917), .B1(n386), .A0N(\ram[205][2] ), .A1N(n6405), 
        .Y(n3864) );
  OAI2BB2XL U1121 ( .B0(n6894), .B1(n386), .A0N(\ram[205][3] ), .A1N(n6405), 
        .Y(n3865) );
  OAI2BB2XL U1122 ( .B0(n6867), .B1(n386), .A0N(\ram[205][4] ), .A1N(n6405), 
        .Y(n3866) );
  OAI2BB2XL U1123 ( .B0(n6844), .B1(n386), .A0N(\ram[205][5] ), .A1N(n6405), 
        .Y(n3867) );
  OAI2BB2XL U1124 ( .B0(n6821), .B1(n386), .A0N(\ram[205][6] ), .A1N(n6405), 
        .Y(n3868) );
  OAI2BB2XL U1125 ( .B0(n6798), .B1(n386), .A0N(\ram[205][7] ), .A1N(n6405), 
        .Y(n3869) );
  OAI2BB2XL U1126 ( .B0(n6775), .B1(n386), .A0N(\ram[205][8] ), .A1N(n6405), 
        .Y(n3870) );
  OAI2BB2XL U1127 ( .B0(n6752), .B1(n386), .A0N(\ram[205][9] ), .A1N(n6405), 
        .Y(n3871) );
  OAI2BB2XL U1128 ( .B0(n6729), .B1(n386), .A0N(\ram[205][10] ), .A1N(n6405), 
        .Y(n3872) );
  OAI2BB2XL U1129 ( .B0(n6706), .B1(n386), .A0N(\ram[205][11] ), .A1N(n6405), 
        .Y(n3873) );
  OAI2BB2XL U1130 ( .B0(n6683), .B1(n386), .A0N(\ram[205][12] ), .A1N(n6405), 
        .Y(n3874) );
  OAI2BB2XL U1131 ( .B0(n6660), .B1(n386), .A0N(\ram[205][13] ), .A1N(n6405), 
        .Y(n3875) );
  OAI2BB2XL U1132 ( .B0(n6637), .B1(n386), .A0N(\ram[205][14] ), .A1N(n6405), 
        .Y(n3876) );
  OAI2BB2XL U1133 ( .B0(n6614), .B1(n386), .A0N(\ram[205][15] ), .A1N(n6405), 
        .Y(n3877) );
  OAI2BB2XL U1134 ( .B0(n6963), .B1(n388), .A0N(\ram[206][0] ), .A1N(n6404), 
        .Y(n3878) );
  OAI2BB2XL U1135 ( .B0(n6940), .B1(n388), .A0N(\ram[206][1] ), .A1N(n6404), 
        .Y(n3879) );
  OAI2BB2XL U1136 ( .B0(n6917), .B1(n388), .A0N(\ram[206][2] ), .A1N(n6404), 
        .Y(n3880) );
  OAI2BB2XL U1137 ( .B0(n6894), .B1(n388), .A0N(\ram[206][3] ), .A1N(n6404), 
        .Y(n3881) );
  OAI2BB2XL U1138 ( .B0(n6867), .B1(n388), .A0N(\ram[206][4] ), .A1N(n6404), 
        .Y(n3882) );
  OAI2BB2XL U1139 ( .B0(n6844), .B1(n388), .A0N(\ram[206][5] ), .A1N(n6404), 
        .Y(n3883) );
  OAI2BB2XL U1140 ( .B0(n6821), .B1(n388), .A0N(\ram[206][6] ), .A1N(n6404), 
        .Y(n3884) );
  OAI2BB2XL U1141 ( .B0(n6798), .B1(n388), .A0N(\ram[206][7] ), .A1N(n6404), 
        .Y(n3885) );
  OAI2BB2XL U1142 ( .B0(n6775), .B1(n388), .A0N(\ram[206][8] ), .A1N(n6404), 
        .Y(n3886) );
  OAI2BB2XL U1143 ( .B0(n6752), .B1(n388), .A0N(\ram[206][9] ), .A1N(n6404), 
        .Y(n3887) );
  OAI2BB2XL U1144 ( .B0(n6729), .B1(n388), .A0N(\ram[206][10] ), .A1N(n6404), 
        .Y(n3888) );
  OAI2BB2XL U1145 ( .B0(n6706), .B1(n388), .A0N(\ram[206][11] ), .A1N(n6404), 
        .Y(n3889) );
  OAI2BB2XL U1146 ( .B0(n6683), .B1(n388), .A0N(\ram[206][12] ), .A1N(n6404), 
        .Y(n3890) );
  OAI2BB2XL U1147 ( .B0(n6660), .B1(n388), .A0N(\ram[206][13] ), .A1N(n6404), 
        .Y(n3891) );
  OAI2BB2XL U1148 ( .B0(n6637), .B1(n388), .A0N(\ram[206][14] ), .A1N(n6404), 
        .Y(n3892) );
  OAI2BB2XL U1149 ( .B0(n6614), .B1(n388), .A0N(\ram[206][15] ), .A1N(n6404), 
        .Y(n3893) );
  OAI2BB2XL U1150 ( .B0(n6963), .B1(n390), .A0N(\ram[207][0] ), .A1N(n6403), 
        .Y(n3894) );
  OAI2BB2XL U1151 ( .B0(n6940), .B1(n390), .A0N(\ram[207][1] ), .A1N(n6403), 
        .Y(n3895) );
  OAI2BB2XL U1152 ( .B0(n6917), .B1(n390), .A0N(\ram[207][2] ), .A1N(n6403), 
        .Y(n3896) );
  OAI2BB2XL U1153 ( .B0(n6894), .B1(n390), .A0N(\ram[207][3] ), .A1N(n6403), 
        .Y(n3897) );
  OAI2BB2XL U1154 ( .B0(n6867), .B1(n390), .A0N(\ram[207][4] ), .A1N(n6403), 
        .Y(n3898) );
  OAI2BB2XL U1155 ( .B0(n6844), .B1(n390), .A0N(\ram[207][5] ), .A1N(n6403), 
        .Y(n3899) );
  OAI2BB2XL U1156 ( .B0(n6821), .B1(n390), .A0N(\ram[207][6] ), .A1N(n6403), 
        .Y(n3900) );
  OAI2BB2XL U1157 ( .B0(n6798), .B1(n390), .A0N(\ram[207][7] ), .A1N(n6403), 
        .Y(n3901) );
  OAI2BB2XL U1158 ( .B0(n6775), .B1(n390), .A0N(\ram[207][8] ), .A1N(n6403), 
        .Y(n3902) );
  OAI2BB2XL U1159 ( .B0(n6752), .B1(n390), .A0N(\ram[207][9] ), .A1N(n6403), 
        .Y(n3903) );
  OAI2BB2XL U1160 ( .B0(n6729), .B1(n390), .A0N(\ram[207][10] ), .A1N(n6403), 
        .Y(n3904) );
  OAI2BB2XL U1161 ( .B0(n6706), .B1(n390), .A0N(\ram[207][11] ), .A1N(n6403), 
        .Y(n3905) );
  OAI2BB2XL U1162 ( .B0(n6683), .B1(n390), .A0N(\ram[207][12] ), .A1N(n6403), 
        .Y(n3906) );
  OAI2BB2XL U1163 ( .B0(n6660), .B1(n390), .A0N(\ram[207][13] ), .A1N(n6403), 
        .Y(n3907) );
  OAI2BB2XL U1164 ( .B0(n6637), .B1(n390), .A0N(\ram[207][14] ), .A1N(n6403), 
        .Y(n3908) );
  OAI2BB2XL U1165 ( .B0(n6614), .B1(n390), .A0N(\ram[207][15] ), .A1N(n6403), 
        .Y(n3909) );
  OAI2BB2XL U1166 ( .B0(n21), .B1(n7), .A0N(\ram[0][0] ), .A1N(n6610), .Y(n582) );
  OAI2BB2XL U1167 ( .B0(n21), .B1(n9), .A0N(\ram[0][1] ), .A1N(n6610), .Y(n583) );
  OAI2BB2XL U1168 ( .B0(n21), .B1(n10), .A0N(\ram[0][2] ), .A1N(n6610), .Y(
        n584) );
  OAI2BB2XL U1169 ( .B0(n21), .B1(n11), .A0N(\ram[0][3] ), .A1N(n6610), .Y(
        n585) );
  OAI2BB2XL U1170 ( .B0(n21), .B1(n6878), .A0N(\ram[0][4] ), .A1N(n6610), .Y(
        n586) );
  OAI2BB2XL U1171 ( .B0(n21), .B1(n6855), .A0N(\ram[0][5] ), .A1N(n6610), .Y(
        n587) );
  OAI2BB2XL U1172 ( .B0(n21), .B1(n6832), .A0N(\ram[0][6] ), .A1N(n6610), .Y(
        n588) );
  OAI2BB2XL U1173 ( .B0(n21), .B1(n6809), .A0N(\ram[0][7] ), .A1N(n6610), .Y(
        n589) );
  OAI2BB2XL U1174 ( .B0(n21), .B1(n6786), .A0N(\ram[0][8] ), .A1N(n6610), .Y(
        n590) );
  OAI2BB2XL U1175 ( .B0(n21), .B1(n6763), .A0N(\ram[0][9] ), .A1N(n6610), .Y(
        n591) );
  OAI2BB2XL U1176 ( .B0(n21), .B1(n6740), .A0N(\ram[0][10] ), .A1N(n6610), .Y(
        n592) );
  OAI2BB2XL U1177 ( .B0(n21), .B1(n6717), .A0N(\ram[0][11] ), .A1N(n6610), .Y(
        n593) );
  OAI2BB2XL U1178 ( .B0(n21), .B1(n6694), .A0N(\ram[0][12] ), .A1N(n6610), .Y(
        n594) );
  OAI2BB2XL U1179 ( .B0(n21), .B1(n6671), .A0N(\ram[0][13] ), .A1N(n6610), .Y(
        n595) );
  OAI2BB2XL U1180 ( .B0(n21), .B1(n6648), .A0N(\ram[0][14] ), .A1N(n6610), .Y(
        n596) );
  OAI2BB2XL U1181 ( .B0(n21), .B1(n6625), .A0N(\ram[0][15] ), .A1N(n6610), .Y(
        n597) );
  OAI2BB2XL U1182 ( .B0(n6969), .B1(n41), .A0N(\ram[5][0] ), .A1N(n6605), .Y(
        n662) );
  OAI2BB2XL U1183 ( .B0(n6946), .B1(n41), .A0N(\ram[5][1] ), .A1N(n6605), .Y(
        n663) );
  OAI2BB2XL U1184 ( .B0(n6923), .B1(n41), .A0N(\ram[5][2] ), .A1N(n6605), .Y(
        n664) );
  OAI2BB2XL U1185 ( .B0(n6900), .B1(n41), .A0N(\ram[5][3] ), .A1N(n6605), .Y(
        n665) );
  OAI2BB2XL U1186 ( .B0(n6882), .B1(n41), .A0N(\ram[5][4] ), .A1N(n6605), .Y(
        n666) );
  OAI2BB2XL U1187 ( .B0(n6859), .B1(n41), .A0N(\ram[5][5] ), .A1N(n6605), .Y(
        n667) );
  OAI2BB2XL U1188 ( .B0(n6836), .B1(n41), .A0N(\ram[5][6] ), .A1N(n6605), .Y(
        n668) );
  OAI2BB2XL U1189 ( .B0(n6813), .B1(n41), .A0N(\ram[5][7] ), .A1N(n6605), .Y(
        n669) );
  OAI2BB2XL U1190 ( .B0(n6790), .B1(n41), .A0N(\ram[5][8] ), .A1N(n6605), .Y(
        n670) );
  OAI2BB2XL U1191 ( .B0(n6767), .B1(n41), .A0N(\ram[5][9] ), .A1N(n6605), .Y(
        n671) );
  OAI2BB2XL U1192 ( .B0(n6744), .B1(n41), .A0N(\ram[5][10] ), .A1N(n6605), .Y(
        n672) );
  OAI2BB2XL U1193 ( .B0(n6721), .B1(n41), .A0N(\ram[5][11] ), .A1N(n6605), .Y(
        n673) );
  OAI2BB2XL U1194 ( .B0(n6698), .B1(n41), .A0N(\ram[5][12] ), .A1N(n6605), .Y(
        n674) );
  OAI2BB2XL U1195 ( .B0(n6675), .B1(n41), .A0N(\ram[5][13] ), .A1N(n6605), .Y(
        n675) );
  OAI2BB2XL U1196 ( .B0(n6652), .B1(n41), .A0N(\ram[5][14] ), .A1N(n6605), .Y(
        n676) );
  OAI2BB2XL U1197 ( .B0(n6629), .B1(n41), .A0N(\ram[5][15] ), .A1N(n6605), .Y(
        n677) );
  OAI2BB2XL U1198 ( .B0(n6960), .B1(n43), .A0N(\ram[6][0] ), .A1N(n6604), .Y(
        n678) );
  OAI2BB2XL U1199 ( .B0(n6937), .B1(n43), .A0N(\ram[6][1] ), .A1N(n6604), .Y(
        n679) );
  OAI2BB2XL U1200 ( .B0(n6914), .B1(n43), .A0N(\ram[6][2] ), .A1N(n6604), .Y(
        n680) );
  OAI2BB2XL U1201 ( .B0(n6891), .B1(n43), .A0N(\ram[6][3] ), .A1N(n6604), .Y(
        n681) );
  OAI2BB2XL U1202 ( .B0(n6882), .B1(n43), .A0N(\ram[6][4] ), .A1N(n6604), .Y(
        n682) );
  OAI2BB2XL U1203 ( .B0(n6859), .B1(n43), .A0N(\ram[6][5] ), .A1N(n6604), .Y(
        n683) );
  OAI2BB2XL U1204 ( .B0(n6836), .B1(n43), .A0N(\ram[6][6] ), .A1N(n6604), .Y(
        n684) );
  OAI2BB2XL U1205 ( .B0(n6813), .B1(n43), .A0N(\ram[6][7] ), .A1N(n6604), .Y(
        n685) );
  OAI2BB2XL U1206 ( .B0(n6790), .B1(n43), .A0N(\ram[6][8] ), .A1N(n6604), .Y(
        n686) );
  OAI2BB2XL U1207 ( .B0(n6767), .B1(n43), .A0N(\ram[6][9] ), .A1N(n6604), .Y(
        n687) );
  OAI2BB2XL U1208 ( .B0(n6744), .B1(n43), .A0N(\ram[6][10] ), .A1N(n6604), .Y(
        n688) );
  OAI2BB2XL U1209 ( .B0(n6721), .B1(n43), .A0N(\ram[6][11] ), .A1N(n6604), .Y(
        n689) );
  OAI2BB2XL U1210 ( .B0(n6698), .B1(n43), .A0N(\ram[6][12] ), .A1N(n6604), .Y(
        n690) );
  OAI2BB2XL U1211 ( .B0(n6675), .B1(n43), .A0N(\ram[6][13] ), .A1N(n6604), .Y(
        n691) );
  OAI2BB2XL U1212 ( .B0(n6652), .B1(n43), .A0N(\ram[6][14] ), .A1N(n6604), .Y(
        n692) );
  OAI2BB2XL U1213 ( .B0(n6629), .B1(n43), .A0N(\ram[6][15] ), .A1N(n6604), .Y(
        n693) );
  OAI2BB2XL U1214 ( .B0(n6959), .B1(n44), .A0N(\ram[7][0] ), .A1N(n6603), .Y(
        n694) );
  OAI2BB2XL U1215 ( .B0(n6936), .B1(n44), .A0N(\ram[7][1] ), .A1N(n6603), .Y(
        n695) );
  OAI2BB2XL U1216 ( .B0(n6913), .B1(n44), .A0N(\ram[7][2] ), .A1N(n6603), .Y(
        n696) );
  OAI2BB2XL U1217 ( .B0(n6890), .B1(n44), .A0N(\ram[7][3] ), .A1N(n6603), .Y(
        n697) );
  OAI2BB2XL U1218 ( .B0(n6882), .B1(n44), .A0N(\ram[7][4] ), .A1N(n6603), .Y(
        n698) );
  OAI2BB2XL U1219 ( .B0(n6859), .B1(n44), .A0N(\ram[7][5] ), .A1N(n6603), .Y(
        n699) );
  OAI2BB2XL U1220 ( .B0(n6836), .B1(n44), .A0N(\ram[7][6] ), .A1N(n6603), .Y(
        n700) );
  OAI2BB2XL U1221 ( .B0(n6813), .B1(n44), .A0N(\ram[7][7] ), .A1N(n6603), .Y(
        n701) );
  OAI2BB2XL U1222 ( .B0(n6790), .B1(n44), .A0N(\ram[7][8] ), .A1N(n6603), .Y(
        n702) );
  OAI2BB2XL U1223 ( .B0(n6767), .B1(n44), .A0N(\ram[7][9] ), .A1N(n6603), .Y(
        n703) );
  OAI2BB2XL U1224 ( .B0(n6744), .B1(n44), .A0N(\ram[7][10] ), .A1N(n6603), .Y(
        n704) );
  OAI2BB2XL U1225 ( .B0(n6721), .B1(n44), .A0N(\ram[7][11] ), .A1N(n6603), .Y(
        n705) );
  OAI2BB2XL U1226 ( .B0(n6698), .B1(n44), .A0N(\ram[7][12] ), .A1N(n6603), .Y(
        n706) );
  OAI2BB2XL U1227 ( .B0(n6675), .B1(n44), .A0N(\ram[7][13] ), .A1N(n6603), .Y(
        n707) );
  OAI2BB2XL U1228 ( .B0(n6652), .B1(n44), .A0N(\ram[7][14] ), .A1N(n6603), .Y(
        n708) );
  OAI2BB2XL U1229 ( .B0(n6629), .B1(n44), .A0N(\ram[7][15] ), .A1N(n6603), .Y(
        n709) );
  OAI2BB2XL U1230 ( .B0(n6974), .B1(n47), .A0N(\ram[9][0] ), .A1N(n6601), .Y(
        n726) );
  OAI2BB2XL U1231 ( .B0(n6951), .B1(n47), .A0N(\ram[9][1] ), .A1N(n6601), .Y(
        n727) );
  OAI2BB2XL U1232 ( .B0(n6928), .B1(n47), .A0N(\ram[9][2] ), .A1N(n6601), .Y(
        n728) );
  OAI2BB2XL U1233 ( .B0(n6905), .B1(n47), .A0N(\ram[9][3] ), .A1N(n6601), .Y(
        n729) );
  OAI2BB2XL U1234 ( .B0(n6882), .B1(n47), .A0N(\ram[9][4] ), .A1N(n6601), .Y(
        n730) );
  OAI2BB2XL U1235 ( .B0(n6859), .B1(n47), .A0N(\ram[9][5] ), .A1N(n6601), .Y(
        n731) );
  OAI2BB2XL U1236 ( .B0(n6836), .B1(n47), .A0N(\ram[9][6] ), .A1N(n6601), .Y(
        n732) );
  OAI2BB2XL U1237 ( .B0(n6813), .B1(n47), .A0N(\ram[9][7] ), .A1N(n6601), .Y(
        n733) );
  OAI2BB2XL U1238 ( .B0(n6790), .B1(n47), .A0N(\ram[9][8] ), .A1N(n6601), .Y(
        n734) );
  OAI2BB2XL U1239 ( .B0(n6767), .B1(n47), .A0N(\ram[9][9] ), .A1N(n6601), .Y(
        n735) );
  OAI2BB2XL U1240 ( .B0(n6744), .B1(n47), .A0N(\ram[9][10] ), .A1N(n6601), .Y(
        n736) );
  OAI2BB2XL U1241 ( .B0(n6721), .B1(n47), .A0N(\ram[9][11] ), .A1N(n6601), .Y(
        n737) );
  OAI2BB2XL U1242 ( .B0(n6698), .B1(n47), .A0N(\ram[9][12] ), .A1N(n6601), .Y(
        n738) );
  OAI2BB2XL U1243 ( .B0(n6675), .B1(n47), .A0N(\ram[9][13] ), .A1N(n6601), .Y(
        n739) );
  OAI2BB2XL U1244 ( .B0(n6652), .B1(n47), .A0N(\ram[9][14] ), .A1N(n6601), .Y(
        n740) );
  OAI2BB2XL U1245 ( .B0(n6629), .B1(n47), .A0N(\ram[9][15] ), .A1N(n6601), .Y(
        n741) );
  OAI2BB2XL U1246 ( .B0(n6973), .B1(n49), .A0N(\ram[10][0] ), .A1N(n6600), .Y(
        n742) );
  OAI2BB2XL U1247 ( .B0(n6950), .B1(n49), .A0N(\ram[10][1] ), .A1N(n6600), .Y(
        n743) );
  OAI2BB2XL U1248 ( .B0(n6927), .B1(n49), .A0N(\ram[10][2] ), .A1N(n6600), .Y(
        n744) );
  OAI2BB2XL U1249 ( .B0(n6904), .B1(n49), .A0N(\ram[10][3] ), .A1N(n6600), .Y(
        n745) );
  OAI2BB2XL U1250 ( .B0(n6882), .B1(n49), .A0N(\ram[10][4] ), .A1N(n6600), .Y(
        n746) );
  OAI2BB2XL U1251 ( .B0(n6859), .B1(n49), .A0N(\ram[10][5] ), .A1N(n6600), .Y(
        n747) );
  OAI2BB2XL U1252 ( .B0(n6836), .B1(n49), .A0N(\ram[10][6] ), .A1N(n6600), .Y(
        n748) );
  OAI2BB2XL U1253 ( .B0(n6813), .B1(n49), .A0N(\ram[10][7] ), .A1N(n6600), .Y(
        n749) );
  OAI2BB2XL U1254 ( .B0(n6790), .B1(n49), .A0N(\ram[10][8] ), .A1N(n6600), .Y(
        n750) );
  OAI2BB2XL U1255 ( .B0(n6767), .B1(n49), .A0N(\ram[10][9] ), .A1N(n6600), .Y(
        n751) );
  OAI2BB2XL U1256 ( .B0(n6744), .B1(n49), .A0N(\ram[10][10] ), .A1N(n6600), 
        .Y(n752) );
  OAI2BB2XL U1257 ( .B0(n6721), .B1(n49), .A0N(\ram[10][11] ), .A1N(n6600), 
        .Y(n753) );
  OAI2BB2XL U1258 ( .B0(n6698), .B1(n49), .A0N(\ram[10][12] ), .A1N(n6600), 
        .Y(n754) );
  OAI2BB2XL U1259 ( .B0(n6675), .B1(n49), .A0N(\ram[10][13] ), .A1N(n6600), 
        .Y(n755) );
  OAI2BB2XL U1260 ( .B0(n6652), .B1(n49), .A0N(\ram[10][14] ), .A1N(n6600), 
        .Y(n756) );
  OAI2BB2XL U1261 ( .B0(n6629), .B1(n49), .A0N(\ram[10][15] ), .A1N(n6600), 
        .Y(n757) );
  OAI2BB2XL U1262 ( .B0(n6972), .B1(n50), .A0N(\ram[11][0] ), .A1N(n6599), .Y(
        n758) );
  OAI2BB2XL U1263 ( .B0(n6949), .B1(n50), .A0N(\ram[11][1] ), .A1N(n6599), .Y(
        n759) );
  OAI2BB2XL U1264 ( .B0(n6926), .B1(n50), .A0N(\ram[11][2] ), .A1N(n6599), .Y(
        n760) );
  OAI2BB2XL U1265 ( .B0(n6903), .B1(n50), .A0N(\ram[11][3] ), .A1N(n6599), .Y(
        n761) );
  OAI2BB2XL U1266 ( .B0(n6882), .B1(n50), .A0N(\ram[11][4] ), .A1N(n6599), .Y(
        n762) );
  OAI2BB2XL U1267 ( .B0(n6859), .B1(n50), .A0N(\ram[11][5] ), .A1N(n6599), .Y(
        n763) );
  OAI2BB2XL U1268 ( .B0(n6836), .B1(n50), .A0N(\ram[11][6] ), .A1N(n6599), .Y(
        n764) );
  OAI2BB2XL U1269 ( .B0(n6813), .B1(n50), .A0N(\ram[11][7] ), .A1N(n6599), .Y(
        n765) );
  OAI2BB2XL U1270 ( .B0(n6790), .B1(n50), .A0N(\ram[11][8] ), .A1N(n6599), .Y(
        n766) );
  OAI2BB2XL U1271 ( .B0(n6767), .B1(n50), .A0N(\ram[11][9] ), .A1N(n6599), .Y(
        n767) );
  OAI2BB2XL U1272 ( .B0(n6744), .B1(n50), .A0N(\ram[11][10] ), .A1N(n6599), 
        .Y(n768) );
  OAI2BB2XL U1273 ( .B0(n6721), .B1(n50), .A0N(\ram[11][11] ), .A1N(n6599), 
        .Y(n769) );
  OAI2BB2XL U1274 ( .B0(n6698), .B1(n50), .A0N(\ram[11][12] ), .A1N(n6599), 
        .Y(n770) );
  OAI2BB2XL U1275 ( .B0(n6675), .B1(n50), .A0N(\ram[11][13] ), .A1N(n6599), 
        .Y(n771) );
  OAI2BB2XL U1276 ( .B0(n6652), .B1(n50), .A0N(\ram[11][14] ), .A1N(n6599), 
        .Y(n772) );
  OAI2BB2XL U1277 ( .B0(n6629), .B1(n50), .A0N(\ram[11][15] ), .A1N(n6599), 
        .Y(n773) );
  OAI2BB2XL U1278 ( .B0(n6971), .B1(n53), .A0N(\ram[13][0] ), .A1N(n6597), .Y(
        n790) );
  OAI2BB2XL U1279 ( .B0(n6948), .B1(n53), .A0N(\ram[13][1] ), .A1N(n6597), .Y(
        n791) );
  OAI2BB2XL U1280 ( .B0(n6925), .B1(n53), .A0N(\ram[13][2] ), .A1N(n6597), .Y(
        n792) );
  OAI2BB2XL U1281 ( .B0(n6902), .B1(n53), .A0N(\ram[13][3] ), .A1N(n6597), .Y(
        n793) );
  OAI2BB2XL U1282 ( .B0(n6882), .B1(n53), .A0N(\ram[13][4] ), .A1N(n6597), .Y(
        n794) );
  OAI2BB2XL U1283 ( .B0(n6859), .B1(n53), .A0N(\ram[13][5] ), .A1N(n6597), .Y(
        n795) );
  OAI2BB2XL U1284 ( .B0(n6836), .B1(n53), .A0N(\ram[13][6] ), .A1N(n6597), .Y(
        n796) );
  OAI2BB2XL U1285 ( .B0(n6813), .B1(n53), .A0N(\ram[13][7] ), .A1N(n6597), .Y(
        n797) );
  OAI2BB2XL U1286 ( .B0(n6790), .B1(n53), .A0N(\ram[13][8] ), .A1N(n6597), .Y(
        n798) );
  OAI2BB2XL U1287 ( .B0(n6767), .B1(n53), .A0N(\ram[13][9] ), .A1N(n6597), .Y(
        n799) );
  OAI2BB2XL U1288 ( .B0(n6744), .B1(n53), .A0N(\ram[13][10] ), .A1N(n6597), 
        .Y(n800) );
  OAI2BB2XL U1289 ( .B0(n6721), .B1(n53), .A0N(\ram[13][11] ), .A1N(n6597), 
        .Y(n801) );
  OAI2BB2XL U1290 ( .B0(n6698), .B1(n53), .A0N(\ram[13][12] ), .A1N(n6597), 
        .Y(n802) );
  OAI2BB2XL U1291 ( .B0(n6675), .B1(n53), .A0N(\ram[13][13] ), .A1N(n6597), 
        .Y(n803) );
  OAI2BB2XL U1292 ( .B0(n6652), .B1(n53), .A0N(\ram[13][14] ), .A1N(n6597), 
        .Y(n804) );
  OAI2BB2XL U1293 ( .B0(n6629), .B1(n53), .A0N(\ram[13][15] ), .A1N(n6597), 
        .Y(n805) );
  OAI2BB2XL U1294 ( .B0(n6970), .B1(n494), .A0N(\ram[14][0] ), .A1N(n6596), 
        .Y(n806) );
  OAI2BB2XL U1295 ( .B0(n6947), .B1(n494), .A0N(\ram[14][1] ), .A1N(n6596), 
        .Y(n807) );
  OAI2BB2XL U1296 ( .B0(n6924), .B1(n494), .A0N(\ram[14][2] ), .A1N(n6596), 
        .Y(n808) );
  OAI2BB2XL U1297 ( .B0(n6901), .B1(n494), .A0N(\ram[14][3] ), .A1N(n6596), 
        .Y(n809) );
  OAI2BB2XL U1298 ( .B0(n6882), .B1(n494), .A0N(\ram[14][4] ), .A1N(n6596), 
        .Y(n810) );
  OAI2BB2XL U1299 ( .B0(n6859), .B1(n494), .A0N(\ram[14][5] ), .A1N(n6596), 
        .Y(n811) );
  OAI2BB2XL U1300 ( .B0(n6836), .B1(n494), .A0N(\ram[14][6] ), .A1N(n6596), 
        .Y(n812) );
  OAI2BB2XL U1301 ( .B0(n6813), .B1(n494), .A0N(\ram[14][7] ), .A1N(n6596), 
        .Y(n813) );
  OAI2BB2XL U1302 ( .B0(n6790), .B1(n494), .A0N(\ram[14][8] ), .A1N(n6596), 
        .Y(n814) );
  OAI2BB2XL U1303 ( .B0(n6767), .B1(n494), .A0N(\ram[14][9] ), .A1N(n6596), 
        .Y(n815) );
  OAI2BB2XL U1304 ( .B0(n6744), .B1(n494), .A0N(\ram[14][10] ), .A1N(n6596), 
        .Y(n816) );
  OAI2BB2XL U1305 ( .B0(n6721), .B1(n494), .A0N(\ram[14][11] ), .A1N(n6596), 
        .Y(n817) );
  OAI2BB2XL U1306 ( .B0(n6698), .B1(n494), .A0N(\ram[14][12] ), .A1N(n6596), 
        .Y(n818) );
  OAI2BB2XL U1307 ( .B0(n6675), .B1(n494), .A0N(\ram[14][13] ), .A1N(n6596), 
        .Y(n819) );
  OAI2BB2XL U1308 ( .B0(n6652), .B1(n494), .A0N(\ram[14][14] ), .A1N(n6596), 
        .Y(n820) );
  OAI2BB2XL U1309 ( .B0(n6629), .B1(n494), .A0N(\ram[14][15] ), .A1N(n6596), 
        .Y(n821) );
  OAI2BB2XL U1310 ( .B0(n6969), .B1(n55), .A0N(\ram[15][0] ), .A1N(n6595), .Y(
        n822) );
  OAI2BB2XL U1311 ( .B0(n6946), .B1(n55), .A0N(\ram[15][1] ), .A1N(n6595), .Y(
        n823) );
  OAI2BB2XL U1312 ( .B0(n6923), .B1(n55), .A0N(\ram[15][2] ), .A1N(n6595), .Y(
        n824) );
  OAI2BB2XL U1313 ( .B0(n6900), .B1(n55), .A0N(\ram[15][3] ), .A1N(n6595), .Y(
        n825) );
  OAI2BB2XL U1314 ( .B0(n6882), .B1(n55), .A0N(\ram[15][4] ), .A1N(n6595), .Y(
        n826) );
  OAI2BB2XL U1315 ( .B0(n6859), .B1(n55), .A0N(\ram[15][5] ), .A1N(n6595), .Y(
        n827) );
  OAI2BB2XL U1316 ( .B0(n6836), .B1(n55), .A0N(\ram[15][6] ), .A1N(n6595), .Y(
        n828) );
  OAI2BB2XL U1317 ( .B0(n6813), .B1(n55), .A0N(\ram[15][7] ), .A1N(n6595), .Y(
        n829) );
  OAI2BB2XL U1318 ( .B0(n6790), .B1(n55), .A0N(\ram[15][8] ), .A1N(n6595), .Y(
        n830) );
  OAI2BB2XL U1319 ( .B0(n6767), .B1(n55), .A0N(\ram[15][9] ), .A1N(n6595), .Y(
        n831) );
  OAI2BB2XL U1320 ( .B0(n6744), .B1(n55), .A0N(\ram[15][10] ), .A1N(n6595), 
        .Y(n832) );
  OAI2BB2XL U1321 ( .B0(n6721), .B1(n55), .A0N(\ram[15][11] ), .A1N(n6595), 
        .Y(n833) );
  OAI2BB2XL U1322 ( .B0(n6698), .B1(n55), .A0N(\ram[15][12] ), .A1N(n6595), 
        .Y(n834) );
  OAI2BB2XL U1323 ( .B0(n6675), .B1(n55), .A0N(\ram[15][13] ), .A1N(n6595), 
        .Y(n835) );
  OAI2BB2XL U1324 ( .B0(n6652), .B1(n55), .A0N(\ram[15][14] ), .A1N(n6595), 
        .Y(n836) );
  OAI2BB2XL U1325 ( .B0(n6629), .B1(n55), .A0N(\ram[15][15] ), .A1N(n6595), 
        .Y(n837) );
  OAI2BB2XL U1326 ( .B0(n6961), .B1(n56), .A0N(\ram[16][0] ), .A1N(n6594), .Y(
        n838) );
  OAI2BB2XL U1327 ( .B0(n6938), .B1(n56), .A0N(\ram[16][1] ), .A1N(n6594), .Y(
        n839) );
  OAI2BB2XL U1328 ( .B0(n6915), .B1(n56), .A0N(\ram[16][2] ), .A1N(n6594), .Y(
        n840) );
  OAI2BB2XL U1329 ( .B0(n6892), .B1(n56), .A0N(\ram[16][3] ), .A1N(n6594), .Y(
        n841) );
  OAI2BB2XL U1330 ( .B0(n6881), .B1(n56), .A0N(\ram[16][4] ), .A1N(n6594), .Y(
        n842) );
  OAI2BB2XL U1331 ( .B0(n6858), .B1(n56), .A0N(\ram[16][5] ), .A1N(n6594), .Y(
        n843) );
  OAI2BB2XL U1332 ( .B0(n6835), .B1(n56), .A0N(\ram[16][6] ), .A1N(n6594), .Y(
        n844) );
  OAI2BB2XL U1333 ( .B0(n6812), .B1(n56), .A0N(\ram[16][7] ), .A1N(n6594), .Y(
        n845) );
  OAI2BB2XL U1334 ( .B0(n6789), .B1(n56), .A0N(\ram[16][8] ), .A1N(n6594), .Y(
        n846) );
  OAI2BB2XL U1335 ( .B0(n6766), .B1(n56), .A0N(\ram[16][9] ), .A1N(n6594), .Y(
        n847) );
  OAI2BB2XL U1336 ( .B0(n6743), .B1(n56), .A0N(\ram[16][10] ), .A1N(n6594), 
        .Y(n848) );
  OAI2BB2XL U1337 ( .B0(n6720), .B1(n56), .A0N(\ram[16][11] ), .A1N(n6594), 
        .Y(n849) );
  OAI2BB2XL U1338 ( .B0(n6697), .B1(n56), .A0N(\ram[16][12] ), .A1N(n6594), 
        .Y(n850) );
  OAI2BB2XL U1339 ( .B0(n6674), .B1(n56), .A0N(\ram[16][13] ), .A1N(n6594), 
        .Y(n851) );
  OAI2BB2XL U1340 ( .B0(n6651), .B1(n56), .A0N(\ram[16][14] ), .A1N(n6594), 
        .Y(n852) );
  OAI2BB2XL U1341 ( .B0(n6628), .B1(n56), .A0N(\ram[16][15] ), .A1N(n6594), 
        .Y(n853) );
  OAI2BB2XL U1342 ( .B0(n6968), .B1(n58), .A0N(\ram[17][0] ), .A1N(n6593), .Y(
        n854) );
  OAI2BB2XL U1343 ( .B0(n6945), .B1(n58), .A0N(\ram[17][1] ), .A1N(n6593), .Y(
        n855) );
  OAI2BB2XL U1344 ( .B0(n6922), .B1(n58), .A0N(\ram[17][2] ), .A1N(n6593), .Y(
        n856) );
  OAI2BB2XL U1345 ( .B0(n6899), .B1(n58), .A0N(\ram[17][3] ), .A1N(n6593), .Y(
        n857) );
  OAI2BB2XL U1346 ( .B0(n6881), .B1(n58), .A0N(\ram[17][4] ), .A1N(n6593), .Y(
        n858) );
  OAI2BB2XL U1347 ( .B0(n6858), .B1(n58), .A0N(\ram[17][5] ), .A1N(n6593), .Y(
        n859) );
  OAI2BB2XL U1348 ( .B0(n6835), .B1(n58), .A0N(\ram[17][6] ), .A1N(n6593), .Y(
        n860) );
  OAI2BB2XL U1349 ( .B0(n6812), .B1(n58), .A0N(\ram[17][7] ), .A1N(n6593), .Y(
        n861) );
  OAI2BB2XL U1350 ( .B0(n6789), .B1(n58), .A0N(\ram[17][8] ), .A1N(n6593), .Y(
        n862) );
  OAI2BB2XL U1351 ( .B0(n6766), .B1(n58), .A0N(\ram[17][9] ), .A1N(n6593), .Y(
        n863) );
  OAI2BB2XL U1352 ( .B0(n6743), .B1(n58), .A0N(\ram[17][10] ), .A1N(n6593), 
        .Y(n864) );
  OAI2BB2XL U1353 ( .B0(n6720), .B1(n58), .A0N(\ram[17][11] ), .A1N(n6593), 
        .Y(n865) );
  OAI2BB2XL U1354 ( .B0(n6697), .B1(n58), .A0N(\ram[17][12] ), .A1N(n6593), 
        .Y(n866) );
  OAI2BB2XL U1355 ( .B0(n6674), .B1(n58), .A0N(\ram[17][13] ), .A1N(n6593), 
        .Y(n867) );
  OAI2BB2XL U1356 ( .B0(n6651), .B1(n58), .A0N(\ram[17][14] ), .A1N(n6593), 
        .Y(n868) );
  OAI2BB2XL U1357 ( .B0(n6628), .B1(n58), .A0N(\ram[17][15] ), .A1N(n6593), 
        .Y(n869) );
  OAI2BB2XL U1358 ( .B0(n6967), .B1(n59), .A0N(\ram[18][0] ), .A1N(n6592), .Y(
        n870) );
  OAI2BB2XL U1359 ( .B0(n6944), .B1(n59), .A0N(\ram[18][1] ), .A1N(n6592), .Y(
        n871) );
  OAI2BB2XL U1360 ( .B0(n6921), .B1(n59), .A0N(\ram[18][2] ), .A1N(n6592), .Y(
        n872) );
  OAI2BB2XL U1361 ( .B0(n6898), .B1(n59), .A0N(\ram[18][3] ), .A1N(n6592), .Y(
        n873) );
  OAI2BB2XL U1362 ( .B0(n6881), .B1(n59), .A0N(\ram[18][4] ), .A1N(n6592), .Y(
        n874) );
  OAI2BB2XL U1363 ( .B0(n6858), .B1(n59), .A0N(\ram[18][5] ), .A1N(n6592), .Y(
        n875) );
  OAI2BB2XL U1364 ( .B0(n6835), .B1(n59), .A0N(\ram[18][6] ), .A1N(n6592), .Y(
        n876) );
  OAI2BB2XL U1365 ( .B0(n6812), .B1(n59), .A0N(\ram[18][7] ), .A1N(n6592), .Y(
        n877) );
  OAI2BB2XL U1366 ( .B0(n6789), .B1(n59), .A0N(\ram[18][8] ), .A1N(n6592), .Y(
        n878) );
  OAI2BB2XL U1367 ( .B0(n6766), .B1(n59), .A0N(\ram[18][9] ), .A1N(n6592), .Y(
        n879) );
  OAI2BB2XL U1368 ( .B0(n6743), .B1(n59), .A0N(\ram[18][10] ), .A1N(n6592), 
        .Y(n880) );
  OAI2BB2XL U1369 ( .B0(n6720), .B1(n59), .A0N(\ram[18][11] ), .A1N(n6592), 
        .Y(n881) );
  OAI2BB2XL U1370 ( .B0(n6697), .B1(n59), .A0N(\ram[18][12] ), .A1N(n6592), 
        .Y(n882) );
  OAI2BB2XL U1371 ( .B0(n6674), .B1(n59), .A0N(\ram[18][13] ), .A1N(n6592), 
        .Y(n883) );
  OAI2BB2XL U1372 ( .B0(n6651), .B1(n59), .A0N(\ram[18][14] ), .A1N(n6592), 
        .Y(n884) );
  OAI2BB2XL U1373 ( .B0(n6628), .B1(n59), .A0N(\ram[18][15] ), .A1N(n6592), 
        .Y(n885) );
  OAI2BB2XL U1374 ( .B0(n6966), .B1(n61), .A0N(\ram[19][0] ), .A1N(n6591), .Y(
        n886) );
  OAI2BB2XL U1375 ( .B0(n6943), .B1(n61), .A0N(\ram[19][1] ), .A1N(n6591), .Y(
        n887) );
  OAI2BB2XL U1376 ( .B0(n6920), .B1(n61), .A0N(\ram[19][2] ), .A1N(n6591), .Y(
        n888) );
  OAI2BB2XL U1377 ( .B0(n6897), .B1(n61), .A0N(\ram[19][3] ), .A1N(n6591), .Y(
        n889) );
  OAI2BB2XL U1378 ( .B0(n6881), .B1(n61), .A0N(\ram[19][4] ), .A1N(n6591), .Y(
        n890) );
  OAI2BB2XL U1379 ( .B0(n6858), .B1(n61), .A0N(\ram[19][5] ), .A1N(n6591), .Y(
        n891) );
  OAI2BB2XL U1380 ( .B0(n6835), .B1(n61), .A0N(\ram[19][6] ), .A1N(n6591), .Y(
        n892) );
  OAI2BB2XL U1381 ( .B0(n6812), .B1(n61), .A0N(\ram[19][7] ), .A1N(n6591), .Y(
        n893) );
  OAI2BB2XL U1382 ( .B0(n6789), .B1(n61), .A0N(\ram[19][8] ), .A1N(n6591), .Y(
        n894) );
  OAI2BB2XL U1383 ( .B0(n6766), .B1(n61), .A0N(\ram[19][9] ), .A1N(n6591), .Y(
        n895) );
  OAI2BB2XL U1384 ( .B0(n6743), .B1(n61), .A0N(\ram[19][10] ), .A1N(n6591), 
        .Y(n896) );
  OAI2BB2XL U1385 ( .B0(n6720), .B1(n61), .A0N(\ram[19][11] ), .A1N(n6591), 
        .Y(n897) );
  OAI2BB2XL U1386 ( .B0(n6697), .B1(n61), .A0N(\ram[19][12] ), .A1N(n6591), 
        .Y(n898) );
  OAI2BB2XL U1387 ( .B0(n6674), .B1(n61), .A0N(\ram[19][13] ), .A1N(n6591), 
        .Y(n899) );
  OAI2BB2XL U1388 ( .B0(n6651), .B1(n61), .A0N(\ram[19][14] ), .A1N(n6591), 
        .Y(n900) );
  OAI2BB2XL U1389 ( .B0(n6628), .B1(n61), .A0N(\ram[19][15] ), .A1N(n6591), 
        .Y(n901) );
  OAI2BB2XL U1390 ( .B0(n6965), .B1(n62), .A0N(\ram[20][0] ), .A1N(n6590), .Y(
        n902) );
  OAI2BB2XL U1391 ( .B0(n6942), .B1(n62), .A0N(\ram[20][1] ), .A1N(n6590), .Y(
        n903) );
  OAI2BB2XL U1392 ( .B0(n6919), .B1(n62), .A0N(\ram[20][2] ), .A1N(n6590), .Y(
        n904) );
  OAI2BB2XL U1393 ( .B0(n6896), .B1(n62), .A0N(\ram[20][3] ), .A1N(n6590), .Y(
        n905) );
  OAI2BB2XL U1394 ( .B0(n6881), .B1(n62), .A0N(\ram[20][4] ), .A1N(n6590), .Y(
        n906) );
  OAI2BB2XL U1395 ( .B0(n6858), .B1(n62), .A0N(\ram[20][5] ), .A1N(n6590), .Y(
        n907) );
  OAI2BB2XL U1396 ( .B0(n6835), .B1(n62), .A0N(\ram[20][6] ), .A1N(n6590), .Y(
        n908) );
  OAI2BB2XL U1397 ( .B0(n6812), .B1(n62), .A0N(\ram[20][7] ), .A1N(n6590), .Y(
        n909) );
  OAI2BB2XL U1398 ( .B0(n6789), .B1(n62), .A0N(\ram[20][8] ), .A1N(n6590), .Y(
        n910) );
  OAI2BB2XL U1399 ( .B0(n6766), .B1(n62), .A0N(\ram[20][9] ), .A1N(n6590), .Y(
        n911) );
  OAI2BB2XL U1400 ( .B0(n6743), .B1(n62), .A0N(\ram[20][10] ), .A1N(n6590), 
        .Y(n912) );
  OAI2BB2XL U1401 ( .B0(n6720), .B1(n62), .A0N(\ram[20][11] ), .A1N(n6590), 
        .Y(n913) );
  OAI2BB2XL U1402 ( .B0(n6697), .B1(n62), .A0N(\ram[20][12] ), .A1N(n6590), 
        .Y(n914) );
  OAI2BB2XL U1403 ( .B0(n6674), .B1(n62), .A0N(\ram[20][13] ), .A1N(n6590), 
        .Y(n915) );
  OAI2BB2XL U1404 ( .B0(n6651), .B1(n62), .A0N(\ram[20][14] ), .A1N(n6590), 
        .Y(n916) );
  OAI2BB2XL U1405 ( .B0(n6628), .B1(n62), .A0N(\ram[20][15] ), .A1N(n6590), 
        .Y(n917) );
  OAI2BB2XL U1406 ( .B0(n6964), .B1(n64), .A0N(\ram[21][0] ), .A1N(n6589), .Y(
        n918) );
  OAI2BB2XL U1407 ( .B0(n6941), .B1(n64), .A0N(\ram[21][1] ), .A1N(n6589), .Y(
        n919) );
  OAI2BB2XL U1408 ( .B0(n6918), .B1(n64), .A0N(\ram[21][2] ), .A1N(n6589), .Y(
        n920) );
  OAI2BB2XL U1409 ( .B0(n6895), .B1(n64), .A0N(\ram[21][3] ), .A1N(n6589), .Y(
        n921) );
  OAI2BB2XL U1410 ( .B0(n6881), .B1(n64), .A0N(\ram[21][4] ), .A1N(n6589), .Y(
        n922) );
  OAI2BB2XL U1411 ( .B0(n6858), .B1(n64), .A0N(\ram[21][5] ), .A1N(n6589), .Y(
        n923) );
  OAI2BB2XL U1412 ( .B0(n6835), .B1(n64), .A0N(\ram[21][6] ), .A1N(n6589), .Y(
        n924) );
  OAI2BB2XL U1413 ( .B0(n6812), .B1(n64), .A0N(\ram[21][7] ), .A1N(n6589), .Y(
        n925) );
  OAI2BB2XL U1414 ( .B0(n6789), .B1(n64), .A0N(\ram[21][8] ), .A1N(n6589), .Y(
        n926) );
  OAI2BB2XL U1415 ( .B0(n6766), .B1(n64), .A0N(\ram[21][9] ), .A1N(n6589), .Y(
        n927) );
  OAI2BB2XL U1416 ( .B0(n6743), .B1(n64), .A0N(\ram[21][10] ), .A1N(n6589), 
        .Y(n928) );
  OAI2BB2XL U1417 ( .B0(n6720), .B1(n64), .A0N(\ram[21][11] ), .A1N(n6589), 
        .Y(n929) );
  OAI2BB2XL U1418 ( .B0(n6697), .B1(n64), .A0N(\ram[21][12] ), .A1N(n6589), 
        .Y(n930) );
  OAI2BB2XL U1419 ( .B0(n6674), .B1(n64), .A0N(\ram[21][13] ), .A1N(n6589), 
        .Y(n931) );
  OAI2BB2XL U1420 ( .B0(n6651), .B1(n64), .A0N(\ram[21][14] ), .A1N(n6589), 
        .Y(n932) );
  OAI2BB2XL U1421 ( .B0(n6628), .B1(n64), .A0N(\ram[21][15] ), .A1N(n6589), 
        .Y(n933) );
  OAI2BB2XL U1422 ( .B0(n6963), .B1(n65), .A0N(\ram[22][0] ), .A1N(n6588), .Y(
        n934) );
  OAI2BB2XL U1423 ( .B0(n6940), .B1(n65), .A0N(\ram[22][1] ), .A1N(n6588), .Y(
        n935) );
  OAI2BB2XL U1424 ( .B0(n6917), .B1(n65), .A0N(\ram[22][2] ), .A1N(n6588), .Y(
        n936) );
  OAI2BB2XL U1425 ( .B0(n6894), .B1(n65), .A0N(\ram[22][3] ), .A1N(n6588), .Y(
        n937) );
  OAI2BB2XL U1426 ( .B0(n6881), .B1(n65), .A0N(\ram[22][4] ), .A1N(n6588), .Y(
        n938) );
  OAI2BB2XL U1427 ( .B0(n6858), .B1(n65), .A0N(\ram[22][5] ), .A1N(n6588), .Y(
        n939) );
  OAI2BB2XL U1428 ( .B0(n6835), .B1(n65), .A0N(\ram[22][6] ), .A1N(n6588), .Y(
        n940) );
  OAI2BB2XL U1429 ( .B0(n6812), .B1(n65), .A0N(\ram[22][7] ), .A1N(n6588), .Y(
        n941) );
  OAI2BB2XL U1430 ( .B0(n6789), .B1(n65), .A0N(\ram[22][8] ), .A1N(n6588), .Y(
        n942) );
  OAI2BB2XL U1431 ( .B0(n6766), .B1(n65), .A0N(\ram[22][9] ), .A1N(n6588), .Y(
        n943) );
  OAI2BB2XL U1432 ( .B0(n6743), .B1(n65), .A0N(\ram[22][10] ), .A1N(n6588), 
        .Y(n944) );
  OAI2BB2XL U1433 ( .B0(n6720), .B1(n65), .A0N(\ram[22][11] ), .A1N(n6588), 
        .Y(n945) );
  OAI2BB2XL U1434 ( .B0(n6697), .B1(n65), .A0N(\ram[22][12] ), .A1N(n6588), 
        .Y(n946) );
  OAI2BB2XL U1435 ( .B0(n6674), .B1(n65), .A0N(\ram[22][13] ), .A1N(n6588), 
        .Y(n947) );
  OAI2BB2XL U1436 ( .B0(n6651), .B1(n65), .A0N(\ram[22][14] ), .A1N(n6588), 
        .Y(n948) );
  OAI2BB2XL U1437 ( .B0(n6628), .B1(n65), .A0N(\ram[22][15] ), .A1N(n6588), 
        .Y(n949) );
  OAI2BB2XL U1438 ( .B0(n6957), .B1(n67), .A0N(\ram[23][0] ), .A1N(n6587), .Y(
        n950) );
  OAI2BB2XL U1439 ( .B0(n6934), .B1(n67), .A0N(\ram[23][1] ), .A1N(n6587), .Y(
        n951) );
  OAI2BB2XL U1440 ( .B0(n6911), .B1(n67), .A0N(\ram[23][2] ), .A1N(n6587), .Y(
        n952) );
  OAI2BB2XL U1441 ( .B0(n6888), .B1(n67), .A0N(\ram[23][3] ), .A1N(n6587), .Y(
        n953) );
  OAI2BB2XL U1442 ( .B0(n6881), .B1(n67), .A0N(\ram[23][4] ), .A1N(n6587), .Y(
        n954) );
  OAI2BB2XL U1443 ( .B0(n6858), .B1(n67), .A0N(\ram[23][5] ), .A1N(n6587), .Y(
        n955) );
  OAI2BB2XL U1444 ( .B0(n6835), .B1(n67), .A0N(\ram[23][6] ), .A1N(n6587), .Y(
        n956) );
  OAI2BB2XL U1445 ( .B0(n6812), .B1(n67), .A0N(\ram[23][7] ), .A1N(n6587), .Y(
        n957) );
  OAI2BB2XL U1446 ( .B0(n6789), .B1(n67), .A0N(\ram[23][8] ), .A1N(n6587), .Y(
        n958) );
  OAI2BB2XL U1447 ( .B0(n6766), .B1(n67), .A0N(\ram[23][9] ), .A1N(n6587), .Y(
        n959) );
  OAI2BB2XL U1448 ( .B0(n6743), .B1(n67), .A0N(\ram[23][10] ), .A1N(n6587), 
        .Y(n960) );
  OAI2BB2XL U1449 ( .B0(n6720), .B1(n67), .A0N(\ram[23][11] ), .A1N(n6587), 
        .Y(n961) );
  OAI2BB2XL U1450 ( .B0(n6697), .B1(n67), .A0N(\ram[23][12] ), .A1N(n6587), 
        .Y(n962) );
  OAI2BB2XL U1451 ( .B0(n6674), .B1(n67), .A0N(\ram[23][13] ), .A1N(n6587), 
        .Y(n963) );
  OAI2BB2XL U1452 ( .B0(n6651), .B1(n67), .A0N(\ram[23][14] ), .A1N(n6587), 
        .Y(n964) );
  OAI2BB2XL U1453 ( .B0(n6628), .B1(n67), .A0N(\ram[23][15] ), .A1N(n6587), 
        .Y(n965) );
  OAI2BB2XL U1454 ( .B0(n6957), .B1(n68), .A0N(\ram[24][0] ), .A1N(n6586), .Y(
        n966) );
  OAI2BB2XL U1455 ( .B0(n6934), .B1(n68), .A0N(\ram[24][1] ), .A1N(n6586), .Y(
        n967) );
  OAI2BB2XL U1456 ( .B0(n6911), .B1(n68), .A0N(\ram[24][2] ), .A1N(n6586), .Y(
        n968) );
  OAI2BB2XL U1457 ( .B0(n6888), .B1(n68), .A0N(\ram[24][3] ), .A1N(n6586), .Y(
        n969) );
  OAI2BB2XL U1458 ( .B0(n6881), .B1(n68), .A0N(\ram[24][4] ), .A1N(n6586), .Y(
        n970) );
  OAI2BB2XL U1459 ( .B0(n6858), .B1(n68), .A0N(\ram[24][5] ), .A1N(n6586), .Y(
        n971) );
  OAI2BB2XL U1460 ( .B0(n6835), .B1(n68), .A0N(\ram[24][6] ), .A1N(n6586), .Y(
        n972) );
  OAI2BB2XL U1461 ( .B0(n6812), .B1(n68), .A0N(\ram[24][7] ), .A1N(n6586), .Y(
        n973) );
  OAI2BB2XL U1462 ( .B0(n6789), .B1(n68), .A0N(\ram[24][8] ), .A1N(n6586), .Y(
        n974) );
  OAI2BB2XL U1463 ( .B0(n6766), .B1(n68), .A0N(\ram[24][9] ), .A1N(n6586), .Y(
        n975) );
  OAI2BB2XL U1464 ( .B0(n6743), .B1(n68), .A0N(\ram[24][10] ), .A1N(n6586), 
        .Y(n976) );
  OAI2BB2XL U1465 ( .B0(n6720), .B1(n68), .A0N(\ram[24][11] ), .A1N(n6586), 
        .Y(n977) );
  OAI2BB2XL U1466 ( .B0(n6697), .B1(n68), .A0N(\ram[24][12] ), .A1N(n6586), 
        .Y(n978) );
  OAI2BB2XL U1467 ( .B0(n6674), .B1(n68), .A0N(\ram[24][13] ), .A1N(n6586), 
        .Y(n979) );
  OAI2BB2XL U1468 ( .B0(n6651), .B1(n68), .A0N(\ram[24][14] ), .A1N(n6586), 
        .Y(n980) );
  OAI2BB2XL U1469 ( .B0(n6628), .B1(n68), .A0N(\ram[24][15] ), .A1N(n6586), 
        .Y(n981) );
  OAI2BB2XL U1470 ( .B0(n6960), .B1(n70), .A0N(\ram[25][0] ), .A1N(n6585), .Y(
        n982) );
  OAI2BB2XL U1471 ( .B0(n6937), .B1(n70), .A0N(\ram[25][1] ), .A1N(n6585), .Y(
        n983) );
  OAI2BB2XL U1472 ( .B0(n6914), .B1(n70), .A0N(\ram[25][2] ), .A1N(n6585), .Y(
        n984) );
  OAI2BB2XL U1473 ( .B0(n6891), .B1(n70), .A0N(\ram[25][3] ), .A1N(n6585), .Y(
        n985) );
  OAI2BB2XL U1474 ( .B0(n6881), .B1(n70), .A0N(\ram[25][4] ), .A1N(n6585), .Y(
        n986) );
  OAI2BB2XL U1475 ( .B0(n6858), .B1(n70), .A0N(\ram[25][5] ), .A1N(n6585), .Y(
        n987) );
  OAI2BB2XL U1476 ( .B0(n6835), .B1(n70), .A0N(\ram[25][6] ), .A1N(n6585), .Y(
        n988) );
  OAI2BB2XL U1477 ( .B0(n6812), .B1(n70), .A0N(\ram[25][7] ), .A1N(n6585), .Y(
        n989) );
  OAI2BB2XL U1478 ( .B0(n6789), .B1(n70), .A0N(\ram[25][8] ), .A1N(n6585), .Y(
        n990) );
  OAI2BB2XL U1479 ( .B0(n6766), .B1(n70), .A0N(\ram[25][9] ), .A1N(n6585), .Y(
        n991) );
  OAI2BB2XL U1480 ( .B0(n6743), .B1(n70), .A0N(\ram[25][10] ), .A1N(n6585), 
        .Y(n992) );
  OAI2BB2XL U1481 ( .B0(n6720), .B1(n70), .A0N(\ram[25][11] ), .A1N(n6585), 
        .Y(n993) );
  OAI2BB2XL U1482 ( .B0(n6697), .B1(n70), .A0N(\ram[25][12] ), .A1N(n6585), 
        .Y(n994) );
  OAI2BB2XL U1483 ( .B0(n6674), .B1(n70), .A0N(\ram[25][13] ), .A1N(n6585), 
        .Y(n995) );
  OAI2BB2XL U1484 ( .B0(n6651), .B1(n70), .A0N(\ram[25][14] ), .A1N(n6585), 
        .Y(n996) );
  OAI2BB2XL U1485 ( .B0(n6628), .B1(n70), .A0N(\ram[25][15] ), .A1N(n6585), 
        .Y(n997) );
  OAI2BB2XL U1486 ( .B0(n6959), .B1(n73), .A0N(\ram[26][0] ), .A1N(n6584), .Y(
        n998) );
  OAI2BB2XL U1487 ( .B0(n6936), .B1(n73), .A0N(\ram[26][1] ), .A1N(n6584), .Y(
        n999) );
  OAI2BB2XL U1488 ( .B0(n6913), .B1(n73), .A0N(\ram[26][2] ), .A1N(n6584), .Y(
        n1000) );
  OAI2BB2XL U1489 ( .B0(n6890), .B1(n73), .A0N(\ram[26][3] ), .A1N(n6584), .Y(
        n1001) );
  OAI2BB2XL U1490 ( .B0(n6881), .B1(n73), .A0N(\ram[26][4] ), .A1N(n6584), .Y(
        n1002) );
  OAI2BB2XL U1491 ( .B0(n6858), .B1(n73), .A0N(\ram[26][5] ), .A1N(n6584), .Y(
        n1003) );
  OAI2BB2XL U1492 ( .B0(n6835), .B1(n73), .A0N(\ram[26][6] ), .A1N(n6584), .Y(
        n1004) );
  OAI2BB2XL U1493 ( .B0(n6812), .B1(n73), .A0N(\ram[26][7] ), .A1N(n6584), .Y(
        n1005) );
  OAI2BB2XL U1494 ( .B0(n6789), .B1(n73), .A0N(\ram[26][8] ), .A1N(n6584), .Y(
        n1006) );
  OAI2BB2XL U1495 ( .B0(n6766), .B1(n73), .A0N(\ram[26][9] ), .A1N(n6584), .Y(
        n1007) );
  OAI2BB2XL U1496 ( .B0(n6743), .B1(n73), .A0N(\ram[26][10] ), .A1N(n6584), 
        .Y(n1008) );
  OAI2BB2XL U1497 ( .B0(n6720), .B1(n73), .A0N(\ram[26][11] ), .A1N(n6584), 
        .Y(n1009) );
  OAI2BB2XL U1498 ( .B0(n6697), .B1(n73), .A0N(\ram[26][12] ), .A1N(n6584), 
        .Y(n1010) );
  OAI2BB2XL U1499 ( .B0(n6674), .B1(n73), .A0N(\ram[26][13] ), .A1N(n6584), 
        .Y(n1011) );
  OAI2BB2XL U1500 ( .B0(n6651), .B1(n73), .A0N(\ram[26][14] ), .A1N(n6584), 
        .Y(n1012) );
  OAI2BB2XL U1501 ( .B0(n6628), .B1(n73), .A0N(\ram[26][15] ), .A1N(n6584), 
        .Y(n1013) );
  OAI2BB2XL U1502 ( .B0(n6974), .B1(n75), .A0N(\ram[27][0] ), .A1N(n6583), .Y(
        n1014) );
  OAI2BB2XL U1503 ( .B0(n6951), .B1(n75), .A0N(\ram[27][1] ), .A1N(n6583), .Y(
        n1015) );
  OAI2BB2XL U1504 ( .B0(n6928), .B1(n75), .A0N(\ram[27][2] ), .A1N(n6583), .Y(
        n1016) );
  OAI2BB2XL U1505 ( .B0(n6905), .B1(n75), .A0N(\ram[27][3] ), .A1N(n6583), .Y(
        n1017) );
  OAI2BB2XL U1506 ( .B0(n6881), .B1(n75), .A0N(\ram[27][4] ), .A1N(n6583), .Y(
        n1018) );
  OAI2BB2XL U1507 ( .B0(n6858), .B1(n75), .A0N(\ram[27][5] ), .A1N(n6583), .Y(
        n1019) );
  OAI2BB2XL U1508 ( .B0(n6835), .B1(n75), .A0N(\ram[27][6] ), .A1N(n6583), .Y(
        n1020) );
  OAI2BB2XL U1509 ( .B0(n6812), .B1(n75), .A0N(\ram[27][7] ), .A1N(n6583), .Y(
        n1021) );
  OAI2BB2XL U1510 ( .B0(n6789), .B1(n75), .A0N(\ram[27][8] ), .A1N(n6583), .Y(
        n1022) );
  OAI2BB2XL U1511 ( .B0(n6766), .B1(n75), .A0N(\ram[27][9] ), .A1N(n6583), .Y(
        n1023) );
  OAI2BB2XL U1512 ( .B0(n6743), .B1(n75), .A0N(\ram[27][10] ), .A1N(n6583), 
        .Y(n1024) );
  OAI2BB2XL U1513 ( .B0(n6720), .B1(n75), .A0N(\ram[27][11] ), .A1N(n6583), 
        .Y(n1025) );
  OAI2BB2XL U1514 ( .B0(n6697), .B1(n75), .A0N(\ram[27][12] ), .A1N(n6583), 
        .Y(n1026) );
  OAI2BB2XL U1515 ( .B0(n6674), .B1(n75), .A0N(\ram[27][13] ), .A1N(n6583), 
        .Y(n1027) );
  OAI2BB2XL U1516 ( .B0(n6651), .B1(n75), .A0N(\ram[27][14] ), .A1N(n6583), 
        .Y(n1028) );
  OAI2BB2XL U1517 ( .B0(n6628), .B1(n75), .A0N(\ram[27][15] ), .A1N(n6583), 
        .Y(n1029) );
  OAI2BB2XL U1518 ( .B0(n6966), .B1(n76), .A0N(\ram[28][0] ), .A1N(n6582), .Y(
        n1030) );
  OAI2BB2XL U1519 ( .B0(n6943), .B1(n76), .A0N(\ram[28][1] ), .A1N(n6582), .Y(
        n1031) );
  OAI2BB2XL U1520 ( .B0(n6920), .B1(n76), .A0N(\ram[28][2] ), .A1N(n6582), .Y(
        n1032) );
  OAI2BB2XL U1521 ( .B0(n6897), .B1(n76), .A0N(\ram[28][3] ), .A1N(n6582), .Y(
        n1033) );
  OAI2BB2XL U1522 ( .B0(n6880), .B1(n76), .A0N(\ram[28][4] ), .A1N(n6582), .Y(
        n1034) );
  OAI2BB2XL U1523 ( .B0(n6857), .B1(n76), .A0N(\ram[28][5] ), .A1N(n6582), .Y(
        n1035) );
  OAI2BB2XL U1524 ( .B0(n6834), .B1(n76), .A0N(\ram[28][6] ), .A1N(n6582), .Y(
        n1036) );
  OAI2BB2XL U1525 ( .B0(n6811), .B1(n76), .A0N(\ram[28][7] ), .A1N(n6582), .Y(
        n1037) );
  OAI2BB2XL U1526 ( .B0(n6788), .B1(n76), .A0N(\ram[28][8] ), .A1N(n6582), .Y(
        n1038) );
  OAI2BB2XL U1527 ( .B0(n6765), .B1(n76), .A0N(\ram[28][9] ), .A1N(n6582), .Y(
        n1039) );
  OAI2BB2XL U1528 ( .B0(n6742), .B1(n76), .A0N(\ram[28][10] ), .A1N(n6582), 
        .Y(n1040) );
  OAI2BB2XL U1529 ( .B0(n6719), .B1(n76), .A0N(\ram[28][11] ), .A1N(n6582), 
        .Y(n1041) );
  OAI2BB2XL U1530 ( .B0(n6696), .B1(n76), .A0N(\ram[28][12] ), .A1N(n6582), 
        .Y(n1042) );
  OAI2BB2XL U1531 ( .B0(n6673), .B1(n76), .A0N(\ram[28][13] ), .A1N(n6582), 
        .Y(n1043) );
  OAI2BB2XL U1532 ( .B0(n6650), .B1(n76), .A0N(\ram[28][14] ), .A1N(n6582), 
        .Y(n1044) );
  OAI2BB2XL U1533 ( .B0(n6627), .B1(n76), .A0N(\ram[28][15] ), .A1N(n6582), 
        .Y(n1045) );
  OAI2BB2XL U1534 ( .B0(n6969), .B1(n541), .A0N(\ram[29][0] ), .A1N(n6581), 
        .Y(n1046) );
  OAI2BB2XL U1535 ( .B0(n6946), .B1(n541), .A0N(\ram[29][1] ), .A1N(n6581), 
        .Y(n1047) );
  OAI2BB2XL U1536 ( .B0(n6923), .B1(n541), .A0N(\ram[29][2] ), .A1N(n6581), 
        .Y(n1048) );
  OAI2BB2XL U1537 ( .B0(n6900), .B1(n541), .A0N(\ram[29][3] ), .A1N(n6581), 
        .Y(n1049) );
  OAI2BB2XL U1538 ( .B0(n6880), .B1(n541), .A0N(\ram[29][4] ), .A1N(n6581), 
        .Y(n1050) );
  OAI2BB2XL U1539 ( .B0(n6857), .B1(n541), .A0N(\ram[29][5] ), .A1N(n6581), 
        .Y(n1051) );
  OAI2BB2XL U1540 ( .B0(n6834), .B1(n541), .A0N(\ram[29][6] ), .A1N(n6581), 
        .Y(n1052) );
  OAI2BB2XL U1541 ( .B0(n6811), .B1(n541), .A0N(\ram[29][7] ), .A1N(n6581), 
        .Y(n1053) );
  OAI2BB2XL U1542 ( .B0(n6788), .B1(n541), .A0N(\ram[29][8] ), .A1N(n6581), 
        .Y(n1054) );
  OAI2BB2XL U1543 ( .B0(n6765), .B1(n541), .A0N(\ram[29][9] ), .A1N(n6581), 
        .Y(n1055) );
  OAI2BB2XL U1544 ( .B0(n6742), .B1(n541), .A0N(\ram[29][10] ), .A1N(n6581), 
        .Y(n1056) );
  OAI2BB2XL U1545 ( .B0(n6719), .B1(n541), .A0N(\ram[29][11] ), .A1N(n6581), 
        .Y(n1057) );
  OAI2BB2XL U1546 ( .B0(n6696), .B1(n541), .A0N(\ram[29][12] ), .A1N(n6581), 
        .Y(n1058) );
  OAI2BB2XL U1547 ( .B0(n6673), .B1(n541), .A0N(\ram[29][13] ), .A1N(n6581), 
        .Y(n1059) );
  OAI2BB2XL U1548 ( .B0(n6650), .B1(n541), .A0N(\ram[29][14] ), .A1N(n6581), 
        .Y(n1060) );
  OAI2BB2XL U1549 ( .B0(n6627), .B1(n541), .A0N(\ram[29][15] ), .A1N(n6581), 
        .Y(n1061) );
  OAI2BB2XL U1550 ( .B0(n6965), .B1(n543), .A0N(\ram[30][0] ), .A1N(n6580), 
        .Y(n1062) );
  OAI2BB2XL U1551 ( .B0(n6942), .B1(n543), .A0N(\ram[30][1] ), .A1N(n6580), 
        .Y(n1063) );
  OAI2BB2XL U1552 ( .B0(n6919), .B1(n543), .A0N(\ram[30][2] ), .A1N(n6580), 
        .Y(n1064) );
  OAI2BB2XL U1553 ( .B0(n6896), .B1(n543), .A0N(\ram[30][3] ), .A1N(n6580), 
        .Y(n1065) );
  OAI2BB2XL U1554 ( .B0(n6880), .B1(n543), .A0N(\ram[30][4] ), .A1N(n6580), 
        .Y(n1066) );
  OAI2BB2XL U1555 ( .B0(n6857), .B1(n543), .A0N(\ram[30][5] ), .A1N(n6580), 
        .Y(n1067) );
  OAI2BB2XL U1556 ( .B0(n6834), .B1(n543), .A0N(\ram[30][6] ), .A1N(n6580), 
        .Y(n1068) );
  OAI2BB2XL U1557 ( .B0(n6811), .B1(n543), .A0N(\ram[30][7] ), .A1N(n6580), 
        .Y(n1069) );
  OAI2BB2XL U1558 ( .B0(n6788), .B1(n543), .A0N(\ram[30][8] ), .A1N(n6580), 
        .Y(n1070) );
  OAI2BB2XL U1559 ( .B0(n6765), .B1(n543), .A0N(\ram[30][9] ), .A1N(n6580), 
        .Y(n1071) );
  OAI2BB2XL U1560 ( .B0(n6742), .B1(n543), .A0N(\ram[30][10] ), .A1N(n6580), 
        .Y(n1072) );
  OAI2BB2XL U1561 ( .B0(n6719), .B1(n543), .A0N(\ram[30][11] ), .A1N(n6580), 
        .Y(n1073) );
  OAI2BB2XL U1562 ( .B0(n6696), .B1(n543), .A0N(\ram[30][12] ), .A1N(n6580), 
        .Y(n1074) );
  OAI2BB2XL U1563 ( .B0(n6673), .B1(n543), .A0N(\ram[30][13] ), .A1N(n6580), 
        .Y(n1075) );
  OAI2BB2XL U1564 ( .B0(n6650), .B1(n543), .A0N(\ram[30][14] ), .A1N(n6580), 
        .Y(n1076) );
  OAI2BB2XL U1565 ( .B0(n6627), .B1(n543), .A0N(\ram[30][15] ), .A1N(n6580), 
        .Y(n1077) );
  OAI2BB2XL U1566 ( .B0(n6960), .B1(n546), .A0N(\ram[31][0] ), .A1N(n6579), 
        .Y(n1078) );
  OAI2BB2XL U1567 ( .B0(n6937), .B1(n546), .A0N(\ram[31][1] ), .A1N(n6579), 
        .Y(n1079) );
  OAI2BB2XL U1568 ( .B0(n6914), .B1(n546), .A0N(\ram[31][2] ), .A1N(n6579), 
        .Y(n1080) );
  OAI2BB2XL U1569 ( .B0(n6891), .B1(n546), .A0N(\ram[31][3] ), .A1N(n6579), 
        .Y(n1081) );
  OAI2BB2XL U1570 ( .B0(n6880), .B1(n546), .A0N(\ram[31][4] ), .A1N(n6579), 
        .Y(n1082) );
  OAI2BB2XL U1571 ( .B0(n6857), .B1(n546), .A0N(\ram[31][5] ), .A1N(n6579), 
        .Y(n1083) );
  OAI2BB2XL U1572 ( .B0(n6834), .B1(n546), .A0N(\ram[31][6] ), .A1N(n6579), 
        .Y(n1084) );
  OAI2BB2XL U1573 ( .B0(n6811), .B1(n546), .A0N(\ram[31][7] ), .A1N(n6579), 
        .Y(n1085) );
  OAI2BB2XL U1574 ( .B0(n6788), .B1(n546), .A0N(\ram[31][8] ), .A1N(n6579), 
        .Y(n1086) );
  OAI2BB2XL U1575 ( .B0(n6765), .B1(n546), .A0N(\ram[31][9] ), .A1N(n6579), 
        .Y(n1087) );
  OAI2BB2XL U1576 ( .B0(n6742), .B1(n546), .A0N(\ram[31][10] ), .A1N(n6579), 
        .Y(n1088) );
  OAI2BB2XL U1577 ( .B0(n6719), .B1(n546), .A0N(\ram[31][11] ), .A1N(n6579), 
        .Y(n1089) );
  OAI2BB2XL U1578 ( .B0(n6696), .B1(n546), .A0N(\ram[31][12] ), .A1N(n6579), 
        .Y(n1090) );
  OAI2BB2XL U1579 ( .B0(n6673), .B1(n546), .A0N(\ram[31][13] ), .A1N(n6579), 
        .Y(n1091) );
  OAI2BB2XL U1580 ( .B0(n6650), .B1(n546), .A0N(\ram[31][14] ), .A1N(n6579), 
        .Y(n1092) );
  OAI2BB2XL U1581 ( .B0(n6627), .B1(n546), .A0N(\ram[31][15] ), .A1N(n6579), 
        .Y(n1093) );
  OAI2BB2XL U1582 ( .B0(n6964), .B1(n78), .A0N(\ram[32][0] ), .A1N(n6578), .Y(
        n1094) );
  OAI2BB2XL U1583 ( .B0(n6941), .B1(n78), .A0N(\ram[32][1] ), .A1N(n6578), .Y(
        n1095) );
  OAI2BB2XL U1584 ( .B0(n6918), .B1(n78), .A0N(\ram[32][2] ), .A1N(n6578), .Y(
        n1096) );
  OAI2BB2XL U1585 ( .B0(n6895), .B1(n78), .A0N(\ram[32][3] ), .A1N(n6578), .Y(
        n1097) );
  OAI2BB2XL U1586 ( .B0(n6880), .B1(n78), .A0N(\ram[32][4] ), .A1N(n6578), .Y(
        n1098) );
  OAI2BB2XL U1587 ( .B0(n6857), .B1(n78), .A0N(\ram[32][5] ), .A1N(n6578), .Y(
        n1099) );
  OAI2BB2XL U1588 ( .B0(n6834), .B1(n78), .A0N(\ram[32][6] ), .A1N(n6578), .Y(
        n1100) );
  OAI2BB2XL U1589 ( .B0(n6811), .B1(n78), .A0N(\ram[32][7] ), .A1N(n6578), .Y(
        n1101) );
  OAI2BB2XL U1590 ( .B0(n6788), .B1(n78), .A0N(\ram[32][8] ), .A1N(n6578), .Y(
        n1102) );
  OAI2BB2XL U1591 ( .B0(n6765), .B1(n78), .A0N(\ram[32][9] ), .A1N(n6578), .Y(
        n1103) );
  OAI2BB2XL U1592 ( .B0(n6742), .B1(n78), .A0N(\ram[32][10] ), .A1N(n6578), 
        .Y(n1104) );
  OAI2BB2XL U1593 ( .B0(n6719), .B1(n78), .A0N(\ram[32][11] ), .A1N(n6578), 
        .Y(n1105) );
  OAI2BB2XL U1594 ( .B0(n6696), .B1(n78), .A0N(\ram[32][12] ), .A1N(n6578), 
        .Y(n1106) );
  OAI2BB2XL U1595 ( .B0(n6673), .B1(n78), .A0N(\ram[32][13] ), .A1N(n6578), 
        .Y(n1107) );
  OAI2BB2XL U1596 ( .B0(n6650), .B1(n78), .A0N(\ram[32][14] ), .A1N(n6578), 
        .Y(n1108) );
  OAI2BB2XL U1597 ( .B0(n6627), .B1(n78), .A0N(\ram[32][15] ), .A1N(n6578), 
        .Y(n1109) );
  OAI2BB2XL U1598 ( .B0(n6959), .B1(n80), .A0N(\ram[33][0] ), .A1N(n6577), .Y(
        n1110) );
  OAI2BB2XL U1599 ( .B0(n6936), .B1(n80), .A0N(\ram[33][1] ), .A1N(n6577), .Y(
        n1111) );
  OAI2BB2XL U1600 ( .B0(n6913), .B1(n80), .A0N(\ram[33][2] ), .A1N(n6577), .Y(
        n1112) );
  OAI2BB2XL U1601 ( .B0(n6890), .B1(n80), .A0N(\ram[33][3] ), .A1N(n6577), .Y(
        n1113) );
  OAI2BB2XL U1602 ( .B0(n6880), .B1(n80), .A0N(\ram[33][4] ), .A1N(n6577), .Y(
        n1114) );
  OAI2BB2XL U1603 ( .B0(n6857), .B1(n80), .A0N(\ram[33][5] ), .A1N(n6577), .Y(
        n1115) );
  OAI2BB2XL U1604 ( .B0(n6834), .B1(n80), .A0N(\ram[33][6] ), .A1N(n6577), .Y(
        n1116) );
  OAI2BB2XL U1605 ( .B0(n6811), .B1(n80), .A0N(\ram[33][7] ), .A1N(n6577), .Y(
        n1117) );
  OAI2BB2XL U1606 ( .B0(n6788), .B1(n80), .A0N(\ram[33][8] ), .A1N(n6577), .Y(
        n1118) );
  OAI2BB2XL U1607 ( .B0(n6765), .B1(n80), .A0N(\ram[33][9] ), .A1N(n6577), .Y(
        n1119) );
  OAI2BB2XL U1608 ( .B0(n6742), .B1(n80), .A0N(\ram[33][10] ), .A1N(n6577), 
        .Y(n1120) );
  OAI2BB2XL U1609 ( .B0(n6719), .B1(n80), .A0N(\ram[33][11] ), .A1N(n6577), 
        .Y(n1121) );
  OAI2BB2XL U1610 ( .B0(n6696), .B1(n80), .A0N(\ram[33][12] ), .A1N(n6577), 
        .Y(n1122) );
  OAI2BB2XL U1611 ( .B0(n6673), .B1(n80), .A0N(\ram[33][13] ), .A1N(n6577), 
        .Y(n1123) );
  OAI2BB2XL U1612 ( .B0(n6650), .B1(n80), .A0N(\ram[33][14] ), .A1N(n6577), 
        .Y(n1124) );
  OAI2BB2XL U1613 ( .B0(n6627), .B1(n80), .A0N(\ram[33][15] ), .A1N(n6577), 
        .Y(n1125) );
  OAI2BB2XL U1614 ( .B0(n6962), .B1(n82), .A0N(\ram[34][0] ), .A1N(n6576), .Y(
        n1126) );
  OAI2BB2XL U1615 ( .B0(n6939), .B1(n82), .A0N(\ram[34][1] ), .A1N(n6576), .Y(
        n1127) );
  OAI2BB2XL U1616 ( .B0(n6916), .B1(n82), .A0N(\ram[34][2] ), .A1N(n6576), .Y(
        n1128) );
  OAI2BB2XL U1617 ( .B0(n6893), .B1(n82), .A0N(\ram[34][3] ), .A1N(n6576), .Y(
        n1129) );
  OAI2BB2XL U1618 ( .B0(n6880), .B1(n82), .A0N(\ram[34][4] ), .A1N(n6576), .Y(
        n1130) );
  OAI2BB2XL U1619 ( .B0(n6857), .B1(n82), .A0N(\ram[34][5] ), .A1N(n6576), .Y(
        n1131) );
  OAI2BB2XL U1620 ( .B0(n6834), .B1(n82), .A0N(\ram[34][6] ), .A1N(n6576), .Y(
        n1132) );
  OAI2BB2XL U1621 ( .B0(n6811), .B1(n82), .A0N(\ram[34][7] ), .A1N(n6576), .Y(
        n1133) );
  OAI2BB2XL U1622 ( .B0(n6788), .B1(n82), .A0N(\ram[34][8] ), .A1N(n6576), .Y(
        n1134) );
  OAI2BB2XL U1623 ( .B0(n6765), .B1(n82), .A0N(\ram[34][9] ), .A1N(n6576), .Y(
        n1135) );
  OAI2BB2XL U1624 ( .B0(n6742), .B1(n82), .A0N(\ram[34][10] ), .A1N(n6576), 
        .Y(n1136) );
  OAI2BB2XL U1625 ( .B0(n6719), .B1(n82), .A0N(\ram[34][11] ), .A1N(n6576), 
        .Y(n1137) );
  OAI2BB2XL U1626 ( .B0(n6696), .B1(n82), .A0N(\ram[34][12] ), .A1N(n6576), 
        .Y(n1138) );
  OAI2BB2XL U1627 ( .B0(n6673), .B1(n82), .A0N(\ram[34][13] ), .A1N(n6576), 
        .Y(n1139) );
  OAI2BB2XL U1628 ( .B0(n6650), .B1(n82), .A0N(\ram[34][14] ), .A1N(n6576), 
        .Y(n1140) );
  OAI2BB2XL U1629 ( .B0(n6627), .B1(n82), .A0N(\ram[34][15] ), .A1N(n6576), 
        .Y(n1141) );
  OAI2BB2XL U1630 ( .B0(n6963), .B1(n84), .A0N(\ram[35][0] ), .A1N(n6575), .Y(
        n1142) );
  OAI2BB2XL U1631 ( .B0(n6940), .B1(n84), .A0N(\ram[35][1] ), .A1N(n6575), .Y(
        n1143) );
  OAI2BB2XL U1632 ( .B0(n6917), .B1(n84), .A0N(\ram[35][2] ), .A1N(n6575), .Y(
        n1144) );
  OAI2BB2XL U1633 ( .B0(n6894), .B1(n84), .A0N(\ram[35][3] ), .A1N(n6575), .Y(
        n1145) );
  OAI2BB2XL U1634 ( .B0(n6880), .B1(n84), .A0N(\ram[35][4] ), .A1N(n6575), .Y(
        n1146) );
  OAI2BB2XL U1635 ( .B0(n6857), .B1(n84), .A0N(\ram[35][5] ), .A1N(n6575), .Y(
        n1147) );
  OAI2BB2XL U1636 ( .B0(n6834), .B1(n84), .A0N(\ram[35][6] ), .A1N(n6575), .Y(
        n1148) );
  OAI2BB2XL U1637 ( .B0(n6811), .B1(n84), .A0N(\ram[35][7] ), .A1N(n6575), .Y(
        n1149) );
  OAI2BB2XL U1638 ( .B0(n6788), .B1(n84), .A0N(\ram[35][8] ), .A1N(n6575), .Y(
        n1150) );
  OAI2BB2XL U1639 ( .B0(n6765), .B1(n84), .A0N(\ram[35][9] ), .A1N(n6575), .Y(
        n1151) );
  OAI2BB2XL U1640 ( .B0(n6742), .B1(n84), .A0N(\ram[35][10] ), .A1N(n6575), 
        .Y(n1152) );
  OAI2BB2XL U1641 ( .B0(n6719), .B1(n84), .A0N(\ram[35][11] ), .A1N(n6575), 
        .Y(n1153) );
  OAI2BB2XL U1642 ( .B0(n6696), .B1(n84), .A0N(\ram[35][12] ), .A1N(n6575), 
        .Y(n1154) );
  OAI2BB2XL U1643 ( .B0(n6673), .B1(n84), .A0N(\ram[35][13] ), .A1N(n6575), 
        .Y(n1155) );
  OAI2BB2XL U1644 ( .B0(n6650), .B1(n84), .A0N(\ram[35][14] ), .A1N(n6575), 
        .Y(n1156) );
  OAI2BB2XL U1645 ( .B0(n6627), .B1(n84), .A0N(\ram[35][15] ), .A1N(n6575), 
        .Y(n1157) );
  OAI2BB2XL U1646 ( .B0(n6974), .B1(n86), .A0N(\ram[36][0] ), .A1N(n6574), .Y(
        n1158) );
  OAI2BB2XL U1647 ( .B0(n6951), .B1(n86), .A0N(\ram[36][1] ), .A1N(n6574), .Y(
        n1159) );
  OAI2BB2XL U1648 ( .B0(n6928), .B1(n86), .A0N(\ram[36][2] ), .A1N(n6574), .Y(
        n1160) );
  OAI2BB2XL U1649 ( .B0(n6905), .B1(n86), .A0N(\ram[36][3] ), .A1N(n6574), .Y(
        n1161) );
  OAI2BB2XL U1650 ( .B0(n6880), .B1(n86), .A0N(\ram[36][4] ), .A1N(n6574), .Y(
        n1162) );
  OAI2BB2XL U1651 ( .B0(n6857), .B1(n86), .A0N(\ram[36][5] ), .A1N(n6574), .Y(
        n1163) );
  OAI2BB2XL U1652 ( .B0(n6834), .B1(n86), .A0N(\ram[36][6] ), .A1N(n6574), .Y(
        n1164) );
  OAI2BB2XL U1653 ( .B0(n6811), .B1(n86), .A0N(\ram[36][7] ), .A1N(n6574), .Y(
        n1165) );
  OAI2BB2XL U1654 ( .B0(n6788), .B1(n86), .A0N(\ram[36][8] ), .A1N(n6574), .Y(
        n1166) );
  OAI2BB2XL U1655 ( .B0(n6765), .B1(n86), .A0N(\ram[36][9] ), .A1N(n6574), .Y(
        n1167) );
  OAI2BB2XL U1656 ( .B0(n6742), .B1(n86), .A0N(\ram[36][10] ), .A1N(n6574), 
        .Y(n1168) );
  OAI2BB2XL U1657 ( .B0(n6719), .B1(n86), .A0N(\ram[36][11] ), .A1N(n6574), 
        .Y(n1169) );
  OAI2BB2XL U1658 ( .B0(n6696), .B1(n86), .A0N(\ram[36][12] ), .A1N(n6574), 
        .Y(n1170) );
  OAI2BB2XL U1659 ( .B0(n6673), .B1(n86), .A0N(\ram[36][13] ), .A1N(n6574), 
        .Y(n1171) );
  OAI2BB2XL U1660 ( .B0(n6650), .B1(n86), .A0N(\ram[36][14] ), .A1N(n6574), 
        .Y(n1172) );
  OAI2BB2XL U1661 ( .B0(n6627), .B1(n86), .A0N(\ram[36][15] ), .A1N(n6574), 
        .Y(n1173) );
  OAI2BB2XL U1662 ( .B0(n6973), .B1(n88), .A0N(\ram[37][0] ), .A1N(n6573), .Y(
        n1174) );
  OAI2BB2XL U1663 ( .B0(n6950), .B1(n88), .A0N(\ram[37][1] ), .A1N(n6573), .Y(
        n1175) );
  OAI2BB2XL U1664 ( .B0(n6927), .B1(n88), .A0N(\ram[37][2] ), .A1N(n6573), .Y(
        n1176) );
  OAI2BB2XL U1665 ( .B0(n6904), .B1(n88), .A0N(\ram[37][3] ), .A1N(n6573), .Y(
        n1177) );
  OAI2BB2XL U1666 ( .B0(n6880), .B1(n88), .A0N(\ram[37][4] ), .A1N(n6573), .Y(
        n1178) );
  OAI2BB2XL U1667 ( .B0(n6857), .B1(n88), .A0N(\ram[37][5] ), .A1N(n6573), .Y(
        n1179) );
  OAI2BB2XL U1668 ( .B0(n6834), .B1(n88), .A0N(\ram[37][6] ), .A1N(n6573), .Y(
        n1180) );
  OAI2BB2XL U1669 ( .B0(n6811), .B1(n88), .A0N(\ram[37][7] ), .A1N(n6573), .Y(
        n1181) );
  OAI2BB2XL U1670 ( .B0(n6788), .B1(n88), .A0N(\ram[37][8] ), .A1N(n6573), .Y(
        n1182) );
  OAI2BB2XL U1671 ( .B0(n6765), .B1(n88), .A0N(\ram[37][9] ), .A1N(n6573), .Y(
        n1183) );
  OAI2BB2XL U1672 ( .B0(n6742), .B1(n88), .A0N(\ram[37][10] ), .A1N(n6573), 
        .Y(n1184) );
  OAI2BB2XL U1673 ( .B0(n6719), .B1(n88), .A0N(\ram[37][11] ), .A1N(n6573), 
        .Y(n1185) );
  OAI2BB2XL U1674 ( .B0(n6696), .B1(n88), .A0N(\ram[37][12] ), .A1N(n6573), 
        .Y(n1186) );
  OAI2BB2XL U1675 ( .B0(n6673), .B1(n88), .A0N(\ram[37][13] ), .A1N(n6573), 
        .Y(n1187) );
  OAI2BB2XL U1676 ( .B0(n6650), .B1(n88), .A0N(\ram[37][14] ), .A1N(n6573), 
        .Y(n1188) );
  OAI2BB2XL U1677 ( .B0(n6627), .B1(n88), .A0N(\ram[37][15] ), .A1N(n6573), 
        .Y(n1189) );
  OAI2BB2XL U1678 ( .B0(n6962), .B1(n90), .A0N(\ram[38][0] ), .A1N(n6572), .Y(
        n1190) );
  OAI2BB2XL U1679 ( .B0(n6939), .B1(n90), .A0N(\ram[38][1] ), .A1N(n6572), .Y(
        n1191) );
  OAI2BB2XL U1680 ( .B0(n6916), .B1(n90), .A0N(\ram[38][2] ), .A1N(n6572), .Y(
        n1192) );
  OAI2BB2XL U1681 ( .B0(n6893), .B1(n90), .A0N(\ram[38][3] ), .A1N(n6572), .Y(
        n1193) );
  OAI2BB2XL U1682 ( .B0(n6880), .B1(n90), .A0N(\ram[38][4] ), .A1N(n6572), .Y(
        n1194) );
  OAI2BB2XL U1683 ( .B0(n6857), .B1(n90), .A0N(\ram[38][5] ), .A1N(n6572), .Y(
        n1195) );
  OAI2BB2XL U1684 ( .B0(n6834), .B1(n90), .A0N(\ram[38][6] ), .A1N(n6572), .Y(
        n1196) );
  OAI2BB2XL U1685 ( .B0(n6811), .B1(n90), .A0N(\ram[38][7] ), .A1N(n6572), .Y(
        n1197) );
  OAI2BB2XL U1686 ( .B0(n6788), .B1(n90), .A0N(\ram[38][8] ), .A1N(n6572), .Y(
        n1198) );
  OAI2BB2XL U1687 ( .B0(n6765), .B1(n90), .A0N(\ram[38][9] ), .A1N(n6572), .Y(
        n1199) );
  OAI2BB2XL U1688 ( .B0(n6742), .B1(n90), .A0N(\ram[38][10] ), .A1N(n6572), 
        .Y(n1200) );
  OAI2BB2XL U1689 ( .B0(n6719), .B1(n90), .A0N(\ram[38][11] ), .A1N(n6572), 
        .Y(n1201) );
  OAI2BB2XL U1690 ( .B0(n6696), .B1(n90), .A0N(\ram[38][12] ), .A1N(n6572), 
        .Y(n1202) );
  OAI2BB2XL U1691 ( .B0(n6673), .B1(n90), .A0N(\ram[38][13] ), .A1N(n6572), 
        .Y(n1203) );
  OAI2BB2XL U1692 ( .B0(n6650), .B1(n90), .A0N(\ram[38][14] ), .A1N(n6572), 
        .Y(n1204) );
  OAI2BB2XL U1693 ( .B0(n6627), .B1(n90), .A0N(\ram[38][15] ), .A1N(n6572), 
        .Y(n1205) );
  OAI2BB2XL U1694 ( .B0(n6973), .B1(n92), .A0N(\ram[39][0] ), .A1N(n6571), .Y(
        n1206) );
  OAI2BB2XL U1695 ( .B0(n6950), .B1(n92), .A0N(\ram[39][1] ), .A1N(n6571), .Y(
        n1207) );
  OAI2BB2XL U1696 ( .B0(n6927), .B1(n92), .A0N(\ram[39][2] ), .A1N(n6571), .Y(
        n1208) );
  OAI2BB2XL U1697 ( .B0(n6904), .B1(n92), .A0N(\ram[39][3] ), .A1N(n6571), .Y(
        n1209) );
  OAI2BB2XL U1698 ( .B0(n6880), .B1(n92), .A0N(\ram[39][4] ), .A1N(n6571), .Y(
        n1210) );
  OAI2BB2XL U1699 ( .B0(n6857), .B1(n92), .A0N(\ram[39][5] ), .A1N(n6571), .Y(
        n1211) );
  OAI2BB2XL U1700 ( .B0(n6834), .B1(n92), .A0N(\ram[39][6] ), .A1N(n6571), .Y(
        n1212) );
  OAI2BB2XL U1701 ( .B0(n6811), .B1(n92), .A0N(\ram[39][7] ), .A1N(n6571), .Y(
        n1213) );
  OAI2BB2XL U1702 ( .B0(n6788), .B1(n92), .A0N(\ram[39][8] ), .A1N(n6571), .Y(
        n1214) );
  OAI2BB2XL U1703 ( .B0(n6765), .B1(n92), .A0N(\ram[39][9] ), .A1N(n6571), .Y(
        n1215) );
  OAI2BB2XL U1704 ( .B0(n6742), .B1(n92), .A0N(\ram[39][10] ), .A1N(n6571), 
        .Y(n1216) );
  OAI2BB2XL U1705 ( .B0(n6719), .B1(n92), .A0N(\ram[39][11] ), .A1N(n6571), 
        .Y(n1217) );
  OAI2BB2XL U1706 ( .B0(n6696), .B1(n92), .A0N(\ram[39][12] ), .A1N(n6571), 
        .Y(n1218) );
  OAI2BB2XL U1707 ( .B0(n6673), .B1(n92), .A0N(\ram[39][13] ), .A1N(n6571), 
        .Y(n1219) );
  OAI2BB2XL U1708 ( .B0(n6650), .B1(n92), .A0N(\ram[39][14] ), .A1N(n6571), 
        .Y(n1220) );
  OAI2BB2XL U1709 ( .B0(n6627), .B1(n92), .A0N(\ram[39][15] ), .A1N(n6571), 
        .Y(n1221) );
  OAI2BB2XL U1710 ( .B0(n6968), .B1(n94), .A0N(\ram[40][0] ), .A1N(n6570), .Y(
        n1222) );
  OAI2BB2XL U1711 ( .B0(n6945), .B1(n94), .A0N(\ram[40][1] ), .A1N(n6570), .Y(
        n1223) );
  OAI2BB2XL U1712 ( .B0(n6922), .B1(n94), .A0N(\ram[40][2] ), .A1N(n6570), .Y(
        n1224) );
  OAI2BB2XL U1713 ( .B0(n6899), .B1(n94), .A0N(\ram[40][3] ), .A1N(n6570), .Y(
        n1225) );
  OAI2BB2XL U1714 ( .B0(n6879), .B1(n94), .A0N(\ram[40][4] ), .A1N(n6570), .Y(
        n1226) );
  OAI2BB2XL U1715 ( .B0(n6856), .B1(n94), .A0N(\ram[40][5] ), .A1N(n6570), .Y(
        n1227) );
  OAI2BB2XL U1716 ( .B0(n6833), .B1(n94), .A0N(\ram[40][6] ), .A1N(n6570), .Y(
        n1228) );
  OAI2BB2XL U1717 ( .B0(n6810), .B1(n94), .A0N(\ram[40][7] ), .A1N(n6570), .Y(
        n1229) );
  OAI2BB2XL U1718 ( .B0(n6787), .B1(n94), .A0N(\ram[40][8] ), .A1N(n6570), .Y(
        n1230) );
  OAI2BB2XL U1719 ( .B0(n6764), .B1(n94), .A0N(\ram[40][9] ), .A1N(n6570), .Y(
        n1231) );
  OAI2BB2XL U1720 ( .B0(n6741), .B1(n94), .A0N(\ram[40][10] ), .A1N(n6570), 
        .Y(n1232) );
  OAI2BB2XL U1721 ( .B0(n6718), .B1(n94), .A0N(\ram[40][11] ), .A1N(n6570), 
        .Y(n1233) );
  OAI2BB2XL U1722 ( .B0(n6695), .B1(n94), .A0N(\ram[40][12] ), .A1N(n6570), 
        .Y(n1234) );
  OAI2BB2XL U1723 ( .B0(n6672), .B1(n94), .A0N(\ram[40][13] ), .A1N(n6570), 
        .Y(n1235) );
  OAI2BB2XL U1724 ( .B0(n6649), .B1(n94), .A0N(\ram[40][14] ), .A1N(n6570), 
        .Y(n1236) );
  OAI2BB2XL U1725 ( .B0(n6626), .B1(n94), .A0N(\ram[40][15] ), .A1N(n6570), 
        .Y(n1237) );
  OAI2BB2XL U1726 ( .B0(n6967), .B1(n96), .A0N(\ram[41][0] ), .A1N(n6569), .Y(
        n1238) );
  OAI2BB2XL U1727 ( .B0(n6944), .B1(n96), .A0N(\ram[41][1] ), .A1N(n6569), .Y(
        n1239) );
  OAI2BB2XL U1728 ( .B0(n6921), .B1(n96), .A0N(\ram[41][2] ), .A1N(n6569), .Y(
        n1240) );
  OAI2BB2XL U1729 ( .B0(n6898), .B1(n96), .A0N(\ram[41][3] ), .A1N(n6569), .Y(
        n1241) );
  OAI2BB2XL U1730 ( .B0(n6879), .B1(n96), .A0N(\ram[41][4] ), .A1N(n6569), .Y(
        n1242) );
  OAI2BB2XL U1731 ( .B0(n6856), .B1(n96), .A0N(\ram[41][5] ), .A1N(n6569), .Y(
        n1243) );
  OAI2BB2XL U1732 ( .B0(n6833), .B1(n96), .A0N(\ram[41][6] ), .A1N(n6569), .Y(
        n1244) );
  OAI2BB2XL U1733 ( .B0(n6810), .B1(n96), .A0N(\ram[41][7] ), .A1N(n6569), .Y(
        n1245) );
  OAI2BB2XL U1734 ( .B0(n6787), .B1(n96), .A0N(\ram[41][8] ), .A1N(n6569), .Y(
        n1246) );
  OAI2BB2XL U1735 ( .B0(n6764), .B1(n96), .A0N(\ram[41][9] ), .A1N(n6569), .Y(
        n1247) );
  OAI2BB2XL U1736 ( .B0(n6741), .B1(n96), .A0N(\ram[41][10] ), .A1N(n6569), 
        .Y(n1248) );
  OAI2BB2XL U1737 ( .B0(n6718), .B1(n96), .A0N(\ram[41][11] ), .A1N(n6569), 
        .Y(n1249) );
  OAI2BB2XL U1738 ( .B0(n6695), .B1(n96), .A0N(\ram[41][12] ), .A1N(n6569), 
        .Y(n1250) );
  OAI2BB2XL U1739 ( .B0(n6672), .B1(n96), .A0N(\ram[41][13] ), .A1N(n6569), 
        .Y(n1251) );
  OAI2BB2XL U1740 ( .B0(n6649), .B1(n96), .A0N(\ram[41][14] ), .A1N(n6569), 
        .Y(n1252) );
  OAI2BB2XL U1741 ( .B0(n6626), .B1(n96), .A0N(\ram[41][15] ), .A1N(n6569), 
        .Y(n1253) );
  OAI2BB2XL U1742 ( .B0(n6966), .B1(n460), .A0N(\ram[42][0] ), .A1N(n6568), 
        .Y(n1254) );
  OAI2BB2XL U1743 ( .B0(n6943), .B1(n460), .A0N(\ram[42][1] ), .A1N(n6568), 
        .Y(n1255) );
  OAI2BB2XL U1744 ( .B0(n6920), .B1(n460), .A0N(\ram[42][2] ), .A1N(n6568), 
        .Y(n1256) );
  OAI2BB2XL U1745 ( .B0(n6897), .B1(n460), .A0N(\ram[42][3] ), .A1N(n6568), 
        .Y(n1257) );
  OAI2BB2XL U1746 ( .B0(n6879), .B1(n460), .A0N(\ram[42][4] ), .A1N(n6568), 
        .Y(n1258) );
  OAI2BB2XL U1747 ( .B0(n6856), .B1(n460), .A0N(\ram[42][5] ), .A1N(n6568), 
        .Y(n1259) );
  OAI2BB2XL U1748 ( .B0(n6833), .B1(n460), .A0N(\ram[42][6] ), .A1N(n6568), 
        .Y(n1260) );
  OAI2BB2XL U1749 ( .B0(n6810), .B1(n460), .A0N(\ram[42][7] ), .A1N(n6568), 
        .Y(n1261) );
  OAI2BB2XL U1750 ( .B0(n6787), .B1(n460), .A0N(\ram[42][8] ), .A1N(n6568), 
        .Y(n1262) );
  OAI2BB2XL U1751 ( .B0(n6764), .B1(n460), .A0N(\ram[42][9] ), .A1N(n6568), 
        .Y(n1263) );
  OAI2BB2XL U1752 ( .B0(n6741), .B1(n460), .A0N(\ram[42][10] ), .A1N(n6568), 
        .Y(n1264) );
  OAI2BB2XL U1753 ( .B0(n6718), .B1(n460), .A0N(\ram[42][11] ), .A1N(n6568), 
        .Y(n1265) );
  OAI2BB2XL U1754 ( .B0(n6695), .B1(n460), .A0N(\ram[42][12] ), .A1N(n6568), 
        .Y(n1266) );
  OAI2BB2XL U1755 ( .B0(n6672), .B1(n460), .A0N(\ram[42][13] ), .A1N(n6568), 
        .Y(n1267) );
  OAI2BB2XL U1756 ( .B0(n6649), .B1(n460), .A0N(\ram[42][14] ), .A1N(n6568), 
        .Y(n1268) );
  OAI2BB2XL U1757 ( .B0(n6626), .B1(n460), .A0N(\ram[42][15] ), .A1N(n6568), 
        .Y(n1269) );
  OAI2BB2XL U1758 ( .B0(n6965), .B1(n98), .A0N(\ram[43][0] ), .A1N(n6567), .Y(
        n1270) );
  OAI2BB2XL U1759 ( .B0(n6942), .B1(n98), .A0N(\ram[43][1] ), .A1N(n6567), .Y(
        n1271) );
  OAI2BB2XL U1760 ( .B0(n6919), .B1(n98), .A0N(\ram[43][2] ), .A1N(n6567), .Y(
        n1272) );
  OAI2BB2XL U1761 ( .B0(n6896), .B1(n98), .A0N(\ram[43][3] ), .A1N(n6567), .Y(
        n1273) );
  OAI2BB2XL U1762 ( .B0(n6879), .B1(n98), .A0N(\ram[43][4] ), .A1N(n6567), .Y(
        n1274) );
  OAI2BB2XL U1763 ( .B0(n6856), .B1(n98), .A0N(\ram[43][5] ), .A1N(n6567), .Y(
        n1275) );
  OAI2BB2XL U1764 ( .B0(n6833), .B1(n98), .A0N(\ram[43][6] ), .A1N(n6567), .Y(
        n1276) );
  OAI2BB2XL U1765 ( .B0(n6810), .B1(n98), .A0N(\ram[43][7] ), .A1N(n6567), .Y(
        n1277) );
  OAI2BB2XL U1766 ( .B0(n6787), .B1(n98), .A0N(\ram[43][8] ), .A1N(n6567), .Y(
        n1278) );
  OAI2BB2XL U1767 ( .B0(n6764), .B1(n98), .A0N(\ram[43][9] ), .A1N(n6567), .Y(
        n1279) );
  OAI2BB2XL U1768 ( .B0(n6741), .B1(n98), .A0N(\ram[43][10] ), .A1N(n6567), 
        .Y(n1280) );
  OAI2BB2XL U1769 ( .B0(n6718), .B1(n98), .A0N(\ram[43][11] ), .A1N(n6567), 
        .Y(n1281) );
  OAI2BB2XL U1770 ( .B0(n6695), .B1(n98), .A0N(\ram[43][12] ), .A1N(n6567), 
        .Y(n1282) );
  OAI2BB2XL U1771 ( .B0(n6672), .B1(n98), .A0N(\ram[43][13] ), .A1N(n6567), 
        .Y(n1283) );
  OAI2BB2XL U1772 ( .B0(n6649), .B1(n98), .A0N(\ram[43][14] ), .A1N(n6567), 
        .Y(n1284) );
  OAI2BB2XL U1773 ( .B0(n6626), .B1(n98), .A0N(\ram[43][15] ), .A1N(n6567), 
        .Y(n1285) );
  OAI2BB2XL U1774 ( .B0(n6964), .B1(n100), .A0N(\ram[44][0] ), .A1N(n6566), 
        .Y(n1286) );
  OAI2BB2XL U1775 ( .B0(n6941), .B1(n100), .A0N(\ram[44][1] ), .A1N(n6566), 
        .Y(n1287) );
  OAI2BB2XL U1776 ( .B0(n6918), .B1(n100), .A0N(\ram[44][2] ), .A1N(n6566), 
        .Y(n1288) );
  OAI2BB2XL U1777 ( .B0(n6895), .B1(n100), .A0N(\ram[44][3] ), .A1N(n6566), 
        .Y(n1289) );
  OAI2BB2XL U1778 ( .B0(n6879), .B1(n100), .A0N(\ram[44][4] ), .A1N(n6566), 
        .Y(n1290) );
  OAI2BB2XL U1779 ( .B0(n6856), .B1(n100), .A0N(\ram[44][5] ), .A1N(n6566), 
        .Y(n1291) );
  OAI2BB2XL U1780 ( .B0(n6833), .B1(n100), .A0N(\ram[44][6] ), .A1N(n6566), 
        .Y(n1292) );
  OAI2BB2XL U1781 ( .B0(n6810), .B1(n100), .A0N(\ram[44][7] ), .A1N(n6566), 
        .Y(n1293) );
  OAI2BB2XL U1782 ( .B0(n6787), .B1(n100), .A0N(\ram[44][8] ), .A1N(n6566), 
        .Y(n1294) );
  OAI2BB2XL U1783 ( .B0(n6764), .B1(n100), .A0N(\ram[44][9] ), .A1N(n6566), 
        .Y(n1295) );
  OAI2BB2XL U1784 ( .B0(n6741), .B1(n100), .A0N(\ram[44][10] ), .A1N(n6566), 
        .Y(n1296) );
  OAI2BB2XL U1785 ( .B0(n6718), .B1(n100), .A0N(\ram[44][11] ), .A1N(n6566), 
        .Y(n1297) );
  OAI2BB2XL U1786 ( .B0(n6695), .B1(n100), .A0N(\ram[44][12] ), .A1N(n6566), 
        .Y(n1298) );
  OAI2BB2XL U1787 ( .B0(n6672), .B1(n100), .A0N(\ram[44][13] ), .A1N(n6566), 
        .Y(n1299) );
  OAI2BB2XL U1788 ( .B0(n6649), .B1(n100), .A0N(\ram[44][14] ), .A1N(n6566), 
        .Y(n1300) );
  OAI2BB2XL U1789 ( .B0(n6626), .B1(n100), .A0N(\ram[44][15] ), .A1N(n6566), 
        .Y(n1301) );
  OAI2BB2XL U1790 ( .B0(n6963), .B1(n102), .A0N(\ram[45][0] ), .A1N(n6565), 
        .Y(n1302) );
  OAI2BB2XL U1791 ( .B0(n6940), .B1(n102), .A0N(\ram[45][1] ), .A1N(n6565), 
        .Y(n1303) );
  OAI2BB2XL U1792 ( .B0(n6917), .B1(n102), .A0N(\ram[45][2] ), .A1N(n6565), 
        .Y(n1304) );
  OAI2BB2XL U1793 ( .B0(n6894), .B1(n102), .A0N(\ram[45][3] ), .A1N(n6565), 
        .Y(n1305) );
  OAI2BB2XL U1794 ( .B0(n6879), .B1(n102), .A0N(\ram[45][4] ), .A1N(n6565), 
        .Y(n1306) );
  OAI2BB2XL U1795 ( .B0(n6856), .B1(n102), .A0N(\ram[45][5] ), .A1N(n6565), 
        .Y(n1307) );
  OAI2BB2XL U1796 ( .B0(n6833), .B1(n102), .A0N(\ram[45][6] ), .A1N(n6565), 
        .Y(n1308) );
  OAI2BB2XL U1797 ( .B0(n6810), .B1(n102), .A0N(\ram[45][7] ), .A1N(n6565), 
        .Y(n1309) );
  OAI2BB2XL U1798 ( .B0(n6787), .B1(n102), .A0N(\ram[45][8] ), .A1N(n6565), 
        .Y(n1310) );
  OAI2BB2XL U1799 ( .B0(n6764), .B1(n102), .A0N(\ram[45][9] ), .A1N(n6565), 
        .Y(n1311) );
  OAI2BB2XL U1800 ( .B0(n6741), .B1(n102), .A0N(\ram[45][10] ), .A1N(n6565), 
        .Y(n1312) );
  OAI2BB2XL U1801 ( .B0(n6718), .B1(n102), .A0N(\ram[45][11] ), .A1N(n6565), 
        .Y(n1313) );
  OAI2BB2XL U1802 ( .B0(n6695), .B1(n102), .A0N(\ram[45][12] ), .A1N(n6565), 
        .Y(n1314) );
  OAI2BB2XL U1803 ( .B0(n6672), .B1(n102), .A0N(\ram[45][13] ), .A1N(n6565), 
        .Y(n1315) );
  OAI2BB2XL U1804 ( .B0(n6649), .B1(n102), .A0N(\ram[45][14] ), .A1N(n6565), 
        .Y(n1316) );
  OAI2BB2XL U1805 ( .B0(n6626), .B1(n102), .A0N(\ram[45][15] ), .A1N(n6565), 
        .Y(n1317) );
  OAI2BB2XL U1806 ( .B0(n6962), .B1(n496), .A0N(\ram[46][0] ), .A1N(n6564), 
        .Y(n1318) );
  OAI2BB2XL U1807 ( .B0(n6939), .B1(n496), .A0N(\ram[46][1] ), .A1N(n6564), 
        .Y(n1319) );
  OAI2BB2XL U1808 ( .B0(n6916), .B1(n496), .A0N(\ram[46][2] ), .A1N(n6564), 
        .Y(n1320) );
  OAI2BB2XL U1809 ( .B0(n6893), .B1(n496), .A0N(\ram[46][3] ), .A1N(n6564), 
        .Y(n1321) );
  OAI2BB2XL U1810 ( .B0(n6879), .B1(n496), .A0N(\ram[46][4] ), .A1N(n6564), 
        .Y(n1322) );
  OAI2BB2XL U1811 ( .B0(n6856), .B1(n496), .A0N(\ram[46][5] ), .A1N(n6564), 
        .Y(n1323) );
  OAI2BB2XL U1812 ( .B0(n6833), .B1(n496), .A0N(\ram[46][6] ), .A1N(n6564), 
        .Y(n1324) );
  OAI2BB2XL U1813 ( .B0(n6810), .B1(n496), .A0N(\ram[46][7] ), .A1N(n6564), 
        .Y(n1325) );
  OAI2BB2XL U1814 ( .B0(n6787), .B1(n496), .A0N(\ram[46][8] ), .A1N(n6564), 
        .Y(n1326) );
  OAI2BB2XL U1815 ( .B0(n6764), .B1(n496), .A0N(\ram[46][9] ), .A1N(n6564), 
        .Y(n1327) );
  OAI2BB2XL U1816 ( .B0(n6741), .B1(n496), .A0N(\ram[46][10] ), .A1N(n6564), 
        .Y(n1328) );
  OAI2BB2XL U1817 ( .B0(n6718), .B1(n496), .A0N(\ram[46][11] ), .A1N(n6564), 
        .Y(n1329) );
  OAI2BB2XL U1818 ( .B0(n6695), .B1(n496), .A0N(\ram[46][12] ), .A1N(n6564), 
        .Y(n1330) );
  OAI2BB2XL U1819 ( .B0(n6672), .B1(n496), .A0N(\ram[46][13] ), .A1N(n6564), 
        .Y(n1331) );
  OAI2BB2XL U1820 ( .B0(n6649), .B1(n496), .A0N(\ram[46][14] ), .A1N(n6564), 
        .Y(n1332) );
  OAI2BB2XL U1821 ( .B0(n6626), .B1(n496), .A0N(\ram[46][15] ), .A1N(n6564), 
        .Y(n1333) );
  OAI2BB2XL U1822 ( .B0(n6961), .B1(n104), .A0N(\ram[47][0] ), .A1N(n6563), 
        .Y(n1334) );
  OAI2BB2XL U1823 ( .B0(n6938), .B1(n104), .A0N(\ram[47][1] ), .A1N(n6563), 
        .Y(n1335) );
  OAI2BB2XL U1824 ( .B0(n6915), .B1(n104), .A0N(\ram[47][2] ), .A1N(n6563), 
        .Y(n1336) );
  OAI2BB2XL U1825 ( .B0(n6892), .B1(n104), .A0N(\ram[47][3] ), .A1N(n6563), 
        .Y(n1337) );
  OAI2BB2XL U1826 ( .B0(n6879), .B1(n104), .A0N(\ram[47][4] ), .A1N(n6563), 
        .Y(n1338) );
  OAI2BB2XL U1827 ( .B0(n6856), .B1(n104), .A0N(\ram[47][5] ), .A1N(n6563), 
        .Y(n1339) );
  OAI2BB2XL U1828 ( .B0(n6833), .B1(n104), .A0N(\ram[47][6] ), .A1N(n6563), 
        .Y(n1340) );
  OAI2BB2XL U1829 ( .B0(n6810), .B1(n104), .A0N(\ram[47][7] ), .A1N(n6563), 
        .Y(n1341) );
  OAI2BB2XL U1830 ( .B0(n6787), .B1(n104), .A0N(\ram[47][8] ), .A1N(n6563), 
        .Y(n1342) );
  OAI2BB2XL U1831 ( .B0(n6764), .B1(n104), .A0N(\ram[47][9] ), .A1N(n6563), 
        .Y(n1343) );
  OAI2BB2XL U1832 ( .B0(n6741), .B1(n104), .A0N(\ram[47][10] ), .A1N(n6563), 
        .Y(n1344) );
  OAI2BB2XL U1833 ( .B0(n6718), .B1(n104), .A0N(\ram[47][11] ), .A1N(n6563), 
        .Y(n1345) );
  OAI2BB2XL U1834 ( .B0(n6695), .B1(n104), .A0N(\ram[47][12] ), .A1N(n6563), 
        .Y(n1346) );
  OAI2BB2XL U1835 ( .B0(n6672), .B1(n104), .A0N(\ram[47][13] ), .A1N(n6563), 
        .Y(n1347) );
  OAI2BB2XL U1836 ( .B0(n6649), .B1(n104), .A0N(\ram[47][14] ), .A1N(n6563), 
        .Y(n1348) );
  OAI2BB2XL U1837 ( .B0(n6626), .B1(n104), .A0N(\ram[47][15] ), .A1N(n6563), 
        .Y(n1349) );
  OAI2BB2XL U1838 ( .B0(n6968), .B1(n107), .A0N(\ram[48][0] ), .A1N(n6562), 
        .Y(n1350) );
  OAI2BB2XL U1839 ( .B0(n6945), .B1(n107), .A0N(\ram[48][1] ), .A1N(n6562), 
        .Y(n1351) );
  OAI2BB2XL U1840 ( .B0(n6922), .B1(n107), .A0N(\ram[48][2] ), .A1N(n6562), 
        .Y(n1352) );
  OAI2BB2XL U1841 ( .B0(n6899), .B1(n107), .A0N(\ram[48][3] ), .A1N(n6562), 
        .Y(n1353) );
  OAI2BB2XL U1842 ( .B0(n6879), .B1(n107), .A0N(\ram[48][4] ), .A1N(n6562), 
        .Y(n1354) );
  OAI2BB2XL U1843 ( .B0(n6856), .B1(n107), .A0N(\ram[48][5] ), .A1N(n6562), 
        .Y(n1355) );
  OAI2BB2XL U1844 ( .B0(n6833), .B1(n107), .A0N(\ram[48][6] ), .A1N(n6562), 
        .Y(n1356) );
  OAI2BB2XL U1845 ( .B0(n6810), .B1(n107), .A0N(\ram[48][7] ), .A1N(n6562), 
        .Y(n1357) );
  OAI2BB2XL U1846 ( .B0(n6787), .B1(n107), .A0N(\ram[48][8] ), .A1N(n6562), 
        .Y(n1358) );
  OAI2BB2XL U1847 ( .B0(n6764), .B1(n107), .A0N(\ram[48][9] ), .A1N(n6562), 
        .Y(n1359) );
  OAI2BB2XL U1848 ( .B0(n6741), .B1(n107), .A0N(\ram[48][10] ), .A1N(n6562), 
        .Y(n1360) );
  OAI2BB2XL U1849 ( .B0(n6718), .B1(n107), .A0N(\ram[48][11] ), .A1N(n6562), 
        .Y(n1361) );
  OAI2BB2XL U1850 ( .B0(n6695), .B1(n107), .A0N(\ram[48][12] ), .A1N(n6562), 
        .Y(n1362) );
  OAI2BB2XL U1851 ( .B0(n6672), .B1(n107), .A0N(\ram[48][13] ), .A1N(n6562), 
        .Y(n1363) );
  OAI2BB2XL U1852 ( .B0(n6649), .B1(n107), .A0N(\ram[48][14] ), .A1N(n6562), 
        .Y(n1364) );
  OAI2BB2XL U1853 ( .B0(n6626), .B1(n107), .A0N(\ram[48][15] ), .A1N(n6562), 
        .Y(n1365) );
  OAI2BB2XL U1854 ( .B0(n6967), .B1(n109), .A0N(\ram[49][0] ), .A1N(n6561), 
        .Y(n1366) );
  OAI2BB2XL U1855 ( .B0(n6944), .B1(n109), .A0N(\ram[49][1] ), .A1N(n6561), 
        .Y(n1367) );
  OAI2BB2XL U1856 ( .B0(n6921), .B1(n109), .A0N(\ram[49][2] ), .A1N(n6561), 
        .Y(n1368) );
  OAI2BB2XL U1857 ( .B0(n6898), .B1(n109), .A0N(\ram[49][3] ), .A1N(n6561), 
        .Y(n1369) );
  OAI2BB2XL U1858 ( .B0(n6879), .B1(n109), .A0N(\ram[49][4] ), .A1N(n6561), 
        .Y(n1370) );
  OAI2BB2XL U1859 ( .B0(n6856), .B1(n109), .A0N(\ram[49][5] ), .A1N(n6561), 
        .Y(n1371) );
  OAI2BB2XL U1860 ( .B0(n6833), .B1(n109), .A0N(\ram[49][6] ), .A1N(n6561), 
        .Y(n1372) );
  OAI2BB2XL U1861 ( .B0(n6810), .B1(n109), .A0N(\ram[49][7] ), .A1N(n6561), 
        .Y(n1373) );
  OAI2BB2XL U1862 ( .B0(n6787), .B1(n109), .A0N(\ram[49][8] ), .A1N(n6561), 
        .Y(n1374) );
  OAI2BB2XL U1863 ( .B0(n6764), .B1(n109), .A0N(\ram[49][9] ), .A1N(n6561), 
        .Y(n1375) );
  OAI2BB2XL U1864 ( .B0(n6741), .B1(n109), .A0N(\ram[49][10] ), .A1N(n6561), 
        .Y(n1376) );
  OAI2BB2XL U1865 ( .B0(n6718), .B1(n109), .A0N(\ram[49][11] ), .A1N(n6561), 
        .Y(n1377) );
  OAI2BB2XL U1866 ( .B0(n6695), .B1(n109), .A0N(\ram[49][12] ), .A1N(n6561), 
        .Y(n1378) );
  OAI2BB2XL U1867 ( .B0(n6672), .B1(n109), .A0N(\ram[49][13] ), .A1N(n6561), 
        .Y(n1379) );
  OAI2BB2XL U1868 ( .B0(n6649), .B1(n109), .A0N(\ram[49][14] ), .A1N(n6561), 
        .Y(n1380) );
  OAI2BB2XL U1869 ( .B0(n6626), .B1(n109), .A0N(\ram[49][15] ), .A1N(n6561), 
        .Y(n1381) );
  OAI2BB2XL U1870 ( .B0(n6966), .B1(n110), .A0N(\ram[50][0] ), .A1N(n6560), 
        .Y(n1382) );
  OAI2BB2XL U1871 ( .B0(n6943), .B1(n110), .A0N(\ram[50][1] ), .A1N(n6560), 
        .Y(n1383) );
  OAI2BB2XL U1872 ( .B0(n6920), .B1(n110), .A0N(\ram[50][2] ), .A1N(n6560), 
        .Y(n1384) );
  OAI2BB2XL U1873 ( .B0(n6897), .B1(n110), .A0N(\ram[50][3] ), .A1N(n6560), 
        .Y(n1385) );
  OAI2BB2XL U1874 ( .B0(n6879), .B1(n110), .A0N(\ram[50][4] ), .A1N(n6560), 
        .Y(n1386) );
  OAI2BB2XL U1875 ( .B0(n6856), .B1(n110), .A0N(\ram[50][5] ), .A1N(n6560), 
        .Y(n1387) );
  OAI2BB2XL U1876 ( .B0(n6833), .B1(n110), .A0N(\ram[50][6] ), .A1N(n6560), 
        .Y(n1388) );
  OAI2BB2XL U1877 ( .B0(n6810), .B1(n110), .A0N(\ram[50][7] ), .A1N(n6560), 
        .Y(n1389) );
  OAI2BB2XL U1878 ( .B0(n6787), .B1(n110), .A0N(\ram[50][8] ), .A1N(n6560), 
        .Y(n1390) );
  OAI2BB2XL U1879 ( .B0(n6764), .B1(n110), .A0N(\ram[50][9] ), .A1N(n6560), 
        .Y(n1391) );
  OAI2BB2XL U1880 ( .B0(n6741), .B1(n110), .A0N(\ram[50][10] ), .A1N(n6560), 
        .Y(n1392) );
  OAI2BB2XL U1881 ( .B0(n6718), .B1(n110), .A0N(\ram[50][11] ), .A1N(n6560), 
        .Y(n1393) );
  OAI2BB2XL U1882 ( .B0(n6695), .B1(n110), .A0N(\ram[50][12] ), .A1N(n6560), 
        .Y(n1394) );
  OAI2BB2XL U1883 ( .B0(n6672), .B1(n110), .A0N(\ram[50][13] ), .A1N(n6560), 
        .Y(n1395) );
  OAI2BB2XL U1884 ( .B0(n6649), .B1(n110), .A0N(\ram[50][14] ), .A1N(n6560), 
        .Y(n1396) );
  OAI2BB2XL U1885 ( .B0(n6626), .B1(n110), .A0N(\ram[50][15] ), .A1N(n6560), 
        .Y(n1397) );
  OAI2BB2XL U1886 ( .B0(n6965), .B1(n112), .A0N(\ram[51][0] ), .A1N(n6559), 
        .Y(n1398) );
  OAI2BB2XL U1887 ( .B0(n6942), .B1(n112), .A0N(\ram[51][1] ), .A1N(n6559), 
        .Y(n1399) );
  OAI2BB2XL U1888 ( .B0(n6919), .B1(n112), .A0N(\ram[51][2] ), .A1N(n6559), 
        .Y(n1400) );
  OAI2BB2XL U1889 ( .B0(n6896), .B1(n112), .A0N(\ram[51][3] ), .A1N(n6559), 
        .Y(n1401) );
  OAI2BB2XL U1890 ( .B0(n6879), .B1(n112), .A0N(\ram[51][4] ), .A1N(n6559), 
        .Y(n1402) );
  OAI2BB2XL U1891 ( .B0(n6856), .B1(n112), .A0N(\ram[51][5] ), .A1N(n6559), 
        .Y(n1403) );
  OAI2BB2XL U1892 ( .B0(n6833), .B1(n112), .A0N(\ram[51][6] ), .A1N(n6559), 
        .Y(n1404) );
  OAI2BB2XL U1893 ( .B0(n6810), .B1(n112), .A0N(\ram[51][7] ), .A1N(n6559), 
        .Y(n1405) );
  OAI2BB2XL U1894 ( .B0(n6787), .B1(n112), .A0N(\ram[51][8] ), .A1N(n6559), 
        .Y(n1406) );
  OAI2BB2XL U1895 ( .B0(n6764), .B1(n112), .A0N(\ram[51][9] ), .A1N(n6559), 
        .Y(n1407) );
  OAI2BB2XL U1896 ( .B0(n6741), .B1(n112), .A0N(\ram[51][10] ), .A1N(n6559), 
        .Y(n1408) );
  OAI2BB2XL U1897 ( .B0(n6718), .B1(n112), .A0N(\ram[51][11] ), .A1N(n6559), 
        .Y(n1409) );
  OAI2BB2XL U1898 ( .B0(n6695), .B1(n112), .A0N(\ram[51][12] ), .A1N(n6559), 
        .Y(n1410) );
  OAI2BB2XL U1899 ( .B0(n6672), .B1(n112), .A0N(\ram[51][13] ), .A1N(n6559), 
        .Y(n1411) );
  OAI2BB2XL U1900 ( .B0(n6649), .B1(n112), .A0N(\ram[51][14] ), .A1N(n6559), 
        .Y(n1412) );
  OAI2BB2XL U1901 ( .B0(n6626), .B1(n112), .A0N(\ram[51][15] ), .A1N(n6559), 
        .Y(n1413) );
  OAI2BB2XL U1902 ( .B0(n6972), .B1(n114), .A0N(\ram[52][0] ), .A1N(n6558), 
        .Y(n1414) );
  OAI2BB2XL U1903 ( .B0(n6949), .B1(n114), .A0N(\ram[52][1] ), .A1N(n6558), 
        .Y(n1415) );
  OAI2BB2XL U1904 ( .B0(n6926), .B1(n114), .A0N(\ram[52][2] ), .A1N(n6558), 
        .Y(n1416) );
  OAI2BB2XL U1905 ( .B0(n6903), .B1(n114), .A0N(\ram[52][3] ), .A1N(n6558), 
        .Y(n1417) );
  OAI2BB2XL U1906 ( .B0(n6878), .B1(n114), .A0N(\ram[52][4] ), .A1N(n6558), 
        .Y(n1418) );
  OAI2BB2XL U1907 ( .B0(n6855), .B1(n114), .A0N(\ram[52][5] ), .A1N(n6558), 
        .Y(n1419) );
  OAI2BB2XL U1908 ( .B0(n6832), .B1(n114), .A0N(\ram[52][6] ), .A1N(n6558), 
        .Y(n1420) );
  OAI2BB2XL U1909 ( .B0(n6809), .B1(n114), .A0N(\ram[52][7] ), .A1N(n6558), 
        .Y(n1421) );
  OAI2BB2XL U1910 ( .B0(n6786), .B1(n114), .A0N(\ram[52][8] ), .A1N(n6558), 
        .Y(n1422) );
  OAI2BB2XL U1911 ( .B0(n6763), .B1(n114), .A0N(\ram[52][9] ), .A1N(n6558), 
        .Y(n1423) );
  OAI2BB2XL U1912 ( .B0(n6740), .B1(n114), .A0N(\ram[52][10] ), .A1N(n6558), 
        .Y(n1424) );
  OAI2BB2XL U1913 ( .B0(n6717), .B1(n114), .A0N(\ram[52][11] ), .A1N(n6558), 
        .Y(n1425) );
  OAI2BB2XL U1914 ( .B0(n6694), .B1(n114), .A0N(\ram[52][12] ), .A1N(n6558), 
        .Y(n1426) );
  OAI2BB2XL U1915 ( .B0(n6671), .B1(n114), .A0N(\ram[52][13] ), .A1N(n6558), 
        .Y(n1427) );
  OAI2BB2XL U1916 ( .B0(n6648), .B1(n114), .A0N(\ram[52][14] ), .A1N(n6558), 
        .Y(n1428) );
  OAI2BB2XL U1917 ( .B0(n6625), .B1(n114), .A0N(\ram[52][15] ), .A1N(n6558), 
        .Y(n1429) );
  OAI2BB2XL U1918 ( .B0(n6968), .B1(n116), .A0N(\ram[53][0] ), .A1N(n6557), 
        .Y(n1430) );
  OAI2BB2XL U1919 ( .B0(n6945), .B1(n116), .A0N(\ram[53][1] ), .A1N(n6557), 
        .Y(n1431) );
  OAI2BB2XL U1920 ( .B0(n6922), .B1(n116), .A0N(\ram[53][2] ), .A1N(n6557), 
        .Y(n1432) );
  OAI2BB2XL U1921 ( .B0(n6899), .B1(n116), .A0N(\ram[53][3] ), .A1N(n6557), 
        .Y(n1433) );
  OAI2BB2XL U1922 ( .B0(n6878), .B1(n116), .A0N(\ram[53][4] ), .A1N(n6557), 
        .Y(n1434) );
  OAI2BB2XL U1923 ( .B0(n6855), .B1(n116), .A0N(\ram[53][5] ), .A1N(n6557), 
        .Y(n1435) );
  OAI2BB2XL U1924 ( .B0(n6832), .B1(n116), .A0N(\ram[53][6] ), .A1N(n6557), 
        .Y(n1436) );
  OAI2BB2XL U1925 ( .B0(n6809), .B1(n116), .A0N(\ram[53][7] ), .A1N(n6557), 
        .Y(n1437) );
  OAI2BB2XL U1926 ( .B0(n6786), .B1(n116), .A0N(\ram[53][8] ), .A1N(n6557), 
        .Y(n1438) );
  OAI2BB2XL U1927 ( .B0(n6763), .B1(n116), .A0N(\ram[53][9] ), .A1N(n6557), 
        .Y(n1439) );
  OAI2BB2XL U1928 ( .B0(n6740), .B1(n116), .A0N(\ram[53][10] ), .A1N(n6557), 
        .Y(n1440) );
  OAI2BB2XL U1929 ( .B0(n6717), .B1(n116), .A0N(\ram[53][11] ), .A1N(n6557), 
        .Y(n1441) );
  OAI2BB2XL U1930 ( .B0(n6694), .B1(n116), .A0N(\ram[53][12] ), .A1N(n6557), 
        .Y(n1442) );
  OAI2BB2XL U1931 ( .B0(n6671), .B1(n116), .A0N(\ram[53][13] ), .A1N(n6557), 
        .Y(n1443) );
  OAI2BB2XL U1932 ( .B0(n6648), .B1(n116), .A0N(\ram[53][14] ), .A1N(n6557), 
        .Y(n1444) );
  OAI2BB2XL U1933 ( .B0(n6625), .B1(n116), .A0N(\ram[53][15] ), .A1N(n6557), 
        .Y(n1445) );
  OAI2BB2XL U1934 ( .B0(n6971), .B1(n118), .A0N(\ram[54][0] ), .A1N(n6556), 
        .Y(n1446) );
  OAI2BB2XL U1935 ( .B0(n6948), .B1(n118), .A0N(\ram[54][1] ), .A1N(n6556), 
        .Y(n1447) );
  OAI2BB2XL U1936 ( .B0(n6925), .B1(n118), .A0N(\ram[54][2] ), .A1N(n6556), 
        .Y(n1448) );
  OAI2BB2XL U1937 ( .B0(n6902), .B1(n118), .A0N(\ram[54][3] ), .A1N(n6556), 
        .Y(n1449) );
  OAI2BB2XL U1938 ( .B0(n6878), .B1(n118), .A0N(\ram[54][4] ), .A1N(n6556), 
        .Y(n1450) );
  OAI2BB2XL U1939 ( .B0(n6855), .B1(n118), .A0N(\ram[54][5] ), .A1N(n6556), 
        .Y(n1451) );
  OAI2BB2XL U1940 ( .B0(n6832), .B1(n118), .A0N(\ram[54][6] ), .A1N(n6556), 
        .Y(n1452) );
  OAI2BB2XL U1941 ( .B0(n6809), .B1(n118), .A0N(\ram[54][7] ), .A1N(n6556), 
        .Y(n1453) );
  OAI2BB2XL U1942 ( .B0(n6786), .B1(n118), .A0N(\ram[54][8] ), .A1N(n6556), 
        .Y(n1454) );
  OAI2BB2XL U1943 ( .B0(n6763), .B1(n118), .A0N(\ram[54][9] ), .A1N(n6556), 
        .Y(n1455) );
  OAI2BB2XL U1944 ( .B0(n6740), .B1(n118), .A0N(\ram[54][10] ), .A1N(n6556), 
        .Y(n1456) );
  OAI2BB2XL U1945 ( .B0(n6717), .B1(n118), .A0N(\ram[54][11] ), .A1N(n6556), 
        .Y(n1457) );
  OAI2BB2XL U1946 ( .B0(n6694), .B1(n118), .A0N(\ram[54][12] ), .A1N(n6556), 
        .Y(n1458) );
  OAI2BB2XL U1947 ( .B0(n6671), .B1(n118), .A0N(\ram[54][13] ), .A1N(n6556), 
        .Y(n1459) );
  OAI2BB2XL U1948 ( .B0(n6648), .B1(n118), .A0N(\ram[54][14] ), .A1N(n6556), 
        .Y(n1460) );
  OAI2BB2XL U1949 ( .B0(n6625), .B1(n118), .A0N(\ram[54][15] ), .A1N(n6556), 
        .Y(n1461) );
  OAI2BB2XL U1950 ( .B0(n6967), .B1(n120), .A0N(\ram[55][0] ), .A1N(n6555), 
        .Y(n1462) );
  OAI2BB2XL U1951 ( .B0(n6944), .B1(n120), .A0N(\ram[55][1] ), .A1N(n6555), 
        .Y(n1463) );
  OAI2BB2XL U1952 ( .B0(n6921), .B1(n120), .A0N(\ram[55][2] ), .A1N(n6555), 
        .Y(n1464) );
  OAI2BB2XL U1953 ( .B0(n6898), .B1(n120), .A0N(\ram[55][3] ), .A1N(n6555), 
        .Y(n1465) );
  OAI2BB2XL U1954 ( .B0(n6878), .B1(n120), .A0N(\ram[55][4] ), .A1N(n6555), 
        .Y(n1466) );
  OAI2BB2XL U1955 ( .B0(n6855), .B1(n120), .A0N(\ram[55][5] ), .A1N(n6555), 
        .Y(n1467) );
  OAI2BB2XL U1956 ( .B0(n6832), .B1(n120), .A0N(\ram[55][6] ), .A1N(n6555), 
        .Y(n1468) );
  OAI2BB2XL U1957 ( .B0(n6809), .B1(n120), .A0N(\ram[55][7] ), .A1N(n6555), 
        .Y(n1469) );
  OAI2BB2XL U1958 ( .B0(n6786), .B1(n120), .A0N(\ram[55][8] ), .A1N(n6555), 
        .Y(n1470) );
  OAI2BB2XL U1959 ( .B0(n6763), .B1(n120), .A0N(\ram[55][9] ), .A1N(n6555), 
        .Y(n1471) );
  OAI2BB2XL U1960 ( .B0(n6740), .B1(n120), .A0N(\ram[55][10] ), .A1N(n6555), 
        .Y(n1472) );
  OAI2BB2XL U1961 ( .B0(n6717), .B1(n120), .A0N(\ram[55][11] ), .A1N(n6555), 
        .Y(n1473) );
  OAI2BB2XL U1962 ( .B0(n6694), .B1(n120), .A0N(\ram[55][12] ), .A1N(n6555), 
        .Y(n1474) );
  OAI2BB2XL U1963 ( .B0(n6671), .B1(n120), .A0N(\ram[55][13] ), .A1N(n6555), 
        .Y(n1475) );
  OAI2BB2XL U1964 ( .B0(n6648), .B1(n120), .A0N(\ram[55][14] ), .A1N(n6555), 
        .Y(n1476) );
  OAI2BB2XL U1965 ( .B0(n6625), .B1(n120), .A0N(\ram[55][15] ), .A1N(n6555), 
        .Y(n1477) );
  OAI2BB2XL U1966 ( .B0(n6970), .B1(n122), .A0N(\ram[56][0] ), .A1N(n6554), 
        .Y(n1478) );
  OAI2BB2XL U1967 ( .B0(n6947), .B1(n122), .A0N(\ram[56][1] ), .A1N(n6554), 
        .Y(n1479) );
  OAI2BB2XL U1968 ( .B0(n6924), .B1(n122), .A0N(\ram[56][2] ), .A1N(n6554), 
        .Y(n1480) );
  OAI2BB2XL U1969 ( .B0(n6901), .B1(n122), .A0N(\ram[56][3] ), .A1N(n6554), 
        .Y(n1481) );
  OAI2BB2XL U1970 ( .B0(n6878), .B1(n122), .A0N(\ram[56][4] ), .A1N(n6554), 
        .Y(n1482) );
  OAI2BB2XL U1971 ( .B0(n6855), .B1(n122), .A0N(\ram[56][5] ), .A1N(n6554), 
        .Y(n1483) );
  OAI2BB2XL U1972 ( .B0(n6832), .B1(n122), .A0N(\ram[56][6] ), .A1N(n6554), 
        .Y(n1484) );
  OAI2BB2XL U1973 ( .B0(n6809), .B1(n122), .A0N(\ram[56][7] ), .A1N(n6554), 
        .Y(n1485) );
  OAI2BB2XL U1974 ( .B0(n6786), .B1(n122), .A0N(\ram[56][8] ), .A1N(n6554), 
        .Y(n1486) );
  OAI2BB2XL U1975 ( .B0(n6763), .B1(n122), .A0N(\ram[56][9] ), .A1N(n6554), 
        .Y(n1487) );
  OAI2BB2XL U1976 ( .B0(n6740), .B1(n122), .A0N(\ram[56][10] ), .A1N(n6554), 
        .Y(n1488) );
  OAI2BB2XL U1977 ( .B0(n6717), .B1(n122), .A0N(\ram[56][11] ), .A1N(n6554), 
        .Y(n1489) );
  OAI2BB2XL U1978 ( .B0(n6694), .B1(n122), .A0N(\ram[56][12] ), .A1N(n6554), 
        .Y(n1490) );
  OAI2BB2XL U1979 ( .B0(n6671), .B1(n122), .A0N(\ram[56][13] ), .A1N(n6554), 
        .Y(n1491) );
  OAI2BB2XL U1980 ( .B0(n6648), .B1(n122), .A0N(\ram[56][14] ), .A1N(n6554), 
        .Y(n1492) );
  OAI2BB2XL U1981 ( .B0(n6625), .B1(n122), .A0N(\ram[56][15] ), .A1N(n6554), 
        .Y(n1493) );
  OAI2BB2XL U1982 ( .B0(n6956), .B1(n124), .A0N(\ram[57][0] ), .A1N(n6553), 
        .Y(n1494) );
  OAI2BB2XL U1983 ( .B0(n6933), .B1(n124), .A0N(\ram[57][1] ), .A1N(n6553), 
        .Y(n1495) );
  OAI2BB2XL U1984 ( .B0(n6910), .B1(n124), .A0N(\ram[57][2] ), .A1N(n6553), 
        .Y(n1496) );
  OAI2BB2XL U1985 ( .B0(n6887), .B1(n124), .A0N(\ram[57][3] ), .A1N(n6553), 
        .Y(n1497) );
  OAI2BB2XL U1986 ( .B0(n6878), .B1(n124), .A0N(\ram[57][4] ), .A1N(n6553), 
        .Y(n1498) );
  OAI2BB2XL U1987 ( .B0(n6855), .B1(n124), .A0N(\ram[57][5] ), .A1N(n6553), 
        .Y(n1499) );
  OAI2BB2XL U1988 ( .B0(n6832), .B1(n124), .A0N(\ram[57][6] ), .A1N(n6553), 
        .Y(n1500) );
  OAI2BB2XL U1989 ( .B0(n6809), .B1(n124), .A0N(\ram[57][7] ), .A1N(n6553), 
        .Y(n1501) );
  OAI2BB2XL U1990 ( .B0(n6786), .B1(n124), .A0N(\ram[57][8] ), .A1N(n6553), 
        .Y(n1502) );
  OAI2BB2XL U1991 ( .B0(n6763), .B1(n124), .A0N(\ram[57][9] ), .A1N(n6553), 
        .Y(n1503) );
  OAI2BB2XL U1992 ( .B0(n6740), .B1(n124), .A0N(\ram[57][10] ), .A1N(n6553), 
        .Y(n1504) );
  OAI2BB2XL U1993 ( .B0(n6717), .B1(n124), .A0N(\ram[57][11] ), .A1N(n6553), 
        .Y(n1505) );
  OAI2BB2XL U1994 ( .B0(n6694), .B1(n124), .A0N(\ram[57][12] ), .A1N(n6553), 
        .Y(n1506) );
  OAI2BB2XL U1995 ( .B0(n6671), .B1(n124), .A0N(\ram[57][13] ), .A1N(n6553), 
        .Y(n1507) );
  OAI2BB2XL U1996 ( .B0(n6648), .B1(n124), .A0N(\ram[57][14] ), .A1N(n6553), 
        .Y(n1508) );
  OAI2BB2XL U1997 ( .B0(n6625), .B1(n124), .A0N(\ram[57][15] ), .A1N(n6553), 
        .Y(n1509) );
  OAI2BB2XL U1998 ( .B0(n6964), .B1(n126), .A0N(\ram[58][0] ), .A1N(n6552), 
        .Y(n1510) );
  OAI2BB2XL U1999 ( .B0(n6941), .B1(n126), .A0N(\ram[58][1] ), .A1N(n6552), 
        .Y(n1511) );
  OAI2BB2XL U2000 ( .B0(n6918), .B1(n126), .A0N(\ram[58][2] ), .A1N(n6552), 
        .Y(n1512) );
  OAI2BB2XL U2001 ( .B0(n6895), .B1(n126), .A0N(\ram[58][3] ), .A1N(n6552), 
        .Y(n1513) );
  OAI2BB2XL U2002 ( .B0(n6878), .B1(n126), .A0N(\ram[58][4] ), .A1N(n6552), 
        .Y(n1514) );
  OAI2BB2XL U2003 ( .B0(n6855), .B1(n126), .A0N(\ram[58][5] ), .A1N(n6552), 
        .Y(n1515) );
  OAI2BB2XL U2004 ( .B0(n6832), .B1(n126), .A0N(\ram[58][6] ), .A1N(n6552), 
        .Y(n1516) );
  OAI2BB2XL U2005 ( .B0(n6809), .B1(n126), .A0N(\ram[58][7] ), .A1N(n6552), 
        .Y(n1517) );
  OAI2BB2XL U2006 ( .B0(n6786), .B1(n126), .A0N(\ram[58][8] ), .A1N(n6552), 
        .Y(n1518) );
  OAI2BB2XL U2007 ( .B0(n6763), .B1(n126), .A0N(\ram[58][9] ), .A1N(n6552), 
        .Y(n1519) );
  OAI2BB2XL U2008 ( .B0(n6740), .B1(n126), .A0N(\ram[58][10] ), .A1N(n6552), 
        .Y(n1520) );
  OAI2BB2XL U2009 ( .B0(n6717), .B1(n126), .A0N(\ram[58][11] ), .A1N(n6552), 
        .Y(n1521) );
  OAI2BB2XL U2010 ( .B0(n6694), .B1(n126), .A0N(\ram[58][12] ), .A1N(n6552), 
        .Y(n1522) );
  OAI2BB2XL U2011 ( .B0(n6671), .B1(n126), .A0N(\ram[58][13] ), .A1N(n6552), 
        .Y(n1523) );
  OAI2BB2XL U2012 ( .B0(n6648), .B1(n126), .A0N(\ram[58][14] ), .A1N(n6552), 
        .Y(n1524) );
  OAI2BB2XL U2013 ( .B0(n6625), .B1(n126), .A0N(\ram[58][15] ), .A1N(n6552), 
        .Y(n1525) );
  OAI2BB2XL U2014 ( .B0(n6963), .B1(n128), .A0N(\ram[59][0] ), .A1N(n6551), 
        .Y(n1526) );
  OAI2BB2XL U2015 ( .B0(n6940), .B1(n128), .A0N(\ram[59][1] ), .A1N(n6551), 
        .Y(n1527) );
  OAI2BB2XL U2016 ( .B0(n6917), .B1(n128), .A0N(\ram[59][2] ), .A1N(n6551), 
        .Y(n1528) );
  OAI2BB2XL U2017 ( .B0(n6894), .B1(n128), .A0N(\ram[59][3] ), .A1N(n6551), 
        .Y(n1529) );
  OAI2BB2XL U2018 ( .B0(n6878), .B1(n128), .A0N(\ram[59][4] ), .A1N(n6551), 
        .Y(n1530) );
  OAI2BB2XL U2019 ( .B0(n6855), .B1(n128), .A0N(\ram[59][5] ), .A1N(n6551), 
        .Y(n1531) );
  OAI2BB2XL U2020 ( .B0(n6832), .B1(n128), .A0N(\ram[59][6] ), .A1N(n6551), 
        .Y(n1532) );
  OAI2BB2XL U2021 ( .B0(n6809), .B1(n128), .A0N(\ram[59][7] ), .A1N(n6551), 
        .Y(n1533) );
  OAI2BB2XL U2022 ( .B0(n6786), .B1(n128), .A0N(\ram[59][8] ), .A1N(n6551), 
        .Y(n1534) );
  OAI2BB2XL U2023 ( .B0(n6763), .B1(n128), .A0N(\ram[59][9] ), .A1N(n6551), 
        .Y(n1535) );
  OAI2BB2XL U2024 ( .B0(n6740), .B1(n128), .A0N(\ram[59][10] ), .A1N(n6551), 
        .Y(n1536) );
  OAI2BB2XL U2025 ( .B0(n6717), .B1(n128), .A0N(\ram[59][11] ), .A1N(n6551), 
        .Y(n1537) );
  OAI2BB2XL U2026 ( .B0(n6694), .B1(n128), .A0N(\ram[59][12] ), .A1N(n6551), 
        .Y(n1538) );
  OAI2BB2XL U2027 ( .B0(n6671), .B1(n128), .A0N(\ram[59][13] ), .A1N(n6551), 
        .Y(n1539) );
  OAI2BB2XL U2028 ( .B0(n6648), .B1(n128), .A0N(\ram[59][14] ), .A1N(n6551), 
        .Y(n1540) );
  OAI2BB2XL U2029 ( .B0(n6625), .B1(n128), .A0N(\ram[59][15] ), .A1N(n6551), 
        .Y(n1541) );
  OAI2BB2XL U2030 ( .B0(n6956), .B1(n130), .A0N(\ram[60][0] ), .A1N(n6550), 
        .Y(n1542) );
  OAI2BB2XL U2031 ( .B0(n6933), .B1(n130), .A0N(\ram[60][1] ), .A1N(n6550), 
        .Y(n1543) );
  OAI2BB2XL U2032 ( .B0(n6910), .B1(n130), .A0N(\ram[60][2] ), .A1N(n6550), 
        .Y(n1544) );
  OAI2BB2XL U2033 ( .B0(n6887), .B1(n130), .A0N(\ram[60][3] ), .A1N(n6550), 
        .Y(n1545) );
  OAI2BB2XL U2034 ( .B0(n6878), .B1(n130), .A0N(\ram[60][4] ), .A1N(n6550), 
        .Y(n1546) );
  OAI2BB2XL U2035 ( .B0(n6855), .B1(n130), .A0N(\ram[60][5] ), .A1N(n6550), 
        .Y(n1547) );
  OAI2BB2XL U2036 ( .B0(n6832), .B1(n130), .A0N(\ram[60][6] ), .A1N(n6550), 
        .Y(n1548) );
  OAI2BB2XL U2037 ( .B0(n6809), .B1(n130), .A0N(\ram[60][7] ), .A1N(n6550), 
        .Y(n1549) );
  OAI2BB2XL U2038 ( .B0(n6786), .B1(n130), .A0N(\ram[60][8] ), .A1N(n6550), 
        .Y(n1550) );
  OAI2BB2XL U2039 ( .B0(n6763), .B1(n130), .A0N(\ram[60][9] ), .A1N(n6550), 
        .Y(n1551) );
  OAI2BB2XL U2040 ( .B0(n6740), .B1(n130), .A0N(\ram[60][10] ), .A1N(n6550), 
        .Y(n1552) );
  OAI2BB2XL U2041 ( .B0(n6717), .B1(n130), .A0N(\ram[60][11] ), .A1N(n6550), 
        .Y(n1553) );
  OAI2BB2XL U2042 ( .B0(n6694), .B1(n130), .A0N(\ram[60][12] ), .A1N(n6550), 
        .Y(n1554) );
  OAI2BB2XL U2043 ( .B0(n6671), .B1(n130), .A0N(\ram[60][13] ), .A1N(n6550), 
        .Y(n1555) );
  OAI2BB2XL U2044 ( .B0(n6648), .B1(n130), .A0N(\ram[60][14] ), .A1N(n6550), 
        .Y(n1556) );
  OAI2BB2XL U2045 ( .B0(n6625), .B1(n130), .A0N(\ram[60][15] ), .A1N(n6550), 
        .Y(n1557) );
  OAI2BB2XL U2046 ( .B0(n6957), .B1(n132), .A0N(\ram[61][0] ), .A1N(n6549), 
        .Y(n1558) );
  OAI2BB2XL U2047 ( .B0(n6934), .B1(n132), .A0N(\ram[61][1] ), .A1N(n6549), 
        .Y(n1559) );
  OAI2BB2XL U2048 ( .B0(n6911), .B1(n132), .A0N(\ram[61][2] ), .A1N(n6549), 
        .Y(n1560) );
  OAI2BB2XL U2049 ( .B0(n6888), .B1(n132), .A0N(\ram[61][3] ), .A1N(n6549), 
        .Y(n1561) );
  OAI2BB2XL U2050 ( .B0(n6878), .B1(n132), .A0N(\ram[61][4] ), .A1N(n6549), 
        .Y(n1562) );
  OAI2BB2XL U2051 ( .B0(n6855), .B1(n132), .A0N(\ram[61][5] ), .A1N(n6549), 
        .Y(n1563) );
  OAI2BB2XL U2052 ( .B0(n6832), .B1(n132), .A0N(\ram[61][6] ), .A1N(n6549), 
        .Y(n1564) );
  OAI2BB2XL U2053 ( .B0(n6809), .B1(n132), .A0N(\ram[61][7] ), .A1N(n6549), 
        .Y(n1565) );
  OAI2BB2XL U2054 ( .B0(n6786), .B1(n132), .A0N(\ram[61][8] ), .A1N(n6549), 
        .Y(n1566) );
  OAI2BB2XL U2055 ( .B0(n6763), .B1(n132), .A0N(\ram[61][9] ), .A1N(n6549), 
        .Y(n1567) );
  OAI2BB2XL U2056 ( .B0(n6740), .B1(n132), .A0N(\ram[61][10] ), .A1N(n6549), 
        .Y(n1568) );
  OAI2BB2XL U2057 ( .B0(n6717), .B1(n132), .A0N(\ram[61][11] ), .A1N(n6549), 
        .Y(n1569) );
  OAI2BB2XL U2058 ( .B0(n6694), .B1(n132), .A0N(\ram[61][12] ), .A1N(n6549), 
        .Y(n1570) );
  OAI2BB2XL U2059 ( .B0(n6671), .B1(n132), .A0N(\ram[61][13] ), .A1N(n6549), 
        .Y(n1571) );
  OAI2BB2XL U2060 ( .B0(n6648), .B1(n132), .A0N(\ram[61][14] ), .A1N(n6549), 
        .Y(n1572) );
  OAI2BB2XL U2061 ( .B0(n6625), .B1(n132), .A0N(\ram[61][15] ), .A1N(n6549), 
        .Y(n1573) );
  OAI2BB2XL U2062 ( .B0(n7), .B1(n498), .A0N(\ram[62][0] ), .A1N(n6548), .Y(
        n1574) );
  OAI2BB2XL U2063 ( .B0(n9), .B1(n498), .A0N(\ram[62][1] ), .A1N(n6548), .Y(
        n1575) );
  OAI2BB2XL U2064 ( .B0(n10), .B1(n498), .A0N(\ram[62][2] ), .A1N(n6548), .Y(
        n1576) );
  OAI2BB2XL U2065 ( .B0(n11), .B1(n498), .A0N(\ram[62][3] ), .A1N(n6548), .Y(
        n1577) );
  OAI2BB2XL U2066 ( .B0(n6878), .B1(n498), .A0N(\ram[62][4] ), .A1N(n6548), 
        .Y(n1578) );
  OAI2BB2XL U2067 ( .B0(n6855), .B1(n498), .A0N(\ram[62][5] ), .A1N(n6548), 
        .Y(n1579) );
  OAI2BB2XL U2068 ( .B0(n6832), .B1(n498), .A0N(\ram[62][6] ), .A1N(n6548), 
        .Y(n1580) );
  OAI2BB2XL U2069 ( .B0(n6809), .B1(n498), .A0N(\ram[62][7] ), .A1N(n6548), 
        .Y(n1581) );
  OAI2BB2XL U2070 ( .B0(n6786), .B1(n498), .A0N(\ram[62][8] ), .A1N(n6548), 
        .Y(n1582) );
  OAI2BB2XL U2071 ( .B0(n6763), .B1(n498), .A0N(\ram[62][9] ), .A1N(n6548), 
        .Y(n1583) );
  OAI2BB2XL U2072 ( .B0(n6740), .B1(n498), .A0N(\ram[62][10] ), .A1N(n6548), 
        .Y(n1584) );
  OAI2BB2XL U2073 ( .B0(n6717), .B1(n498), .A0N(\ram[62][11] ), .A1N(n6548), 
        .Y(n1585) );
  OAI2BB2XL U2074 ( .B0(n6694), .B1(n498), .A0N(\ram[62][12] ), .A1N(n6548), 
        .Y(n1586) );
  OAI2BB2XL U2075 ( .B0(n6671), .B1(n498), .A0N(\ram[62][13] ), .A1N(n6548), 
        .Y(n1587) );
  OAI2BB2XL U2076 ( .B0(n6648), .B1(n498), .A0N(\ram[62][14] ), .A1N(n6548), 
        .Y(n1588) );
  OAI2BB2XL U2077 ( .B0(n6625), .B1(n498), .A0N(\ram[62][15] ), .A1N(n6548), 
        .Y(n1589) );
  OAI2BB2XL U2078 ( .B0(n7), .B1(n134), .A0N(\ram[63][0] ), .A1N(n6547), .Y(
        n1590) );
  OAI2BB2XL U2079 ( .B0(n9), .B1(n134), .A0N(\ram[63][1] ), .A1N(n6547), .Y(
        n1591) );
  OAI2BB2XL U2080 ( .B0(n10), .B1(n134), .A0N(\ram[63][2] ), .A1N(n6547), .Y(
        n1592) );
  OAI2BB2XL U2081 ( .B0(n11), .B1(n134), .A0N(\ram[63][3] ), .A1N(n6547), .Y(
        n1593) );
  OAI2BB2XL U2082 ( .B0(n6878), .B1(n134), .A0N(\ram[63][4] ), .A1N(n6547), 
        .Y(n1594) );
  OAI2BB2XL U2083 ( .B0(n6855), .B1(n134), .A0N(\ram[63][5] ), .A1N(n6547), 
        .Y(n1595) );
  OAI2BB2XL U2084 ( .B0(n6832), .B1(n134), .A0N(\ram[63][6] ), .A1N(n6547), 
        .Y(n1596) );
  OAI2BB2XL U2085 ( .B0(n6809), .B1(n134), .A0N(\ram[63][7] ), .A1N(n6547), 
        .Y(n1597) );
  OAI2BB2XL U2086 ( .B0(n6786), .B1(n134), .A0N(\ram[63][8] ), .A1N(n6547), 
        .Y(n1598) );
  OAI2BB2XL U2087 ( .B0(n6763), .B1(n134), .A0N(\ram[63][9] ), .A1N(n6547), 
        .Y(n1599) );
  OAI2BB2XL U2088 ( .B0(n6740), .B1(n134), .A0N(\ram[63][10] ), .A1N(n6547), 
        .Y(n1600) );
  OAI2BB2XL U2089 ( .B0(n6717), .B1(n134), .A0N(\ram[63][11] ), .A1N(n6547), 
        .Y(n1601) );
  OAI2BB2XL U2090 ( .B0(n6694), .B1(n134), .A0N(\ram[63][12] ), .A1N(n6547), 
        .Y(n1602) );
  OAI2BB2XL U2091 ( .B0(n6671), .B1(n134), .A0N(\ram[63][13] ), .A1N(n6547), 
        .Y(n1603) );
  OAI2BB2XL U2092 ( .B0(n6648), .B1(n134), .A0N(\ram[63][14] ), .A1N(n6547), 
        .Y(n1604) );
  OAI2BB2XL U2093 ( .B0(n6625), .B1(n134), .A0N(\ram[63][15] ), .A1N(n6547), 
        .Y(n1605) );
  OAI2BB2XL U2094 ( .B0(n6973), .B1(n168), .A0N(\ram[80][0] ), .A1N(n6530), 
        .Y(n1862) );
  OAI2BB2XL U2095 ( .B0(n6950), .B1(n168), .A0N(\ram[80][1] ), .A1N(n6530), 
        .Y(n1863) );
  OAI2BB2XL U2096 ( .B0(n6927), .B1(n168), .A0N(\ram[80][2] ), .A1N(n6530), 
        .Y(n1864) );
  OAI2BB2XL U2097 ( .B0(n6904), .B1(n168), .A0N(\ram[80][3] ), .A1N(n6530), 
        .Y(n1865) );
  OAI2BB2XL U2098 ( .B0(n6876), .B1(n168), .A0N(\ram[80][4] ), .A1N(n6530), 
        .Y(n1866) );
  OAI2BB2XL U2099 ( .B0(n6853), .B1(n168), .A0N(\ram[80][5] ), .A1N(n6530), 
        .Y(n1867) );
  OAI2BB2XL U2100 ( .B0(n6830), .B1(n168), .A0N(\ram[80][6] ), .A1N(n6530), 
        .Y(n1868) );
  OAI2BB2XL U2101 ( .B0(n6807), .B1(n168), .A0N(\ram[80][7] ), .A1N(n6530), 
        .Y(n1869) );
  OAI2BB2XL U2102 ( .B0(n6784), .B1(n168), .A0N(\ram[80][8] ), .A1N(n6530), 
        .Y(n1870) );
  OAI2BB2XL U2103 ( .B0(n6761), .B1(n168), .A0N(\ram[80][9] ), .A1N(n6530), 
        .Y(n1871) );
  OAI2BB2XL U2104 ( .B0(n6738), .B1(n168), .A0N(\ram[80][10] ), .A1N(n6530), 
        .Y(n1872) );
  OAI2BB2XL U2105 ( .B0(n6715), .B1(n168), .A0N(\ram[80][11] ), .A1N(n6530), 
        .Y(n1873) );
  OAI2BB2XL U2106 ( .B0(n6692), .B1(n168), .A0N(\ram[80][12] ), .A1N(n6530), 
        .Y(n1874) );
  OAI2BB2XL U2107 ( .B0(n6669), .B1(n168), .A0N(\ram[80][13] ), .A1N(n6530), 
        .Y(n1875) );
  OAI2BB2XL U2108 ( .B0(n6646), .B1(n168), .A0N(\ram[80][14] ), .A1N(n6530), 
        .Y(n1876) );
  OAI2BB2XL U2109 ( .B0(n6623), .B1(n168), .A0N(\ram[80][15] ), .A1N(n6530), 
        .Y(n1877) );
  OAI2BB2XL U2110 ( .B0(n6973), .B1(n170), .A0N(\ram[81][0] ), .A1N(n6529), 
        .Y(n1878) );
  OAI2BB2XL U2111 ( .B0(n6950), .B1(n170), .A0N(\ram[81][1] ), .A1N(n6529), 
        .Y(n1879) );
  OAI2BB2XL U2112 ( .B0(n6927), .B1(n170), .A0N(\ram[81][2] ), .A1N(n6529), 
        .Y(n1880) );
  OAI2BB2XL U2113 ( .B0(n6904), .B1(n170), .A0N(\ram[81][3] ), .A1N(n6529), 
        .Y(n1881) );
  OAI2BB2XL U2114 ( .B0(n6876), .B1(n170), .A0N(\ram[81][4] ), .A1N(n6529), 
        .Y(n1882) );
  OAI2BB2XL U2115 ( .B0(n6853), .B1(n170), .A0N(\ram[81][5] ), .A1N(n6529), 
        .Y(n1883) );
  OAI2BB2XL U2116 ( .B0(n6830), .B1(n170), .A0N(\ram[81][6] ), .A1N(n6529), 
        .Y(n1884) );
  OAI2BB2XL U2117 ( .B0(n6807), .B1(n170), .A0N(\ram[81][7] ), .A1N(n6529), 
        .Y(n1885) );
  OAI2BB2XL U2118 ( .B0(n6784), .B1(n170), .A0N(\ram[81][8] ), .A1N(n6529), 
        .Y(n1886) );
  OAI2BB2XL U2119 ( .B0(n6761), .B1(n170), .A0N(\ram[81][9] ), .A1N(n6529), 
        .Y(n1887) );
  OAI2BB2XL U2120 ( .B0(n6738), .B1(n170), .A0N(\ram[81][10] ), .A1N(n6529), 
        .Y(n1888) );
  OAI2BB2XL U2121 ( .B0(n6715), .B1(n170), .A0N(\ram[81][11] ), .A1N(n6529), 
        .Y(n1889) );
  OAI2BB2XL U2122 ( .B0(n6692), .B1(n170), .A0N(\ram[81][12] ), .A1N(n6529), 
        .Y(n1890) );
  OAI2BB2XL U2123 ( .B0(n6669), .B1(n170), .A0N(\ram[81][13] ), .A1N(n6529), 
        .Y(n1891) );
  OAI2BB2XL U2124 ( .B0(n6646), .B1(n170), .A0N(\ram[81][14] ), .A1N(n6529), 
        .Y(n1892) );
  OAI2BB2XL U2125 ( .B0(n6623), .B1(n170), .A0N(\ram[81][15] ), .A1N(n6529), 
        .Y(n1893) );
  OAI2BB2XL U2126 ( .B0(n6973), .B1(n172), .A0N(\ram[82][0] ), .A1N(n6528), 
        .Y(n1894) );
  OAI2BB2XL U2127 ( .B0(n6950), .B1(n172), .A0N(\ram[82][1] ), .A1N(n6528), 
        .Y(n1895) );
  OAI2BB2XL U2128 ( .B0(n6927), .B1(n172), .A0N(\ram[82][2] ), .A1N(n6528), 
        .Y(n1896) );
  OAI2BB2XL U2129 ( .B0(n6904), .B1(n172), .A0N(\ram[82][3] ), .A1N(n6528), 
        .Y(n1897) );
  OAI2BB2XL U2130 ( .B0(n6876), .B1(n172), .A0N(\ram[82][4] ), .A1N(n6528), 
        .Y(n1898) );
  OAI2BB2XL U2131 ( .B0(n6853), .B1(n172), .A0N(\ram[82][5] ), .A1N(n6528), 
        .Y(n1899) );
  OAI2BB2XL U2132 ( .B0(n6830), .B1(n172), .A0N(\ram[82][6] ), .A1N(n6528), 
        .Y(n1900) );
  OAI2BB2XL U2133 ( .B0(n6807), .B1(n172), .A0N(\ram[82][7] ), .A1N(n6528), 
        .Y(n1901) );
  OAI2BB2XL U2134 ( .B0(n6784), .B1(n172), .A0N(\ram[82][8] ), .A1N(n6528), 
        .Y(n1902) );
  OAI2BB2XL U2135 ( .B0(n6761), .B1(n172), .A0N(\ram[82][9] ), .A1N(n6528), 
        .Y(n1903) );
  OAI2BB2XL U2136 ( .B0(n6738), .B1(n172), .A0N(\ram[82][10] ), .A1N(n6528), 
        .Y(n1904) );
  OAI2BB2XL U2137 ( .B0(n6715), .B1(n172), .A0N(\ram[82][11] ), .A1N(n6528), 
        .Y(n1905) );
  OAI2BB2XL U2138 ( .B0(n6692), .B1(n172), .A0N(\ram[82][12] ), .A1N(n6528), 
        .Y(n1906) );
  OAI2BB2XL U2139 ( .B0(n6669), .B1(n172), .A0N(\ram[82][13] ), .A1N(n6528), 
        .Y(n1907) );
  OAI2BB2XL U2140 ( .B0(n6646), .B1(n172), .A0N(\ram[82][14] ), .A1N(n6528), 
        .Y(n1908) );
  OAI2BB2XL U2141 ( .B0(n6623), .B1(n172), .A0N(\ram[82][15] ), .A1N(n6528), 
        .Y(n1909) );
  OAI2BB2XL U2142 ( .B0(n6973), .B1(n175), .A0N(\ram[83][0] ), .A1N(n6527), 
        .Y(n1910) );
  OAI2BB2XL U2143 ( .B0(n6950), .B1(n175), .A0N(\ram[83][1] ), .A1N(n6527), 
        .Y(n1911) );
  OAI2BB2XL U2144 ( .B0(n6927), .B1(n175), .A0N(\ram[83][2] ), .A1N(n6527), 
        .Y(n1912) );
  OAI2BB2XL U2145 ( .B0(n6904), .B1(n175), .A0N(\ram[83][3] ), .A1N(n6527), 
        .Y(n1913) );
  OAI2BB2XL U2146 ( .B0(n6876), .B1(n175), .A0N(\ram[83][4] ), .A1N(n6527), 
        .Y(n1914) );
  OAI2BB2XL U2147 ( .B0(n6853), .B1(n175), .A0N(\ram[83][5] ), .A1N(n6527), 
        .Y(n1915) );
  OAI2BB2XL U2148 ( .B0(n6830), .B1(n175), .A0N(\ram[83][6] ), .A1N(n6527), 
        .Y(n1916) );
  OAI2BB2XL U2149 ( .B0(n6807), .B1(n175), .A0N(\ram[83][7] ), .A1N(n6527), 
        .Y(n1917) );
  OAI2BB2XL U2150 ( .B0(n6784), .B1(n175), .A0N(\ram[83][8] ), .A1N(n6527), 
        .Y(n1918) );
  OAI2BB2XL U2151 ( .B0(n6761), .B1(n175), .A0N(\ram[83][9] ), .A1N(n6527), 
        .Y(n1919) );
  OAI2BB2XL U2152 ( .B0(n6738), .B1(n175), .A0N(\ram[83][10] ), .A1N(n6527), 
        .Y(n1920) );
  OAI2BB2XL U2153 ( .B0(n6715), .B1(n175), .A0N(\ram[83][11] ), .A1N(n6527), 
        .Y(n1921) );
  OAI2BB2XL U2154 ( .B0(n6692), .B1(n175), .A0N(\ram[83][12] ), .A1N(n6527), 
        .Y(n1922) );
  OAI2BB2XL U2155 ( .B0(n6669), .B1(n175), .A0N(\ram[83][13] ), .A1N(n6527), 
        .Y(n1923) );
  OAI2BB2XL U2156 ( .B0(n6646), .B1(n175), .A0N(\ram[83][14] ), .A1N(n6527), 
        .Y(n1924) );
  OAI2BB2XL U2157 ( .B0(n6623), .B1(n175), .A0N(\ram[83][15] ), .A1N(n6527), 
        .Y(n1925) );
  OAI2BB2XL U2158 ( .B0(n6973), .B1(n177), .A0N(\ram[84][0] ), .A1N(n6526), 
        .Y(n1926) );
  OAI2BB2XL U2159 ( .B0(n6950), .B1(n177), .A0N(\ram[84][1] ), .A1N(n6526), 
        .Y(n1927) );
  OAI2BB2XL U2160 ( .B0(n6927), .B1(n177), .A0N(\ram[84][2] ), .A1N(n6526), 
        .Y(n1928) );
  OAI2BB2XL U2161 ( .B0(n6904), .B1(n177), .A0N(\ram[84][3] ), .A1N(n6526), 
        .Y(n1929) );
  OAI2BB2XL U2162 ( .B0(n6876), .B1(n177), .A0N(\ram[84][4] ), .A1N(n6526), 
        .Y(n1930) );
  OAI2BB2XL U2163 ( .B0(n6853), .B1(n177), .A0N(\ram[84][5] ), .A1N(n6526), 
        .Y(n1931) );
  OAI2BB2XL U2164 ( .B0(n6830), .B1(n177), .A0N(\ram[84][6] ), .A1N(n6526), 
        .Y(n1932) );
  OAI2BB2XL U2165 ( .B0(n6807), .B1(n177), .A0N(\ram[84][7] ), .A1N(n6526), 
        .Y(n1933) );
  OAI2BB2XL U2166 ( .B0(n6784), .B1(n177), .A0N(\ram[84][8] ), .A1N(n6526), 
        .Y(n1934) );
  OAI2BB2XL U2167 ( .B0(n6761), .B1(n177), .A0N(\ram[84][9] ), .A1N(n6526), 
        .Y(n1935) );
  OAI2BB2XL U2168 ( .B0(n6738), .B1(n177), .A0N(\ram[84][10] ), .A1N(n6526), 
        .Y(n1936) );
  OAI2BB2XL U2169 ( .B0(n6715), .B1(n177), .A0N(\ram[84][11] ), .A1N(n6526), 
        .Y(n1937) );
  OAI2BB2XL U2170 ( .B0(n6692), .B1(n177), .A0N(\ram[84][12] ), .A1N(n6526), 
        .Y(n1938) );
  OAI2BB2XL U2171 ( .B0(n6669), .B1(n177), .A0N(\ram[84][13] ), .A1N(n6526), 
        .Y(n1939) );
  OAI2BB2XL U2172 ( .B0(n6646), .B1(n177), .A0N(\ram[84][14] ), .A1N(n6526), 
        .Y(n1940) );
  OAI2BB2XL U2173 ( .B0(n6623), .B1(n177), .A0N(\ram[84][15] ), .A1N(n6526), 
        .Y(n1941) );
  OAI2BB2XL U2174 ( .B0(n6973), .B1(n178), .A0N(\ram[85][0] ), .A1N(n6525), 
        .Y(n1942) );
  OAI2BB2XL U2175 ( .B0(n6950), .B1(n178), .A0N(\ram[85][1] ), .A1N(n6525), 
        .Y(n1943) );
  OAI2BB2XL U2176 ( .B0(n6927), .B1(n178), .A0N(\ram[85][2] ), .A1N(n6525), 
        .Y(n1944) );
  OAI2BB2XL U2177 ( .B0(n6904), .B1(n178), .A0N(\ram[85][3] ), .A1N(n6525), 
        .Y(n1945) );
  OAI2BB2XL U2178 ( .B0(n6876), .B1(n178), .A0N(\ram[85][4] ), .A1N(n6525), 
        .Y(n1946) );
  OAI2BB2XL U2179 ( .B0(n6853), .B1(n178), .A0N(\ram[85][5] ), .A1N(n6525), 
        .Y(n1947) );
  OAI2BB2XL U2180 ( .B0(n6830), .B1(n178), .A0N(\ram[85][6] ), .A1N(n6525), 
        .Y(n1948) );
  OAI2BB2XL U2181 ( .B0(n6807), .B1(n178), .A0N(\ram[85][7] ), .A1N(n6525), 
        .Y(n1949) );
  OAI2BB2XL U2182 ( .B0(n6784), .B1(n178), .A0N(\ram[85][8] ), .A1N(n6525), 
        .Y(n1950) );
  OAI2BB2XL U2183 ( .B0(n6761), .B1(n178), .A0N(\ram[85][9] ), .A1N(n6525), 
        .Y(n1951) );
  OAI2BB2XL U2184 ( .B0(n6738), .B1(n178), .A0N(\ram[85][10] ), .A1N(n6525), 
        .Y(n1952) );
  OAI2BB2XL U2185 ( .B0(n6715), .B1(n178), .A0N(\ram[85][11] ), .A1N(n6525), 
        .Y(n1953) );
  OAI2BB2XL U2186 ( .B0(n6692), .B1(n178), .A0N(\ram[85][12] ), .A1N(n6525), 
        .Y(n1954) );
  OAI2BB2XL U2187 ( .B0(n6669), .B1(n178), .A0N(\ram[85][13] ), .A1N(n6525), 
        .Y(n1955) );
  OAI2BB2XL U2188 ( .B0(n6646), .B1(n178), .A0N(\ram[85][14] ), .A1N(n6525), 
        .Y(n1956) );
  OAI2BB2XL U2189 ( .B0(n6623), .B1(n178), .A0N(\ram[85][15] ), .A1N(n6525), 
        .Y(n1957) );
  OAI2BB2XL U2190 ( .B0(n6973), .B1(n180), .A0N(\ram[86][0] ), .A1N(n6524), 
        .Y(n1958) );
  OAI2BB2XL U2191 ( .B0(n6950), .B1(n180), .A0N(\ram[86][1] ), .A1N(n6524), 
        .Y(n1959) );
  OAI2BB2XL U2192 ( .B0(n6927), .B1(n180), .A0N(\ram[86][2] ), .A1N(n6524), 
        .Y(n1960) );
  OAI2BB2XL U2193 ( .B0(n6904), .B1(n180), .A0N(\ram[86][3] ), .A1N(n6524), 
        .Y(n1961) );
  OAI2BB2XL U2194 ( .B0(n6876), .B1(n180), .A0N(\ram[86][4] ), .A1N(n6524), 
        .Y(n1962) );
  OAI2BB2XL U2195 ( .B0(n6853), .B1(n180), .A0N(\ram[86][5] ), .A1N(n6524), 
        .Y(n1963) );
  OAI2BB2XL U2196 ( .B0(n6830), .B1(n180), .A0N(\ram[86][6] ), .A1N(n6524), 
        .Y(n1964) );
  OAI2BB2XL U2197 ( .B0(n6807), .B1(n180), .A0N(\ram[86][7] ), .A1N(n6524), 
        .Y(n1965) );
  OAI2BB2XL U2198 ( .B0(n6784), .B1(n180), .A0N(\ram[86][8] ), .A1N(n6524), 
        .Y(n1966) );
  OAI2BB2XL U2199 ( .B0(n6761), .B1(n180), .A0N(\ram[86][9] ), .A1N(n6524), 
        .Y(n1967) );
  OAI2BB2XL U2200 ( .B0(n6738), .B1(n180), .A0N(\ram[86][10] ), .A1N(n6524), 
        .Y(n1968) );
  OAI2BB2XL U2201 ( .B0(n6715), .B1(n180), .A0N(\ram[86][11] ), .A1N(n6524), 
        .Y(n1969) );
  OAI2BB2XL U2202 ( .B0(n6692), .B1(n180), .A0N(\ram[86][12] ), .A1N(n6524), 
        .Y(n1970) );
  OAI2BB2XL U2203 ( .B0(n6669), .B1(n180), .A0N(\ram[86][13] ), .A1N(n6524), 
        .Y(n1971) );
  OAI2BB2XL U2204 ( .B0(n6646), .B1(n180), .A0N(\ram[86][14] ), .A1N(n6524), 
        .Y(n1972) );
  OAI2BB2XL U2205 ( .B0(n6623), .B1(n180), .A0N(\ram[86][15] ), .A1N(n6524), 
        .Y(n1973) );
  OAI2BB2XL U2206 ( .B0(n6973), .B1(n182), .A0N(\ram[87][0] ), .A1N(n6523), 
        .Y(n1974) );
  OAI2BB2XL U2207 ( .B0(n6950), .B1(n182), .A0N(\ram[87][1] ), .A1N(n6523), 
        .Y(n1975) );
  OAI2BB2XL U2208 ( .B0(n6927), .B1(n182), .A0N(\ram[87][2] ), .A1N(n6523), 
        .Y(n1976) );
  OAI2BB2XL U2209 ( .B0(n6904), .B1(n182), .A0N(\ram[87][3] ), .A1N(n6523), 
        .Y(n1977) );
  OAI2BB2XL U2210 ( .B0(n6876), .B1(n182), .A0N(\ram[87][4] ), .A1N(n6523), 
        .Y(n1978) );
  OAI2BB2XL U2211 ( .B0(n6853), .B1(n182), .A0N(\ram[87][5] ), .A1N(n6523), 
        .Y(n1979) );
  OAI2BB2XL U2212 ( .B0(n6830), .B1(n182), .A0N(\ram[87][6] ), .A1N(n6523), 
        .Y(n1980) );
  OAI2BB2XL U2213 ( .B0(n6807), .B1(n182), .A0N(\ram[87][7] ), .A1N(n6523), 
        .Y(n1981) );
  OAI2BB2XL U2214 ( .B0(n6784), .B1(n182), .A0N(\ram[87][8] ), .A1N(n6523), 
        .Y(n1982) );
  OAI2BB2XL U2215 ( .B0(n6761), .B1(n182), .A0N(\ram[87][9] ), .A1N(n6523), 
        .Y(n1983) );
  OAI2BB2XL U2216 ( .B0(n6738), .B1(n182), .A0N(\ram[87][10] ), .A1N(n6523), 
        .Y(n1984) );
  OAI2BB2XL U2217 ( .B0(n6715), .B1(n182), .A0N(\ram[87][11] ), .A1N(n6523), 
        .Y(n1985) );
  OAI2BB2XL U2218 ( .B0(n6692), .B1(n182), .A0N(\ram[87][12] ), .A1N(n6523), 
        .Y(n1986) );
  OAI2BB2XL U2219 ( .B0(n6669), .B1(n182), .A0N(\ram[87][13] ), .A1N(n6523), 
        .Y(n1987) );
  OAI2BB2XL U2220 ( .B0(n6646), .B1(n182), .A0N(\ram[87][14] ), .A1N(n6523), 
        .Y(n1988) );
  OAI2BB2XL U2221 ( .B0(n6623), .B1(n182), .A0N(\ram[87][15] ), .A1N(n6523), 
        .Y(n1989) );
  OAI2BB2XL U2222 ( .B0(n6972), .B1(n184), .A0N(\ram[88][0] ), .A1N(n6522), 
        .Y(n1990) );
  OAI2BB2XL U2223 ( .B0(n6949), .B1(n184), .A0N(\ram[88][1] ), .A1N(n6522), 
        .Y(n1991) );
  OAI2BB2XL U2224 ( .B0(n6926), .B1(n184), .A0N(\ram[88][2] ), .A1N(n6522), 
        .Y(n1992) );
  OAI2BB2XL U2225 ( .B0(n6903), .B1(n184), .A0N(\ram[88][3] ), .A1N(n6522), 
        .Y(n1993) );
  OAI2BB2XL U2226 ( .B0(n6875), .B1(n184), .A0N(\ram[88][4] ), .A1N(n6522), 
        .Y(n1994) );
  OAI2BB2XL U2227 ( .B0(n6852), .B1(n184), .A0N(\ram[88][5] ), .A1N(n6522), 
        .Y(n1995) );
  OAI2BB2XL U2228 ( .B0(n6829), .B1(n184), .A0N(\ram[88][6] ), .A1N(n6522), 
        .Y(n1996) );
  OAI2BB2XL U2229 ( .B0(n6806), .B1(n184), .A0N(\ram[88][7] ), .A1N(n6522), 
        .Y(n1997) );
  OAI2BB2XL U2230 ( .B0(n6783), .B1(n184), .A0N(\ram[88][8] ), .A1N(n6522), 
        .Y(n1998) );
  OAI2BB2XL U2231 ( .B0(n6760), .B1(n184), .A0N(\ram[88][9] ), .A1N(n6522), 
        .Y(n1999) );
  OAI2BB2XL U2232 ( .B0(n6737), .B1(n184), .A0N(\ram[88][10] ), .A1N(n6522), 
        .Y(n2000) );
  OAI2BB2XL U2233 ( .B0(n6714), .B1(n184), .A0N(\ram[88][11] ), .A1N(n6522), 
        .Y(n2001) );
  OAI2BB2XL U2234 ( .B0(n6691), .B1(n184), .A0N(\ram[88][12] ), .A1N(n6522), 
        .Y(n2002) );
  OAI2BB2XL U2235 ( .B0(n6668), .B1(n184), .A0N(\ram[88][13] ), .A1N(n6522), 
        .Y(n2003) );
  OAI2BB2XL U2236 ( .B0(n6645), .B1(n184), .A0N(\ram[88][14] ), .A1N(n6522), 
        .Y(n2004) );
  OAI2BB2XL U2237 ( .B0(n6622), .B1(n184), .A0N(\ram[88][15] ), .A1N(n6522), 
        .Y(n2005) );
  OAI2BB2XL U2238 ( .B0(n6972), .B1(n186), .A0N(\ram[89][0] ), .A1N(n6521), 
        .Y(n2006) );
  OAI2BB2XL U2239 ( .B0(n6949), .B1(n186), .A0N(\ram[89][1] ), .A1N(n6521), 
        .Y(n2007) );
  OAI2BB2XL U2240 ( .B0(n6926), .B1(n186), .A0N(\ram[89][2] ), .A1N(n6521), 
        .Y(n2008) );
  OAI2BB2XL U2241 ( .B0(n6903), .B1(n186), .A0N(\ram[89][3] ), .A1N(n6521), 
        .Y(n2009) );
  OAI2BB2XL U2242 ( .B0(n6875), .B1(n186), .A0N(\ram[89][4] ), .A1N(n6521), 
        .Y(n2010) );
  OAI2BB2XL U2243 ( .B0(n6852), .B1(n186), .A0N(\ram[89][5] ), .A1N(n6521), 
        .Y(n2011) );
  OAI2BB2XL U2244 ( .B0(n6829), .B1(n186), .A0N(\ram[89][6] ), .A1N(n6521), 
        .Y(n2012) );
  OAI2BB2XL U2245 ( .B0(n6806), .B1(n186), .A0N(\ram[89][7] ), .A1N(n6521), 
        .Y(n2013) );
  OAI2BB2XL U2246 ( .B0(n6783), .B1(n186), .A0N(\ram[89][8] ), .A1N(n6521), 
        .Y(n2014) );
  OAI2BB2XL U2247 ( .B0(n6760), .B1(n186), .A0N(\ram[89][9] ), .A1N(n6521), 
        .Y(n2015) );
  OAI2BB2XL U2248 ( .B0(n6737), .B1(n186), .A0N(\ram[89][10] ), .A1N(n6521), 
        .Y(n2016) );
  OAI2BB2XL U2249 ( .B0(n6714), .B1(n186), .A0N(\ram[89][11] ), .A1N(n6521), 
        .Y(n2017) );
  OAI2BB2XL U2250 ( .B0(n6691), .B1(n186), .A0N(\ram[89][12] ), .A1N(n6521), 
        .Y(n2018) );
  OAI2BB2XL U2251 ( .B0(n6668), .B1(n186), .A0N(\ram[89][13] ), .A1N(n6521), 
        .Y(n2019) );
  OAI2BB2XL U2252 ( .B0(n6645), .B1(n186), .A0N(\ram[89][14] ), .A1N(n6521), 
        .Y(n2020) );
  OAI2BB2XL U2253 ( .B0(n6622), .B1(n186), .A0N(\ram[89][15] ), .A1N(n6521), 
        .Y(n2021) );
  OAI2BB2XL U2254 ( .B0(n6972), .B1(n188), .A0N(\ram[90][0] ), .A1N(n6520), 
        .Y(n2022) );
  OAI2BB2XL U2255 ( .B0(n6949), .B1(n188), .A0N(\ram[90][1] ), .A1N(n6520), 
        .Y(n2023) );
  OAI2BB2XL U2256 ( .B0(n6926), .B1(n188), .A0N(\ram[90][2] ), .A1N(n6520), 
        .Y(n2024) );
  OAI2BB2XL U2257 ( .B0(n6903), .B1(n188), .A0N(\ram[90][3] ), .A1N(n6520), 
        .Y(n2025) );
  OAI2BB2XL U2258 ( .B0(n6875), .B1(n188), .A0N(\ram[90][4] ), .A1N(n6520), 
        .Y(n2026) );
  OAI2BB2XL U2259 ( .B0(n6852), .B1(n188), .A0N(\ram[90][5] ), .A1N(n6520), 
        .Y(n2027) );
  OAI2BB2XL U2260 ( .B0(n6829), .B1(n188), .A0N(\ram[90][6] ), .A1N(n6520), 
        .Y(n2028) );
  OAI2BB2XL U2261 ( .B0(n6806), .B1(n188), .A0N(\ram[90][7] ), .A1N(n6520), 
        .Y(n2029) );
  OAI2BB2XL U2262 ( .B0(n6783), .B1(n188), .A0N(\ram[90][8] ), .A1N(n6520), 
        .Y(n2030) );
  OAI2BB2XL U2263 ( .B0(n6760), .B1(n188), .A0N(\ram[90][9] ), .A1N(n6520), 
        .Y(n2031) );
  OAI2BB2XL U2264 ( .B0(n6737), .B1(n188), .A0N(\ram[90][10] ), .A1N(n6520), 
        .Y(n2032) );
  OAI2BB2XL U2265 ( .B0(n6714), .B1(n188), .A0N(\ram[90][11] ), .A1N(n6520), 
        .Y(n2033) );
  OAI2BB2XL U2266 ( .B0(n6691), .B1(n188), .A0N(\ram[90][12] ), .A1N(n6520), 
        .Y(n2034) );
  OAI2BB2XL U2267 ( .B0(n6668), .B1(n188), .A0N(\ram[90][13] ), .A1N(n6520), 
        .Y(n2035) );
  OAI2BB2XL U2268 ( .B0(n6645), .B1(n188), .A0N(\ram[90][14] ), .A1N(n6520), 
        .Y(n2036) );
  OAI2BB2XL U2269 ( .B0(n6622), .B1(n188), .A0N(\ram[90][15] ), .A1N(n6520), 
        .Y(n2037) );
  OAI2BB2XL U2270 ( .B0(n6972), .B1(n190), .A0N(\ram[91][0] ), .A1N(n6519), 
        .Y(n2038) );
  OAI2BB2XL U2271 ( .B0(n6949), .B1(n190), .A0N(\ram[91][1] ), .A1N(n6519), 
        .Y(n2039) );
  OAI2BB2XL U2272 ( .B0(n6926), .B1(n190), .A0N(\ram[91][2] ), .A1N(n6519), 
        .Y(n2040) );
  OAI2BB2XL U2273 ( .B0(n6903), .B1(n190), .A0N(\ram[91][3] ), .A1N(n6519), 
        .Y(n2041) );
  OAI2BB2XL U2274 ( .B0(n6875), .B1(n190), .A0N(\ram[91][4] ), .A1N(n6519), 
        .Y(n2042) );
  OAI2BB2XL U2275 ( .B0(n6852), .B1(n190), .A0N(\ram[91][5] ), .A1N(n6519), 
        .Y(n2043) );
  OAI2BB2XL U2276 ( .B0(n6829), .B1(n190), .A0N(\ram[91][6] ), .A1N(n6519), 
        .Y(n2044) );
  OAI2BB2XL U2277 ( .B0(n6806), .B1(n190), .A0N(\ram[91][7] ), .A1N(n6519), 
        .Y(n2045) );
  OAI2BB2XL U2278 ( .B0(n6783), .B1(n190), .A0N(\ram[91][8] ), .A1N(n6519), 
        .Y(n2046) );
  OAI2BB2XL U2279 ( .B0(n6760), .B1(n190), .A0N(\ram[91][9] ), .A1N(n6519), 
        .Y(n2047) );
  OAI2BB2XL U2280 ( .B0(n6737), .B1(n190), .A0N(\ram[91][10] ), .A1N(n6519), 
        .Y(n2048) );
  OAI2BB2XL U2281 ( .B0(n6714), .B1(n190), .A0N(\ram[91][11] ), .A1N(n6519), 
        .Y(n2049) );
  OAI2BB2XL U2282 ( .B0(n6691), .B1(n190), .A0N(\ram[91][12] ), .A1N(n6519), 
        .Y(n2050) );
  OAI2BB2XL U2283 ( .B0(n6668), .B1(n190), .A0N(\ram[91][13] ), .A1N(n6519), 
        .Y(n2051) );
  OAI2BB2XL U2284 ( .B0(n6645), .B1(n190), .A0N(\ram[91][14] ), .A1N(n6519), 
        .Y(n2052) );
  OAI2BB2XL U2285 ( .B0(n6622), .B1(n190), .A0N(\ram[91][15] ), .A1N(n6519), 
        .Y(n2053) );
  OAI2BB2XL U2286 ( .B0(n6972), .B1(n192), .A0N(\ram[92][0] ), .A1N(n6518), 
        .Y(n2054) );
  OAI2BB2XL U2287 ( .B0(n6949), .B1(n192), .A0N(\ram[92][1] ), .A1N(n6518), 
        .Y(n2055) );
  OAI2BB2XL U2288 ( .B0(n6926), .B1(n192), .A0N(\ram[92][2] ), .A1N(n6518), 
        .Y(n2056) );
  OAI2BB2XL U2289 ( .B0(n6903), .B1(n192), .A0N(\ram[92][3] ), .A1N(n6518), 
        .Y(n2057) );
  OAI2BB2XL U2290 ( .B0(n6875), .B1(n192), .A0N(\ram[92][4] ), .A1N(n6518), 
        .Y(n2058) );
  OAI2BB2XL U2291 ( .B0(n6852), .B1(n192), .A0N(\ram[92][5] ), .A1N(n6518), 
        .Y(n2059) );
  OAI2BB2XL U2292 ( .B0(n6829), .B1(n192), .A0N(\ram[92][6] ), .A1N(n6518), 
        .Y(n2060) );
  OAI2BB2XL U2293 ( .B0(n6806), .B1(n192), .A0N(\ram[92][7] ), .A1N(n6518), 
        .Y(n2061) );
  OAI2BB2XL U2294 ( .B0(n6783), .B1(n192), .A0N(\ram[92][8] ), .A1N(n6518), 
        .Y(n2062) );
  OAI2BB2XL U2295 ( .B0(n6760), .B1(n192), .A0N(\ram[92][9] ), .A1N(n6518), 
        .Y(n2063) );
  OAI2BB2XL U2296 ( .B0(n6737), .B1(n192), .A0N(\ram[92][10] ), .A1N(n6518), 
        .Y(n2064) );
  OAI2BB2XL U2297 ( .B0(n6714), .B1(n192), .A0N(\ram[92][11] ), .A1N(n6518), 
        .Y(n2065) );
  OAI2BB2XL U2298 ( .B0(n6691), .B1(n192), .A0N(\ram[92][12] ), .A1N(n6518), 
        .Y(n2066) );
  OAI2BB2XL U2299 ( .B0(n6668), .B1(n192), .A0N(\ram[92][13] ), .A1N(n6518), 
        .Y(n2067) );
  OAI2BB2XL U2300 ( .B0(n6645), .B1(n192), .A0N(\ram[92][14] ), .A1N(n6518), 
        .Y(n2068) );
  OAI2BB2XL U2301 ( .B0(n6622), .B1(n192), .A0N(\ram[92][15] ), .A1N(n6518), 
        .Y(n2069) );
  OAI2BB2XL U2302 ( .B0(n6972), .B1(n194), .A0N(\ram[93][0] ), .A1N(n6517), 
        .Y(n2070) );
  OAI2BB2XL U2303 ( .B0(n6949), .B1(n194), .A0N(\ram[93][1] ), .A1N(n6517), 
        .Y(n2071) );
  OAI2BB2XL U2304 ( .B0(n6926), .B1(n194), .A0N(\ram[93][2] ), .A1N(n6517), 
        .Y(n2072) );
  OAI2BB2XL U2305 ( .B0(n6903), .B1(n194), .A0N(\ram[93][3] ), .A1N(n6517), 
        .Y(n2073) );
  OAI2BB2XL U2306 ( .B0(n6875), .B1(n194), .A0N(\ram[93][4] ), .A1N(n6517), 
        .Y(n2074) );
  OAI2BB2XL U2307 ( .B0(n6852), .B1(n194), .A0N(\ram[93][5] ), .A1N(n6517), 
        .Y(n2075) );
  OAI2BB2XL U2308 ( .B0(n6829), .B1(n194), .A0N(\ram[93][6] ), .A1N(n6517), 
        .Y(n2076) );
  OAI2BB2XL U2309 ( .B0(n6806), .B1(n194), .A0N(\ram[93][7] ), .A1N(n6517), 
        .Y(n2077) );
  OAI2BB2XL U2310 ( .B0(n6783), .B1(n194), .A0N(\ram[93][8] ), .A1N(n6517), 
        .Y(n2078) );
  OAI2BB2XL U2311 ( .B0(n6760), .B1(n194), .A0N(\ram[93][9] ), .A1N(n6517), 
        .Y(n2079) );
  OAI2BB2XL U2312 ( .B0(n6737), .B1(n194), .A0N(\ram[93][10] ), .A1N(n6517), 
        .Y(n2080) );
  OAI2BB2XL U2313 ( .B0(n6714), .B1(n194), .A0N(\ram[93][11] ), .A1N(n6517), 
        .Y(n2081) );
  OAI2BB2XL U2314 ( .B0(n6691), .B1(n194), .A0N(\ram[93][12] ), .A1N(n6517), 
        .Y(n2082) );
  OAI2BB2XL U2315 ( .B0(n6668), .B1(n194), .A0N(\ram[93][13] ), .A1N(n6517), 
        .Y(n2083) );
  OAI2BB2XL U2316 ( .B0(n6645), .B1(n194), .A0N(\ram[93][14] ), .A1N(n6517), 
        .Y(n2084) );
  OAI2BB2XL U2317 ( .B0(n6622), .B1(n194), .A0N(\ram[93][15] ), .A1N(n6517), 
        .Y(n2085) );
  OAI2BB2XL U2318 ( .B0(n6972), .B1(n196), .A0N(\ram[94][0] ), .A1N(n6516), 
        .Y(n2086) );
  OAI2BB2XL U2319 ( .B0(n6949), .B1(n196), .A0N(\ram[94][1] ), .A1N(n6516), 
        .Y(n2087) );
  OAI2BB2XL U2320 ( .B0(n6926), .B1(n196), .A0N(\ram[94][2] ), .A1N(n6516), 
        .Y(n2088) );
  OAI2BB2XL U2321 ( .B0(n6903), .B1(n196), .A0N(\ram[94][3] ), .A1N(n6516), 
        .Y(n2089) );
  OAI2BB2XL U2322 ( .B0(n6875), .B1(n196), .A0N(\ram[94][4] ), .A1N(n6516), 
        .Y(n2090) );
  OAI2BB2XL U2323 ( .B0(n6852), .B1(n196), .A0N(\ram[94][5] ), .A1N(n6516), 
        .Y(n2091) );
  OAI2BB2XL U2324 ( .B0(n6829), .B1(n196), .A0N(\ram[94][6] ), .A1N(n6516), 
        .Y(n2092) );
  OAI2BB2XL U2325 ( .B0(n6806), .B1(n196), .A0N(\ram[94][7] ), .A1N(n6516), 
        .Y(n2093) );
  OAI2BB2XL U2326 ( .B0(n6783), .B1(n196), .A0N(\ram[94][8] ), .A1N(n6516), 
        .Y(n2094) );
  OAI2BB2XL U2327 ( .B0(n6760), .B1(n196), .A0N(\ram[94][9] ), .A1N(n6516), 
        .Y(n2095) );
  OAI2BB2XL U2328 ( .B0(n6737), .B1(n196), .A0N(\ram[94][10] ), .A1N(n6516), 
        .Y(n2096) );
  OAI2BB2XL U2329 ( .B0(n6714), .B1(n196), .A0N(\ram[94][11] ), .A1N(n6516), 
        .Y(n2097) );
  OAI2BB2XL U2330 ( .B0(n6691), .B1(n196), .A0N(\ram[94][12] ), .A1N(n6516), 
        .Y(n2098) );
  OAI2BB2XL U2331 ( .B0(n6668), .B1(n196), .A0N(\ram[94][13] ), .A1N(n6516), 
        .Y(n2099) );
  OAI2BB2XL U2332 ( .B0(n6645), .B1(n196), .A0N(\ram[94][14] ), .A1N(n6516), 
        .Y(n2100) );
  OAI2BB2XL U2333 ( .B0(n6622), .B1(n196), .A0N(\ram[94][15] ), .A1N(n6516), 
        .Y(n2101) );
  OAI2BB2XL U2334 ( .B0(n6972), .B1(n198), .A0N(\ram[95][0] ), .A1N(n6515), 
        .Y(n2102) );
  OAI2BB2XL U2335 ( .B0(n6949), .B1(n198), .A0N(\ram[95][1] ), .A1N(n6515), 
        .Y(n2103) );
  OAI2BB2XL U2336 ( .B0(n6926), .B1(n198), .A0N(\ram[95][2] ), .A1N(n6515), 
        .Y(n2104) );
  OAI2BB2XL U2337 ( .B0(n6903), .B1(n198), .A0N(\ram[95][3] ), .A1N(n6515), 
        .Y(n2105) );
  OAI2BB2XL U2338 ( .B0(n6875), .B1(n198), .A0N(\ram[95][4] ), .A1N(n6515), 
        .Y(n2106) );
  OAI2BB2XL U2339 ( .B0(n6852), .B1(n198), .A0N(\ram[95][5] ), .A1N(n6515), 
        .Y(n2107) );
  OAI2BB2XL U2340 ( .B0(n6829), .B1(n198), .A0N(\ram[95][6] ), .A1N(n6515), 
        .Y(n2108) );
  OAI2BB2XL U2341 ( .B0(n6806), .B1(n198), .A0N(\ram[95][7] ), .A1N(n6515), 
        .Y(n2109) );
  OAI2BB2XL U2342 ( .B0(n6783), .B1(n198), .A0N(\ram[95][8] ), .A1N(n6515), 
        .Y(n2110) );
  OAI2BB2XL U2343 ( .B0(n6760), .B1(n198), .A0N(\ram[95][9] ), .A1N(n6515), 
        .Y(n2111) );
  OAI2BB2XL U2344 ( .B0(n6737), .B1(n198), .A0N(\ram[95][10] ), .A1N(n6515), 
        .Y(n2112) );
  OAI2BB2XL U2345 ( .B0(n6714), .B1(n198), .A0N(\ram[95][11] ), .A1N(n6515), 
        .Y(n2113) );
  OAI2BB2XL U2346 ( .B0(n6691), .B1(n198), .A0N(\ram[95][12] ), .A1N(n6515), 
        .Y(n2114) );
  OAI2BB2XL U2347 ( .B0(n6668), .B1(n198), .A0N(\ram[95][13] ), .A1N(n6515), 
        .Y(n2115) );
  OAI2BB2XL U2348 ( .B0(n6645), .B1(n198), .A0N(\ram[95][14] ), .A1N(n6515), 
        .Y(n2116) );
  OAI2BB2XL U2349 ( .B0(n6622), .B1(n198), .A0N(\ram[95][15] ), .A1N(n6515), 
        .Y(n2117) );
  OAI2BB2XL U2350 ( .B0(n6972), .B1(n200), .A0N(\ram[96][0] ), .A1N(n6514), 
        .Y(n2118) );
  OAI2BB2XL U2351 ( .B0(n6949), .B1(n200), .A0N(\ram[96][1] ), .A1N(n6514), 
        .Y(n2119) );
  OAI2BB2XL U2352 ( .B0(n6926), .B1(n200), .A0N(\ram[96][2] ), .A1N(n6514), 
        .Y(n2120) );
  OAI2BB2XL U2353 ( .B0(n6903), .B1(n200), .A0N(\ram[96][3] ), .A1N(n6514), 
        .Y(n2121) );
  OAI2BB2XL U2354 ( .B0(n6875), .B1(n200), .A0N(\ram[96][4] ), .A1N(n6514), 
        .Y(n2122) );
  OAI2BB2XL U2355 ( .B0(n6852), .B1(n200), .A0N(\ram[96][5] ), .A1N(n6514), 
        .Y(n2123) );
  OAI2BB2XL U2356 ( .B0(n6829), .B1(n200), .A0N(\ram[96][6] ), .A1N(n6514), 
        .Y(n2124) );
  OAI2BB2XL U2357 ( .B0(n6806), .B1(n200), .A0N(\ram[96][7] ), .A1N(n6514), 
        .Y(n2125) );
  OAI2BB2XL U2358 ( .B0(n6783), .B1(n200), .A0N(\ram[96][8] ), .A1N(n6514), 
        .Y(n2126) );
  OAI2BB2XL U2359 ( .B0(n6760), .B1(n200), .A0N(\ram[96][9] ), .A1N(n6514), 
        .Y(n2127) );
  OAI2BB2XL U2360 ( .B0(n6737), .B1(n200), .A0N(\ram[96][10] ), .A1N(n6514), 
        .Y(n2128) );
  OAI2BB2XL U2361 ( .B0(n6714), .B1(n200), .A0N(\ram[96][11] ), .A1N(n6514), 
        .Y(n2129) );
  OAI2BB2XL U2362 ( .B0(n6691), .B1(n200), .A0N(\ram[96][12] ), .A1N(n6514), 
        .Y(n2130) );
  OAI2BB2XL U2363 ( .B0(n6668), .B1(n200), .A0N(\ram[96][13] ), .A1N(n6514), 
        .Y(n2131) );
  OAI2BB2XL U2364 ( .B0(n6645), .B1(n200), .A0N(\ram[96][14] ), .A1N(n6514), 
        .Y(n2132) );
  OAI2BB2XL U2365 ( .B0(n6622), .B1(n200), .A0N(\ram[96][15] ), .A1N(n6514), 
        .Y(n2133) );
  OAI2BB2XL U2366 ( .B0(n6972), .B1(n202), .A0N(\ram[97][0] ), .A1N(n6513), 
        .Y(n2134) );
  OAI2BB2XL U2367 ( .B0(n6949), .B1(n202), .A0N(\ram[97][1] ), .A1N(n6513), 
        .Y(n2135) );
  OAI2BB2XL U2368 ( .B0(n6926), .B1(n202), .A0N(\ram[97][2] ), .A1N(n6513), 
        .Y(n2136) );
  OAI2BB2XL U2369 ( .B0(n6903), .B1(n202), .A0N(\ram[97][3] ), .A1N(n6513), 
        .Y(n2137) );
  OAI2BB2XL U2370 ( .B0(n6875), .B1(n202), .A0N(\ram[97][4] ), .A1N(n6513), 
        .Y(n2138) );
  OAI2BB2XL U2371 ( .B0(n6852), .B1(n202), .A0N(\ram[97][5] ), .A1N(n6513), 
        .Y(n2139) );
  OAI2BB2XL U2372 ( .B0(n6829), .B1(n202), .A0N(\ram[97][6] ), .A1N(n6513), 
        .Y(n2140) );
  OAI2BB2XL U2373 ( .B0(n6806), .B1(n202), .A0N(\ram[97][7] ), .A1N(n6513), 
        .Y(n2141) );
  OAI2BB2XL U2374 ( .B0(n6783), .B1(n202), .A0N(\ram[97][8] ), .A1N(n6513), 
        .Y(n2142) );
  OAI2BB2XL U2375 ( .B0(n6760), .B1(n202), .A0N(\ram[97][9] ), .A1N(n6513), 
        .Y(n2143) );
  OAI2BB2XL U2376 ( .B0(n6737), .B1(n202), .A0N(\ram[97][10] ), .A1N(n6513), 
        .Y(n2144) );
  OAI2BB2XL U2377 ( .B0(n6714), .B1(n202), .A0N(\ram[97][11] ), .A1N(n6513), 
        .Y(n2145) );
  OAI2BB2XL U2378 ( .B0(n6691), .B1(n202), .A0N(\ram[97][12] ), .A1N(n6513), 
        .Y(n2146) );
  OAI2BB2XL U2379 ( .B0(n6668), .B1(n202), .A0N(\ram[97][13] ), .A1N(n6513), 
        .Y(n2147) );
  OAI2BB2XL U2380 ( .B0(n6645), .B1(n202), .A0N(\ram[97][14] ), .A1N(n6513), 
        .Y(n2148) );
  OAI2BB2XL U2381 ( .B0(n6622), .B1(n202), .A0N(\ram[97][15] ), .A1N(n6513), 
        .Y(n2149) );
  OAI2BB2XL U2382 ( .B0(n6972), .B1(n204), .A0N(\ram[98][0] ), .A1N(n6512), 
        .Y(n2150) );
  OAI2BB2XL U2383 ( .B0(n6949), .B1(n204), .A0N(\ram[98][1] ), .A1N(n6512), 
        .Y(n2151) );
  OAI2BB2XL U2384 ( .B0(n6926), .B1(n204), .A0N(\ram[98][2] ), .A1N(n6512), 
        .Y(n2152) );
  OAI2BB2XL U2385 ( .B0(n6903), .B1(n204), .A0N(\ram[98][3] ), .A1N(n6512), 
        .Y(n2153) );
  OAI2BB2XL U2386 ( .B0(n6875), .B1(n204), .A0N(\ram[98][4] ), .A1N(n6512), 
        .Y(n2154) );
  OAI2BB2XL U2387 ( .B0(n6852), .B1(n204), .A0N(\ram[98][5] ), .A1N(n6512), 
        .Y(n2155) );
  OAI2BB2XL U2388 ( .B0(n6829), .B1(n204), .A0N(\ram[98][6] ), .A1N(n6512), 
        .Y(n2156) );
  OAI2BB2XL U2389 ( .B0(n6806), .B1(n204), .A0N(\ram[98][7] ), .A1N(n6512), 
        .Y(n2157) );
  OAI2BB2XL U2390 ( .B0(n6783), .B1(n204), .A0N(\ram[98][8] ), .A1N(n6512), 
        .Y(n2158) );
  OAI2BB2XL U2391 ( .B0(n6760), .B1(n204), .A0N(\ram[98][9] ), .A1N(n6512), 
        .Y(n2159) );
  OAI2BB2XL U2392 ( .B0(n6737), .B1(n204), .A0N(\ram[98][10] ), .A1N(n6512), 
        .Y(n2160) );
  OAI2BB2XL U2393 ( .B0(n6714), .B1(n204), .A0N(\ram[98][11] ), .A1N(n6512), 
        .Y(n2161) );
  OAI2BB2XL U2394 ( .B0(n6691), .B1(n204), .A0N(\ram[98][12] ), .A1N(n6512), 
        .Y(n2162) );
  OAI2BB2XL U2395 ( .B0(n6668), .B1(n204), .A0N(\ram[98][13] ), .A1N(n6512), 
        .Y(n2163) );
  OAI2BB2XL U2396 ( .B0(n6645), .B1(n204), .A0N(\ram[98][14] ), .A1N(n6512), 
        .Y(n2164) );
  OAI2BB2XL U2397 ( .B0(n6622), .B1(n204), .A0N(\ram[98][15] ), .A1N(n6512), 
        .Y(n2165) );
  OAI2BB2XL U2398 ( .B0(n6972), .B1(n206), .A0N(\ram[99][0] ), .A1N(n6511), 
        .Y(n2166) );
  OAI2BB2XL U2399 ( .B0(n6949), .B1(n206), .A0N(\ram[99][1] ), .A1N(n6511), 
        .Y(n2167) );
  OAI2BB2XL U2400 ( .B0(n6926), .B1(n206), .A0N(\ram[99][2] ), .A1N(n6511), 
        .Y(n2168) );
  OAI2BB2XL U2401 ( .B0(n6903), .B1(n206), .A0N(\ram[99][3] ), .A1N(n6511), 
        .Y(n2169) );
  OAI2BB2XL U2402 ( .B0(n6875), .B1(n206), .A0N(\ram[99][4] ), .A1N(n6511), 
        .Y(n2170) );
  OAI2BB2XL U2403 ( .B0(n6852), .B1(n206), .A0N(\ram[99][5] ), .A1N(n6511), 
        .Y(n2171) );
  OAI2BB2XL U2404 ( .B0(n6829), .B1(n206), .A0N(\ram[99][6] ), .A1N(n6511), 
        .Y(n2172) );
  OAI2BB2XL U2405 ( .B0(n6806), .B1(n206), .A0N(\ram[99][7] ), .A1N(n6511), 
        .Y(n2173) );
  OAI2BB2XL U2406 ( .B0(n6783), .B1(n206), .A0N(\ram[99][8] ), .A1N(n6511), 
        .Y(n2174) );
  OAI2BB2XL U2407 ( .B0(n6760), .B1(n206), .A0N(\ram[99][9] ), .A1N(n6511), 
        .Y(n2175) );
  OAI2BB2XL U2408 ( .B0(n6737), .B1(n206), .A0N(\ram[99][10] ), .A1N(n6511), 
        .Y(n2176) );
  OAI2BB2XL U2409 ( .B0(n6714), .B1(n206), .A0N(\ram[99][11] ), .A1N(n6511), 
        .Y(n2177) );
  OAI2BB2XL U2410 ( .B0(n6691), .B1(n206), .A0N(\ram[99][12] ), .A1N(n6511), 
        .Y(n2178) );
  OAI2BB2XL U2411 ( .B0(n6668), .B1(n206), .A0N(\ram[99][13] ), .A1N(n6511), 
        .Y(n2179) );
  OAI2BB2XL U2412 ( .B0(n6645), .B1(n206), .A0N(\ram[99][14] ), .A1N(n6511), 
        .Y(n2180) );
  OAI2BB2XL U2413 ( .B0(n6622), .B1(n206), .A0N(\ram[99][15] ), .A1N(n6511), 
        .Y(n2181) );
  OAI2BB2XL U2414 ( .B0(n6971), .B1(n209), .A0N(\ram[100][0] ), .A1N(n6510), 
        .Y(n2182) );
  OAI2BB2XL U2415 ( .B0(n6948), .B1(n209), .A0N(\ram[100][1] ), .A1N(n6510), 
        .Y(n2183) );
  OAI2BB2XL U2416 ( .B0(n6925), .B1(n209), .A0N(\ram[100][2] ), .A1N(n6510), 
        .Y(n2184) );
  OAI2BB2XL U2417 ( .B0(n6902), .B1(n209), .A0N(\ram[100][3] ), .A1N(n6510), 
        .Y(n2185) );
  OAI2BB2XL U2418 ( .B0(n6874), .B1(n209), .A0N(\ram[100][4] ), .A1N(n6510), 
        .Y(n2186) );
  OAI2BB2XL U2419 ( .B0(n6851), .B1(n209), .A0N(\ram[100][5] ), .A1N(n6510), 
        .Y(n2187) );
  OAI2BB2XL U2420 ( .B0(n6828), .B1(n209), .A0N(\ram[100][6] ), .A1N(n6510), 
        .Y(n2188) );
  OAI2BB2XL U2421 ( .B0(n6805), .B1(n209), .A0N(\ram[100][7] ), .A1N(n6510), 
        .Y(n2189) );
  OAI2BB2XL U2422 ( .B0(n6782), .B1(n209), .A0N(\ram[100][8] ), .A1N(n6510), 
        .Y(n2190) );
  OAI2BB2XL U2423 ( .B0(n6759), .B1(n209), .A0N(\ram[100][9] ), .A1N(n6510), 
        .Y(n2191) );
  OAI2BB2XL U2424 ( .B0(n6736), .B1(n209), .A0N(\ram[100][10] ), .A1N(n6510), 
        .Y(n2192) );
  OAI2BB2XL U2425 ( .B0(n6713), .B1(n209), .A0N(\ram[100][11] ), .A1N(n6510), 
        .Y(n2193) );
  OAI2BB2XL U2426 ( .B0(n6690), .B1(n209), .A0N(\ram[100][12] ), .A1N(n6510), 
        .Y(n2194) );
  OAI2BB2XL U2427 ( .B0(n6667), .B1(n209), .A0N(\ram[100][13] ), .A1N(n6510), 
        .Y(n2195) );
  OAI2BB2XL U2428 ( .B0(n6644), .B1(n209), .A0N(\ram[100][14] ), .A1N(n6510), 
        .Y(n2196) );
  OAI2BB2XL U2429 ( .B0(n6621), .B1(n209), .A0N(\ram[100][15] ), .A1N(n6510), 
        .Y(n2197) );
  OAI2BB2XL U2430 ( .B0(n6971), .B1(n211), .A0N(\ram[101][0] ), .A1N(n6509), 
        .Y(n2198) );
  OAI2BB2XL U2431 ( .B0(n6948), .B1(n211), .A0N(\ram[101][1] ), .A1N(n6509), 
        .Y(n2199) );
  OAI2BB2XL U2432 ( .B0(n6925), .B1(n211), .A0N(\ram[101][2] ), .A1N(n6509), 
        .Y(n2200) );
  OAI2BB2XL U2433 ( .B0(n6902), .B1(n211), .A0N(\ram[101][3] ), .A1N(n6509), 
        .Y(n2201) );
  OAI2BB2XL U2434 ( .B0(n6874), .B1(n211), .A0N(\ram[101][4] ), .A1N(n6509), 
        .Y(n2202) );
  OAI2BB2XL U2435 ( .B0(n6851), .B1(n211), .A0N(\ram[101][5] ), .A1N(n6509), 
        .Y(n2203) );
  OAI2BB2XL U2436 ( .B0(n6828), .B1(n211), .A0N(\ram[101][6] ), .A1N(n6509), 
        .Y(n2204) );
  OAI2BB2XL U2437 ( .B0(n6805), .B1(n211), .A0N(\ram[101][7] ), .A1N(n6509), 
        .Y(n2205) );
  OAI2BB2XL U2438 ( .B0(n6782), .B1(n211), .A0N(\ram[101][8] ), .A1N(n6509), 
        .Y(n2206) );
  OAI2BB2XL U2439 ( .B0(n6759), .B1(n211), .A0N(\ram[101][9] ), .A1N(n6509), 
        .Y(n2207) );
  OAI2BB2XL U2440 ( .B0(n6736), .B1(n211), .A0N(\ram[101][10] ), .A1N(n6509), 
        .Y(n2208) );
  OAI2BB2XL U2441 ( .B0(n6713), .B1(n211), .A0N(\ram[101][11] ), .A1N(n6509), 
        .Y(n2209) );
  OAI2BB2XL U2442 ( .B0(n6690), .B1(n211), .A0N(\ram[101][12] ), .A1N(n6509), 
        .Y(n2210) );
  OAI2BB2XL U2443 ( .B0(n6667), .B1(n211), .A0N(\ram[101][13] ), .A1N(n6509), 
        .Y(n2211) );
  OAI2BB2XL U2444 ( .B0(n6644), .B1(n211), .A0N(\ram[101][14] ), .A1N(n6509), 
        .Y(n2212) );
  OAI2BB2XL U2445 ( .B0(n6621), .B1(n211), .A0N(\ram[101][15] ), .A1N(n6509), 
        .Y(n2213) );
  OAI2BB2XL U2446 ( .B0(n6971), .B1(n212), .A0N(\ram[102][0] ), .A1N(n6508), 
        .Y(n2214) );
  OAI2BB2XL U2447 ( .B0(n6948), .B1(n212), .A0N(\ram[102][1] ), .A1N(n6508), 
        .Y(n2215) );
  OAI2BB2XL U2448 ( .B0(n6925), .B1(n212), .A0N(\ram[102][2] ), .A1N(n6508), 
        .Y(n2216) );
  OAI2BB2XL U2449 ( .B0(n6902), .B1(n212), .A0N(\ram[102][3] ), .A1N(n6508), 
        .Y(n2217) );
  OAI2BB2XL U2450 ( .B0(n6874), .B1(n212), .A0N(\ram[102][4] ), .A1N(n6508), 
        .Y(n2218) );
  OAI2BB2XL U2451 ( .B0(n6851), .B1(n212), .A0N(\ram[102][5] ), .A1N(n6508), 
        .Y(n2219) );
  OAI2BB2XL U2452 ( .B0(n6828), .B1(n212), .A0N(\ram[102][6] ), .A1N(n6508), 
        .Y(n2220) );
  OAI2BB2XL U2453 ( .B0(n6805), .B1(n212), .A0N(\ram[102][7] ), .A1N(n6508), 
        .Y(n2221) );
  OAI2BB2XL U2454 ( .B0(n6782), .B1(n212), .A0N(\ram[102][8] ), .A1N(n6508), 
        .Y(n2222) );
  OAI2BB2XL U2455 ( .B0(n6759), .B1(n212), .A0N(\ram[102][9] ), .A1N(n6508), 
        .Y(n2223) );
  OAI2BB2XL U2456 ( .B0(n6736), .B1(n212), .A0N(\ram[102][10] ), .A1N(n6508), 
        .Y(n2224) );
  OAI2BB2XL U2457 ( .B0(n6713), .B1(n212), .A0N(\ram[102][11] ), .A1N(n6508), 
        .Y(n2225) );
  OAI2BB2XL U2458 ( .B0(n6690), .B1(n212), .A0N(\ram[102][12] ), .A1N(n6508), 
        .Y(n2226) );
  OAI2BB2XL U2459 ( .B0(n6667), .B1(n212), .A0N(\ram[102][13] ), .A1N(n6508), 
        .Y(n2227) );
  OAI2BB2XL U2460 ( .B0(n6644), .B1(n212), .A0N(\ram[102][14] ), .A1N(n6508), 
        .Y(n2228) );
  OAI2BB2XL U2461 ( .B0(n6621), .B1(n212), .A0N(\ram[102][15] ), .A1N(n6508), 
        .Y(n2229) );
  OAI2BB2XL U2462 ( .B0(n6971), .B1(n214), .A0N(\ram[103][0] ), .A1N(n6507), 
        .Y(n2230) );
  OAI2BB2XL U2463 ( .B0(n6948), .B1(n214), .A0N(\ram[103][1] ), .A1N(n6507), 
        .Y(n2231) );
  OAI2BB2XL U2464 ( .B0(n6925), .B1(n214), .A0N(\ram[103][2] ), .A1N(n6507), 
        .Y(n2232) );
  OAI2BB2XL U2465 ( .B0(n6902), .B1(n214), .A0N(\ram[103][3] ), .A1N(n6507), 
        .Y(n2233) );
  OAI2BB2XL U2466 ( .B0(n6874), .B1(n214), .A0N(\ram[103][4] ), .A1N(n6507), 
        .Y(n2234) );
  OAI2BB2XL U2467 ( .B0(n6851), .B1(n214), .A0N(\ram[103][5] ), .A1N(n6507), 
        .Y(n2235) );
  OAI2BB2XL U2468 ( .B0(n6828), .B1(n214), .A0N(\ram[103][6] ), .A1N(n6507), 
        .Y(n2236) );
  OAI2BB2XL U2469 ( .B0(n6805), .B1(n214), .A0N(\ram[103][7] ), .A1N(n6507), 
        .Y(n2237) );
  OAI2BB2XL U2470 ( .B0(n6782), .B1(n214), .A0N(\ram[103][8] ), .A1N(n6507), 
        .Y(n2238) );
  OAI2BB2XL U2471 ( .B0(n6759), .B1(n214), .A0N(\ram[103][9] ), .A1N(n6507), 
        .Y(n2239) );
  OAI2BB2XL U2472 ( .B0(n6736), .B1(n214), .A0N(\ram[103][10] ), .A1N(n6507), 
        .Y(n2240) );
  OAI2BB2XL U2473 ( .B0(n6713), .B1(n214), .A0N(\ram[103][11] ), .A1N(n6507), 
        .Y(n2241) );
  OAI2BB2XL U2474 ( .B0(n6690), .B1(n214), .A0N(\ram[103][12] ), .A1N(n6507), 
        .Y(n2242) );
  OAI2BB2XL U2475 ( .B0(n6667), .B1(n214), .A0N(\ram[103][13] ), .A1N(n6507), 
        .Y(n2243) );
  OAI2BB2XL U2476 ( .B0(n6644), .B1(n214), .A0N(\ram[103][14] ), .A1N(n6507), 
        .Y(n2244) );
  OAI2BB2XL U2477 ( .B0(n6621), .B1(n214), .A0N(\ram[103][15] ), .A1N(n6507), 
        .Y(n2245) );
  OAI2BB2XL U2478 ( .B0(n6971), .B1(n216), .A0N(\ram[104][0] ), .A1N(n6506), 
        .Y(n2246) );
  OAI2BB2XL U2479 ( .B0(n6948), .B1(n216), .A0N(\ram[104][1] ), .A1N(n6506), 
        .Y(n2247) );
  OAI2BB2XL U2480 ( .B0(n6925), .B1(n216), .A0N(\ram[104][2] ), .A1N(n6506), 
        .Y(n2248) );
  OAI2BB2XL U2481 ( .B0(n6902), .B1(n216), .A0N(\ram[104][3] ), .A1N(n6506), 
        .Y(n2249) );
  OAI2BB2XL U2482 ( .B0(n6874), .B1(n216), .A0N(\ram[104][4] ), .A1N(n6506), 
        .Y(n2250) );
  OAI2BB2XL U2483 ( .B0(n6851), .B1(n216), .A0N(\ram[104][5] ), .A1N(n6506), 
        .Y(n2251) );
  OAI2BB2XL U2484 ( .B0(n6828), .B1(n216), .A0N(\ram[104][6] ), .A1N(n6506), 
        .Y(n2252) );
  OAI2BB2XL U2485 ( .B0(n6805), .B1(n216), .A0N(\ram[104][7] ), .A1N(n6506), 
        .Y(n2253) );
  OAI2BB2XL U2486 ( .B0(n6782), .B1(n216), .A0N(\ram[104][8] ), .A1N(n6506), 
        .Y(n2254) );
  OAI2BB2XL U2487 ( .B0(n6759), .B1(n216), .A0N(\ram[104][9] ), .A1N(n6506), 
        .Y(n2255) );
  OAI2BB2XL U2488 ( .B0(n6736), .B1(n216), .A0N(\ram[104][10] ), .A1N(n6506), 
        .Y(n2256) );
  OAI2BB2XL U2489 ( .B0(n6713), .B1(n216), .A0N(\ram[104][11] ), .A1N(n6506), 
        .Y(n2257) );
  OAI2BB2XL U2490 ( .B0(n6690), .B1(n216), .A0N(\ram[104][12] ), .A1N(n6506), 
        .Y(n2258) );
  OAI2BB2XL U2491 ( .B0(n6667), .B1(n216), .A0N(\ram[104][13] ), .A1N(n6506), 
        .Y(n2259) );
  OAI2BB2XL U2492 ( .B0(n6644), .B1(n216), .A0N(\ram[104][14] ), .A1N(n6506), 
        .Y(n2260) );
  OAI2BB2XL U2493 ( .B0(n6621), .B1(n216), .A0N(\ram[104][15] ), .A1N(n6506), 
        .Y(n2261) );
  OAI2BB2XL U2494 ( .B0(n6971), .B1(n218), .A0N(\ram[105][0] ), .A1N(n6505), 
        .Y(n2262) );
  OAI2BB2XL U2495 ( .B0(n6948), .B1(n218), .A0N(\ram[105][1] ), .A1N(n6505), 
        .Y(n2263) );
  OAI2BB2XL U2496 ( .B0(n6925), .B1(n218), .A0N(\ram[105][2] ), .A1N(n6505), 
        .Y(n2264) );
  OAI2BB2XL U2497 ( .B0(n6902), .B1(n218), .A0N(\ram[105][3] ), .A1N(n6505), 
        .Y(n2265) );
  OAI2BB2XL U2498 ( .B0(n6874), .B1(n218), .A0N(\ram[105][4] ), .A1N(n6505), 
        .Y(n2266) );
  OAI2BB2XL U2499 ( .B0(n6851), .B1(n218), .A0N(\ram[105][5] ), .A1N(n6505), 
        .Y(n2267) );
  OAI2BB2XL U2500 ( .B0(n6828), .B1(n218), .A0N(\ram[105][6] ), .A1N(n6505), 
        .Y(n2268) );
  OAI2BB2XL U2501 ( .B0(n6805), .B1(n218), .A0N(\ram[105][7] ), .A1N(n6505), 
        .Y(n2269) );
  OAI2BB2XL U2502 ( .B0(n6782), .B1(n218), .A0N(\ram[105][8] ), .A1N(n6505), 
        .Y(n2270) );
  OAI2BB2XL U2503 ( .B0(n6759), .B1(n218), .A0N(\ram[105][9] ), .A1N(n6505), 
        .Y(n2271) );
  OAI2BB2XL U2504 ( .B0(n6736), .B1(n218), .A0N(\ram[105][10] ), .A1N(n6505), 
        .Y(n2272) );
  OAI2BB2XL U2505 ( .B0(n6713), .B1(n218), .A0N(\ram[105][11] ), .A1N(n6505), 
        .Y(n2273) );
  OAI2BB2XL U2506 ( .B0(n6690), .B1(n218), .A0N(\ram[105][12] ), .A1N(n6505), 
        .Y(n2274) );
  OAI2BB2XL U2507 ( .B0(n6667), .B1(n218), .A0N(\ram[105][13] ), .A1N(n6505), 
        .Y(n2275) );
  OAI2BB2XL U2508 ( .B0(n6644), .B1(n218), .A0N(\ram[105][14] ), .A1N(n6505), 
        .Y(n2276) );
  OAI2BB2XL U2509 ( .B0(n6621), .B1(n218), .A0N(\ram[105][15] ), .A1N(n6505), 
        .Y(n2277) );
  OAI2BB2XL U2510 ( .B0(n6971), .B1(n462), .A0N(\ram[106][0] ), .A1N(n6504), 
        .Y(n2278) );
  OAI2BB2XL U2511 ( .B0(n6948), .B1(n462), .A0N(\ram[106][1] ), .A1N(n6504), 
        .Y(n2279) );
  OAI2BB2XL U2512 ( .B0(n6925), .B1(n462), .A0N(\ram[106][2] ), .A1N(n6504), 
        .Y(n2280) );
  OAI2BB2XL U2513 ( .B0(n6902), .B1(n462), .A0N(\ram[106][3] ), .A1N(n6504), 
        .Y(n2281) );
  OAI2BB2XL U2514 ( .B0(n6874), .B1(n462), .A0N(\ram[106][4] ), .A1N(n6504), 
        .Y(n2282) );
  OAI2BB2XL U2515 ( .B0(n6851), .B1(n462), .A0N(\ram[106][5] ), .A1N(n6504), 
        .Y(n2283) );
  OAI2BB2XL U2516 ( .B0(n6828), .B1(n462), .A0N(\ram[106][6] ), .A1N(n6504), 
        .Y(n2284) );
  OAI2BB2XL U2517 ( .B0(n6805), .B1(n462), .A0N(\ram[106][7] ), .A1N(n6504), 
        .Y(n2285) );
  OAI2BB2XL U2518 ( .B0(n6782), .B1(n462), .A0N(\ram[106][8] ), .A1N(n6504), 
        .Y(n2286) );
  OAI2BB2XL U2519 ( .B0(n6759), .B1(n462), .A0N(\ram[106][9] ), .A1N(n6504), 
        .Y(n2287) );
  OAI2BB2XL U2520 ( .B0(n6736), .B1(n462), .A0N(\ram[106][10] ), .A1N(n6504), 
        .Y(n2288) );
  OAI2BB2XL U2521 ( .B0(n6713), .B1(n462), .A0N(\ram[106][11] ), .A1N(n6504), 
        .Y(n2289) );
  OAI2BB2XL U2522 ( .B0(n6690), .B1(n462), .A0N(\ram[106][12] ), .A1N(n6504), 
        .Y(n2290) );
  OAI2BB2XL U2523 ( .B0(n6667), .B1(n462), .A0N(\ram[106][13] ), .A1N(n6504), 
        .Y(n2291) );
  OAI2BB2XL U2524 ( .B0(n6644), .B1(n462), .A0N(\ram[106][14] ), .A1N(n6504), 
        .Y(n2292) );
  OAI2BB2XL U2525 ( .B0(n6621), .B1(n462), .A0N(\ram[106][15] ), .A1N(n6504), 
        .Y(n2293) );
  OAI2BB2XL U2526 ( .B0(n6971), .B1(n220), .A0N(\ram[107][0] ), .A1N(n6503), 
        .Y(n2294) );
  OAI2BB2XL U2527 ( .B0(n6948), .B1(n220), .A0N(\ram[107][1] ), .A1N(n6503), 
        .Y(n2295) );
  OAI2BB2XL U2528 ( .B0(n6925), .B1(n220), .A0N(\ram[107][2] ), .A1N(n6503), 
        .Y(n2296) );
  OAI2BB2XL U2529 ( .B0(n6902), .B1(n220), .A0N(\ram[107][3] ), .A1N(n6503), 
        .Y(n2297) );
  OAI2BB2XL U2530 ( .B0(n6874), .B1(n220), .A0N(\ram[107][4] ), .A1N(n6503), 
        .Y(n2298) );
  OAI2BB2XL U2531 ( .B0(n6851), .B1(n220), .A0N(\ram[107][5] ), .A1N(n6503), 
        .Y(n2299) );
  OAI2BB2XL U2532 ( .B0(n6828), .B1(n220), .A0N(\ram[107][6] ), .A1N(n6503), 
        .Y(n2300) );
  OAI2BB2XL U2533 ( .B0(n6805), .B1(n220), .A0N(\ram[107][7] ), .A1N(n6503), 
        .Y(n2301) );
  OAI2BB2XL U2534 ( .B0(n6782), .B1(n220), .A0N(\ram[107][8] ), .A1N(n6503), 
        .Y(n2302) );
  OAI2BB2XL U2535 ( .B0(n6759), .B1(n220), .A0N(\ram[107][9] ), .A1N(n6503), 
        .Y(n2303) );
  OAI2BB2XL U2536 ( .B0(n6736), .B1(n220), .A0N(\ram[107][10] ), .A1N(n6503), 
        .Y(n2304) );
  OAI2BB2XL U2537 ( .B0(n6713), .B1(n220), .A0N(\ram[107][11] ), .A1N(n6503), 
        .Y(n2305) );
  OAI2BB2XL U2538 ( .B0(n6690), .B1(n220), .A0N(\ram[107][12] ), .A1N(n6503), 
        .Y(n2306) );
  OAI2BB2XL U2539 ( .B0(n6667), .B1(n220), .A0N(\ram[107][13] ), .A1N(n6503), 
        .Y(n2307) );
  OAI2BB2XL U2540 ( .B0(n6644), .B1(n220), .A0N(\ram[107][14] ), .A1N(n6503), 
        .Y(n2308) );
  OAI2BB2XL U2541 ( .B0(n6621), .B1(n220), .A0N(\ram[107][15] ), .A1N(n6503), 
        .Y(n2309) );
  OAI2BB2XL U2542 ( .B0(n6971), .B1(n222), .A0N(\ram[108][0] ), .A1N(n6502), 
        .Y(n2310) );
  OAI2BB2XL U2543 ( .B0(n6948), .B1(n222), .A0N(\ram[108][1] ), .A1N(n6502), 
        .Y(n2311) );
  OAI2BB2XL U2544 ( .B0(n6925), .B1(n222), .A0N(\ram[108][2] ), .A1N(n6502), 
        .Y(n2312) );
  OAI2BB2XL U2545 ( .B0(n6902), .B1(n222), .A0N(\ram[108][3] ), .A1N(n6502), 
        .Y(n2313) );
  OAI2BB2XL U2546 ( .B0(n6874), .B1(n222), .A0N(\ram[108][4] ), .A1N(n6502), 
        .Y(n2314) );
  OAI2BB2XL U2547 ( .B0(n6851), .B1(n222), .A0N(\ram[108][5] ), .A1N(n6502), 
        .Y(n2315) );
  OAI2BB2XL U2548 ( .B0(n6828), .B1(n222), .A0N(\ram[108][6] ), .A1N(n6502), 
        .Y(n2316) );
  OAI2BB2XL U2549 ( .B0(n6805), .B1(n222), .A0N(\ram[108][7] ), .A1N(n6502), 
        .Y(n2317) );
  OAI2BB2XL U2550 ( .B0(n6782), .B1(n222), .A0N(\ram[108][8] ), .A1N(n6502), 
        .Y(n2318) );
  OAI2BB2XL U2551 ( .B0(n6759), .B1(n222), .A0N(\ram[108][9] ), .A1N(n6502), 
        .Y(n2319) );
  OAI2BB2XL U2552 ( .B0(n6736), .B1(n222), .A0N(\ram[108][10] ), .A1N(n6502), 
        .Y(n2320) );
  OAI2BB2XL U2553 ( .B0(n6713), .B1(n222), .A0N(\ram[108][11] ), .A1N(n6502), 
        .Y(n2321) );
  OAI2BB2XL U2554 ( .B0(n6690), .B1(n222), .A0N(\ram[108][12] ), .A1N(n6502), 
        .Y(n2322) );
  OAI2BB2XL U2555 ( .B0(n6667), .B1(n222), .A0N(\ram[108][13] ), .A1N(n6502), 
        .Y(n2323) );
  OAI2BB2XL U2556 ( .B0(n6644), .B1(n222), .A0N(\ram[108][14] ), .A1N(n6502), 
        .Y(n2324) );
  OAI2BB2XL U2557 ( .B0(n6621), .B1(n222), .A0N(\ram[108][15] ), .A1N(n6502), 
        .Y(n2325) );
  OAI2BB2XL U2558 ( .B0(n6971), .B1(n224), .A0N(\ram[109][0] ), .A1N(n6501), 
        .Y(n2326) );
  OAI2BB2XL U2559 ( .B0(n6948), .B1(n224), .A0N(\ram[109][1] ), .A1N(n6501), 
        .Y(n2327) );
  OAI2BB2XL U2560 ( .B0(n6925), .B1(n224), .A0N(\ram[109][2] ), .A1N(n6501), 
        .Y(n2328) );
  OAI2BB2XL U2561 ( .B0(n6902), .B1(n224), .A0N(\ram[109][3] ), .A1N(n6501), 
        .Y(n2329) );
  OAI2BB2XL U2562 ( .B0(n6874), .B1(n224), .A0N(\ram[109][4] ), .A1N(n6501), 
        .Y(n2330) );
  OAI2BB2XL U2563 ( .B0(n6851), .B1(n224), .A0N(\ram[109][5] ), .A1N(n6501), 
        .Y(n2331) );
  OAI2BB2XL U2564 ( .B0(n6828), .B1(n224), .A0N(\ram[109][6] ), .A1N(n6501), 
        .Y(n2332) );
  OAI2BB2XL U2565 ( .B0(n6805), .B1(n224), .A0N(\ram[109][7] ), .A1N(n6501), 
        .Y(n2333) );
  OAI2BB2XL U2566 ( .B0(n6782), .B1(n224), .A0N(\ram[109][8] ), .A1N(n6501), 
        .Y(n2334) );
  OAI2BB2XL U2567 ( .B0(n6759), .B1(n224), .A0N(\ram[109][9] ), .A1N(n6501), 
        .Y(n2335) );
  OAI2BB2XL U2568 ( .B0(n6736), .B1(n224), .A0N(\ram[109][10] ), .A1N(n6501), 
        .Y(n2336) );
  OAI2BB2XL U2569 ( .B0(n6713), .B1(n224), .A0N(\ram[109][11] ), .A1N(n6501), 
        .Y(n2337) );
  OAI2BB2XL U2570 ( .B0(n6690), .B1(n224), .A0N(\ram[109][12] ), .A1N(n6501), 
        .Y(n2338) );
  OAI2BB2XL U2571 ( .B0(n6667), .B1(n224), .A0N(\ram[109][13] ), .A1N(n6501), 
        .Y(n2339) );
  OAI2BB2XL U2572 ( .B0(n6644), .B1(n224), .A0N(\ram[109][14] ), .A1N(n6501), 
        .Y(n2340) );
  OAI2BB2XL U2573 ( .B0(n6621), .B1(n224), .A0N(\ram[109][15] ), .A1N(n6501), 
        .Y(n2341) );
  OAI2BB2XL U2574 ( .B0(n6971), .B1(n226), .A0N(\ram[110][0] ), .A1N(n6500), 
        .Y(n2342) );
  OAI2BB2XL U2575 ( .B0(n6948), .B1(n226), .A0N(\ram[110][1] ), .A1N(n6500), 
        .Y(n2343) );
  OAI2BB2XL U2576 ( .B0(n6925), .B1(n226), .A0N(\ram[110][2] ), .A1N(n6500), 
        .Y(n2344) );
  OAI2BB2XL U2577 ( .B0(n6902), .B1(n226), .A0N(\ram[110][3] ), .A1N(n6500), 
        .Y(n2345) );
  OAI2BB2XL U2578 ( .B0(n6874), .B1(n226), .A0N(\ram[110][4] ), .A1N(n6500), 
        .Y(n2346) );
  OAI2BB2XL U2579 ( .B0(n6851), .B1(n226), .A0N(\ram[110][5] ), .A1N(n6500), 
        .Y(n2347) );
  OAI2BB2XL U2580 ( .B0(n6828), .B1(n226), .A0N(\ram[110][6] ), .A1N(n6500), 
        .Y(n2348) );
  OAI2BB2XL U2581 ( .B0(n6805), .B1(n226), .A0N(\ram[110][7] ), .A1N(n6500), 
        .Y(n2349) );
  OAI2BB2XL U2582 ( .B0(n6782), .B1(n226), .A0N(\ram[110][8] ), .A1N(n6500), 
        .Y(n2350) );
  OAI2BB2XL U2583 ( .B0(n6759), .B1(n226), .A0N(\ram[110][9] ), .A1N(n6500), 
        .Y(n2351) );
  OAI2BB2XL U2584 ( .B0(n6736), .B1(n226), .A0N(\ram[110][10] ), .A1N(n6500), 
        .Y(n2352) );
  OAI2BB2XL U2585 ( .B0(n6713), .B1(n226), .A0N(\ram[110][11] ), .A1N(n6500), 
        .Y(n2353) );
  OAI2BB2XL U2586 ( .B0(n6690), .B1(n226), .A0N(\ram[110][12] ), .A1N(n6500), 
        .Y(n2354) );
  OAI2BB2XL U2587 ( .B0(n6667), .B1(n226), .A0N(\ram[110][13] ), .A1N(n6500), 
        .Y(n2355) );
  OAI2BB2XL U2588 ( .B0(n6644), .B1(n226), .A0N(\ram[110][14] ), .A1N(n6500), 
        .Y(n2356) );
  OAI2BB2XL U2589 ( .B0(n6621), .B1(n226), .A0N(\ram[110][15] ), .A1N(n6500), 
        .Y(n2357) );
  OAI2BB2XL U2590 ( .B0(n6971), .B1(n228), .A0N(\ram[111][0] ), .A1N(n6499), 
        .Y(n2358) );
  OAI2BB2XL U2591 ( .B0(n6948), .B1(n228), .A0N(\ram[111][1] ), .A1N(n6499), 
        .Y(n2359) );
  OAI2BB2XL U2592 ( .B0(n6925), .B1(n228), .A0N(\ram[111][2] ), .A1N(n6499), 
        .Y(n2360) );
  OAI2BB2XL U2593 ( .B0(n6902), .B1(n228), .A0N(\ram[111][3] ), .A1N(n6499), 
        .Y(n2361) );
  OAI2BB2XL U2594 ( .B0(n6874), .B1(n228), .A0N(\ram[111][4] ), .A1N(n6499), 
        .Y(n2362) );
  OAI2BB2XL U2595 ( .B0(n6851), .B1(n228), .A0N(\ram[111][5] ), .A1N(n6499), 
        .Y(n2363) );
  OAI2BB2XL U2596 ( .B0(n6828), .B1(n228), .A0N(\ram[111][6] ), .A1N(n6499), 
        .Y(n2364) );
  OAI2BB2XL U2597 ( .B0(n6805), .B1(n228), .A0N(\ram[111][7] ), .A1N(n6499), 
        .Y(n2365) );
  OAI2BB2XL U2598 ( .B0(n6782), .B1(n228), .A0N(\ram[111][8] ), .A1N(n6499), 
        .Y(n2366) );
  OAI2BB2XL U2599 ( .B0(n6759), .B1(n228), .A0N(\ram[111][9] ), .A1N(n6499), 
        .Y(n2367) );
  OAI2BB2XL U2600 ( .B0(n6736), .B1(n228), .A0N(\ram[111][10] ), .A1N(n6499), 
        .Y(n2368) );
  OAI2BB2XL U2601 ( .B0(n6713), .B1(n228), .A0N(\ram[111][11] ), .A1N(n6499), 
        .Y(n2369) );
  OAI2BB2XL U2602 ( .B0(n6690), .B1(n228), .A0N(\ram[111][12] ), .A1N(n6499), 
        .Y(n2370) );
  OAI2BB2XL U2603 ( .B0(n6667), .B1(n228), .A0N(\ram[111][13] ), .A1N(n6499), 
        .Y(n2371) );
  OAI2BB2XL U2604 ( .B0(n6644), .B1(n228), .A0N(\ram[111][14] ), .A1N(n6499), 
        .Y(n2372) );
  OAI2BB2XL U2605 ( .B0(n6621), .B1(n228), .A0N(\ram[111][15] ), .A1N(n6499), 
        .Y(n2373) );
  OAI2BB2XL U2606 ( .B0(n6970), .B1(n230), .A0N(\ram[112][0] ), .A1N(n6498), 
        .Y(n2374) );
  OAI2BB2XL U2607 ( .B0(n6947), .B1(n230), .A0N(\ram[112][1] ), .A1N(n6498), 
        .Y(n2375) );
  OAI2BB2XL U2608 ( .B0(n6924), .B1(n230), .A0N(\ram[112][2] ), .A1N(n6498), 
        .Y(n2376) );
  OAI2BB2XL U2609 ( .B0(n6901), .B1(n230), .A0N(\ram[112][3] ), .A1N(n6498), 
        .Y(n2377) );
  OAI2BB2XL U2610 ( .B0(n6873), .B1(n230), .A0N(\ram[112][4] ), .A1N(n6498), 
        .Y(n2378) );
  OAI2BB2XL U2611 ( .B0(n6850), .B1(n230), .A0N(\ram[112][5] ), .A1N(n6498), 
        .Y(n2379) );
  OAI2BB2XL U2612 ( .B0(n6827), .B1(n230), .A0N(\ram[112][6] ), .A1N(n6498), 
        .Y(n2380) );
  OAI2BB2XL U2613 ( .B0(n6804), .B1(n230), .A0N(\ram[112][7] ), .A1N(n6498), 
        .Y(n2381) );
  OAI2BB2XL U2614 ( .B0(n6781), .B1(n230), .A0N(\ram[112][8] ), .A1N(n6498), 
        .Y(n2382) );
  OAI2BB2XL U2615 ( .B0(n6758), .B1(n230), .A0N(\ram[112][9] ), .A1N(n6498), 
        .Y(n2383) );
  OAI2BB2XL U2616 ( .B0(n6735), .B1(n230), .A0N(\ram[112][10] ), .A1N(n6498), 
        .Y(n2384) );
  OAI2BB2XL U2617 ( .B0(n6712), .B1(n230), .A0N(\ram[112][11] ), .A1N(n6498), 
        .Y(n2385) );
  OAI2BB2XL U2618 ( .B0(n6689), .B1(n230), .A0N(\ram[112][12] ), .A1N(n6498), 
        .Y(n2386) );
  OAI2BB2XL U2619 ( .B0(n6666), .B1(n230), .A0N(\ram[112][13] ), .A1N(n6498), 
        .Y(n2387) );
  OAI2BB2XL U2620 ( .B0(n6643), .B1(n230), .A0N(\ram[112][14] ), .A1N(n6498), 
        .Y(n2388) );
  OAI2BB2XL U2621 ( .B0(n6620), .B1(n230), .A0N(\ram[112][15] ), .A1N(n6498), 
        .Y(n2389) );
  OAI2BB2XL U2622 ( .B0(n6970), .B1(n232), .A0N(\ram[113][0] ), .A1N(n6497), 
        .Y(n2390) );
  OAI2BB2XL U2623 ( .B0(n6947), .B1(n232), .A0N(\ram[113][1] ), .A1N(n6497), 
        .Y(n2391) );
  OAI2BB2XL U2624 ( .B0(n6924), .B1(n232), .A0N(\ram[113][2] ), .A1N(n6497), 
        .Y(n2392) );
  OAI2BB2XL U2625 ( .B0(n6901), .B1(n232), .A0N(\ram[113][3] ), .A1N(n6497), 
        .Y(n2393) );
  OAI2BB2XL U2626 ( .B0(n6873), .B1(n232), .A0N(\ram[113][4] ), .A1N(n6497), 
        .Y(n2394) );
  OAI2BB2XL U2627 ( .B0(n6850), .B1(n232), .A0N(\ram[113][5] ), .A1N(n6497), 
        .Y(n2395) );
  OAI2BB2XL U2628 ( .B0(n6827), .B1(n232), .A0N(\ram[113][6] ), .A1N(n6497), 
        .Y(n2396) );
  OAI2BB2XL U2629 ( .B0(n6804), .B1(n232), .A0N(\ram[113][7] ), .A1N(n6497), 
        .Y(n2397) );
  OAI2BB2XL U2630 ( .B0(n6781), .B1(n232), .A0N(\ram[113][8] ), .A1N(n6497), 
        .Y(n2398) );
  OAI2BB2XL U2631 ( .B0(n6758), .B1(n232), .A0N(\ram[113][9] ), .A1N(n6497), 
        .Y(n2399) );
  OAI2BB2XL U2632 ( .B0(n6735), .B1(n232), .A0N(\ram[113][10] ), .A1N(n6497), 
        .Y(n2400) );
  OAI2BB2XL U2633 ( .B0(n6712), .B1(n232), .A0N(\ram[113][11] ), .A1N(n6497), 
        .Y(n2401) );
  OAI2BB2XL U2634 ( .B0(n6689), .B1(n232), .A0N(\ram[113][12] ), .A1N(n6497), 
        .Y(n2402) );
  OAI2BB2XL U2635 ( .B0(n6666), .B1(n232), .A0N(\ram[113][13] ), .A1N(n6497), 
        .Y(n2403) );
  OAI2BB2XL U2636 ( .B0(n6643), .B1(n232), .A0N(\ram[113][14] ), .A1N(n6497), 
        .Y(n2404) );
  OAI2BB2XL U2637 ( .B0(n6620), .B1(n232), .A0N(\ram[113][15] ), .A1N(n6497), 
        .Y(n2405) );
  OAI2BB2XL U2638 ( .B0(n6970), .B1(n234), .A0N(\ram[114][0] ), .A1N(n6496), 
        .Y(n2406) );
  OAI2BB2XL U2639 ( .B0(n6947), .B1(n234), .A0N(\ram[114][1] ), .A1N(n6496), 
        .Y(n2407) );
  OAI2BB2XL U2640 ( .B0(n6924), .B1(n234), .A0N(\ram[114][2] ), .A1N(n6496), 
        .Y(n2408) );
  OAI2BB2XL U2641 ( .B0(n6901), .B1(n234), .A0N(\ram[114][3] ), .A1N(n6496), 
        .Y(n2409) );
  OAI2BB2XL U2642 ( .B0(n6873), .B1(n234), .A0N(\ram[114][4] ), .A1N(n6496), 
        .Y(n2410) );
  OAI2BB2XL U2643 ( .B0(n6850), .B1(n234), .A0N(\ram[114][5] ), .A1N(n6496), 
        .Y(n2411) );
  OAI2BB2XL U2644 ( .B0(n6827), .B1(n234), .A0N(\ram[114][6] ), .A1N(n6496), 
        .Y(n2412) );
  OAI2BB2XL U2645 ( .B0(n6804), .B1(n234), .A0N(\ram[114][7] ), .A1N(n6496), 
        .Y(n2413) );
  OAI2BB2XL U2646 ( .B0(n6781), .B1(n234), .A0N(\ram[114][8] ), .A1N(n6496), 
        .Y(n2414) );
  OAI2BB2XL U2647 ( .B0(n6758), .B1(n234), .A0N(\ram[114][9] ), .A1N(n6496), 
        .Y(n2415) );
  OAI2BB2XL U2648 ( .B0(n6735), .B1(n234), .A0N(\ram[114][10] ), .A1N(n6496), 
        .Y(n2416) );
  OAI2BB2XL U2649 ( .B0(n6712), .B1(n234), .A0N(\ram[114][11] ), .A1N(n6496), 
        .Y(n2417) );
  OAI2BB2XL U2650 ( .B0(n6689), .B1(n234), .A0N(\ram[114][12] ), .A1N(n6496), 
        .Y(n2418) );
  OAI2BB2XL U2651 ( .B0(n6666), .B1(n234), .A0N(\ram[114][13] ), .A1N(n6496), 
        .Y(n2419) );
  OAI2BB2XL U2652 ( .B0(n6643), .B1(n234), .A0N(\ram[114][14] ), .A1N(n6496), 
        .Y(n2420) );
  OAI2BB2XL U2653 ( .B0(n6620), .B1(n234), .A0N(\ram[114][15] ), .A1N(n6496), 
        .Y(n2421) );
  OAI2BB2XL U2654 ( .B0(n6970), .B1(n236), .A0N(\ram[115][0] ), .A1N(n6495), 
        .Y(n2422) );
  OAI2BB2XL U2655 ( .B0(n6947), .B1(n236), .A0N(\ram[115][1] ), .A1N(n6495), 
        .Y(n2423) );
  OAI2BB2XL U2656 ( .B0(n6924), .B1(n236), .A0N(\ram[115][2] ), .A1N(n6495), 
        .Y(n2424) );
  OAI2BB2XL U2657 ( .B0(n6901), .B1(n236), .A0N(\ram[115][3] ), .A1N(n6495), 
        .Y(n2425) );
  OAI2BB2XL U2658 ( .B0(n6873), .B1(n236), .A0N(\ram[115][4] ), .A1N(n6495), 
        .Y(n2426) );
  OAI2BB2XL U2659 ( .B0(n6850), .B1(n236), .A0N(\ram[115][5] ), .A1N(n6495), 
        .Y(n2427) );
  OAI2BB2XL U2660 ( .B0(n6827), .B1(n236), .A0N(\ram[115][6] ), .A1N(n6495), 
        .Y(n2428) );
  OAI2BB2XL U2661 ( .B0(n6804), .B1(n236), .A0N(\ram[115][7] ), .A1N(n6495), 
        .Y(n2429) );
  OAI2BB2XL U2662 ( .B0(n6781), .B1(n236), .A0N(\ram[115][8] ), .A1N(n6495), 
        .Y(n2430) );
  OAI2BB2XL U2663 ( .B0(n6758), .B1(n236), .A0N(\ram[115][9] ), .A1N(n6495), 
        .Y(n2431) );
  OAI2BB2XL U2664 ( .B0(n6735), .B1(n236), .A0N(\ram[115][10] ), .A1N(n6495), 
        .Y(n2432) );
  OAI2BB2XL U2665 ( .B0(n6712), .B1(n236), .A0N(\ram[115][11] ), .A1N(n6495), 
        .Y(n2433) );
  OAI2BB2XL U2666 ( .B0(n6689), .B1(n236), .A0N(\ram[115][12] ), .A1N(n6495), 
        .Y(n2434) );
  OAI2BB2XL U2667 ( .B0(n6666), .B1(n236), .A0N(\ram[115][13] ), .A1N(n6495), 
        .Y(n2435) );
  OAI2BB2XL U2668 ( .B0(n6643), .B1(n236), .A0N(\ram[115][14] ), .A1N(n6495), 
        .Y(n2436) );
  OAI2BB2XL U2669 ( .B0(n6620), .B1(n236), .A0N(\ram[115][15] ), .A1N(n6495), 
        .Y(n2437) );
  OAI2BB2XL U2670 ( .B0(n6970), .B1(n238), .A0N(\ram[116][0] ), .A1N(n6494), 
        .Y(n2438) );
  OAI2BB2XL U2671 ( .B0(n6947), .B1(n238), .A0N(\ram[116][1] ), .A1N(n6494), 
        .Y(n2439) );
  OAI2BB2XL U2672 ( .B0(n6924), .B1(n238), .A0N(\ram[116][2] ), .A1N(n6494), 
        .Y(n2440) );
  OAI2BB2XL U2673 ( .B0(n6901), .B1(n238), .A0N(\ram[116][3] ), .A1N(n6494), 
        .Y(n2441) );
  OAI2BB2XL U2674 ( .B0(n6873), .B1(n238), .A0N(\ram[116][4] ), .A1N(n6494), 
        .Y(n2442) );
  OAI2BB2XL U2675 ( .B0(n6850), .B1(n238), .A0N(\ram[116][5] ), .A1N(n6494), 
        .Y(n2443) );
  OAI2BB2XL U2676 ( .B0(n6827), .B1(n238), .A0N(\ram[116][6] ), .A1N(n6494), 
        .Y(n2444) );
  OAI2BB2XL U2677 ( .B0(n6804), .B1(n238), .A0N(\ram[116][7] ), .A1N(n6494), 
        .Y(n2445) );
  OAI2BB2XL U2678 ( .B0(n6781), .B1(n238), .A0N(\ram[116][8] ), .A1N(n6494), 
        .Y(n2446) );
  OAI2BB2XL U2679 ( .B0(n6758), .B1(n238), .A0N(\ram[116][9] ), .A1N(n6494), 
        .Y(n2447) );
  OAI2BB2XL U2680 ( .B0(n6735), .B1(n238), .A0N(\ram[116][10] ), .A1N(n6494), 
        .Y(n2448) );
  OAI2BB2XL U2681 ( .B0(n6712), .B1(n238), .A0N(\ram[116][11] ), .A1N(n6494), 
        .Y(n2449) );
  OAI2BB2XL U2682 ( .B0(n6689), .B1(n238), .A0N(\ram[116][12] ), .A1N(n6494), 
        .Y(n2450) );
  OAI2BB2XL U2683 ( .B0(n6666), .B1(n238), .A0N(\ram[116][13] ), .A1N(n6494), 
        .Y(n2451) );
  OAI2BB2XL U2684 ( .B0(n6643), .B1(n238), .A0N(\ram[116][14] ), .A1N(n6494), 
        .Y(n2452) );
  OAI2BB2XL U2685 ( .B0(n6620), .B1(n238), .A0N(\ram[116][15] ), .A1N(n6494), 
        .Y(n2453) );
  OAI2BB2XL U2686 ( .B0(n6970), .B1(n240), .A0N(\ram[117][0] ), .A1N(n6493), 
        .Y(n2454) );
  OAI2BB2XL U2687 ( .B0(n6947), .B1(n240), .A0N(\ram[117][1] ), .A1N(n6493), 
        .Y(n2455) );
  OAI2BB2XL U2688 ( .B0(n6924), .B1(n240), .A0N(\ram[117][2] ), .A1N(n6493), 
        .Y(n2456) );
  OAI2BB2XL U2689 ( .B0(n6901), .B1(n240), .A0N(\ram[117][3] ), .A1N(n6493), 
        .Y(n2457) );
  OAI2BB2XL U2690 ( .B0(n6873), .B1(n240), .A0N(\ram[117][4] ), .A1N(n6493), 
        .Y(n2458) );
  OAI2BB2XL U2691 ( .B0(n6850), .B1(n240), .A0N(\ram[117][5] ), .A1N(n6493), 
        .Y(n2459) );
  OAI2BB2XL U2692 ( .B0(n6827), .B1(n240), .A0N(\ram[117][6] ), .A1N(n6493), 
        .Y(n2460) );
  OAI2BB2XL U2693 ( .B0(n6804), .B1(n240), .A0N(\ram[117][7] ), .A1N(n6493), 
        .Y(n2461) );
  OAI2BB2XL U2694 ( .B0(n6781), .B1(n240), .A0N(\ram[117][8] ), .A1N(n6493), 
        .Y(n2462) );
  OAI2BB2XL U2695 ( .B0(n6758), .B1(n240), .A0N(\ram[117][9] ), .A1N(n6493), 
        .Y(n2463) );
  OAI2BB2XL U2696 ( .B0(n6735), .B1(n240), .A0N(\ram[117][10] ), .A1N(n6493), 
        .Y(n2464) );
  OAI2BB2XL U2697 ( .B0(n6712), .B1(n240), .A0N(\ram[117][11] ), .A1N(n6493), 
        .Y(n2465) );
  OAI2BB2XL U2698 ( .B0(n6689), .B1(n240), .A0N(\ram[117][12] ), .A1N(n6493), 
        .Y(n2466) );
  OAI2BB2XL U2699 ( .B0(n6666), .B1(n240), .A0N(\ram[117][13] ), .A1N(n6493), 
        .Y(n2467) );
  OAI2BB2XL U2700 ( .B0(n6643), .B1(n240), .A0N(\ram[117][14] ), .A1N(n6493), 
        .Y(n2468) );
  OAI2BB2XL U2701 ( .B0(n6620), .B1(n240), .A0N(\ram[117][15] ), .A1N(n6493), 
        .Y(n2469) );
  OAI2BB2XL U2702 ( .B0(n6970), .B1(n242), .A0N(\ram[118][0] ), .A1N(n6492), 
        .Y(n2470) );
  OAI2BB2XL U2703 ( .B0(n6947), .B1(n242), .A0N(\ram[118][1] ), .A1N(n6492), 
        .Y(n2471) );
  OAI2BB2XL U2704 ( .B0(n6924), .B1(n242), .A0N(\ram[118][2] ), .A1N(n6492), 
        .Y(n2472) );
  OAI2BB2XL U2705 ( .B0(n6901), .B1(n242), .A0N(\ram[118][3] ), .A1N(n6492), 
        .Y(n2473) );
  OAI2BB2XL U2706 ( .B0(n6873), .B1(n242), .A0N(\ram[118][4] ), .A1N(n6492), 
        .Y(n2474) );
  OAI2BB2XL U2707 ( .B0(n6850), .B1(n242), .A0N(\ram[118][5] ), .A1N(n6492), 
        .Y(n2475) );
  OAI2BB2XL U2708 ( .B0(n6827), .B1(n242), .A0N(\ram[118][6] ), .A1N(n6492), 
        .Y(n2476) );
  OAI2BB2XL U2709 ( .B0(n6804), .B1(n242), .A0N(\ram[118][7] ), .A1N(n6492), 
        .Y(n2477) );
  OAI2BB2XL U2710 ( .B0(n6781), .B1(n242), .A0N(\ram[118][8] ), .A1N(n6492), 
        .Y(n2478) );
  OAI2BB2XL U2711 ( .B0(n6758), .B1(n242), .A0N(\ram[118][9] ), .A1N(n6492), 
        .Y(n2479) );
  OAI2BB2XL U2712 ( .B0(n6735), .B1(n242), .A0N(\ram[118][10] ), .A1N(n6492), 
        .Y(n2480) );
  OAI2BB2XL U2713 ( .B0(n6712), .B1(n242), .A0N(\ram[118][11] ), .A1N(n6492), 
        .Y(n2481) );
  OAI2BB2XL U2714 ( .B0(n6689), .B1(n242), .A0N(\ram[118][12] ), .A1N(n6492), 
        .Y(n2482) );
  OAI2BB2XL U2715 ( .B0(n6666), .B1(n242), .A0N(\ram[118][13] ), .A1N(n6492), 
        .Y(n2483) );
  OAI2BB2XL U2716 ( .B0(n6643), .B1(n242), .A0N(\ram[118][14] ), .A1N(n6492), 
        .Y(n2484) );
  OAI2BB2XL U2717 ( .B0(n6620), .B1(n242), .A0N(\ram[118][15] ), .A1N(n6492), 
        .Y(n2485) );
  OAI2BB2XL U2718 ( .B0(n6970), .B1(n244), .A0N(\ram[119][0] ), .A1N(n6491), 
        .Y(n2486) );
  OAI2BB2XL U2719 ( .B0(n6947), .B1(n244), .A0N(\ram[119][1] ), .A1N(n6491), 
        .Y(n2487) );
  OAI2BB2XL U2720 ( .B0(n6924), .B1(n244), .A0N(\ram[119][2] ), .A1N(n6491), 
        .Y(n2488) );
  OAI2BB2XL U2721 ( .B0(n6901), .B1(n244), .A0N(\ram[119][3] ), .A1N(n6491), 
        .Y(n2489) );
  OAI2BB2XL U2722 ( .B0(n6873), .B1(n244), .A0N(\ram[119][4] ), .A1N(n6491), 
        .Y(n2490) );
  OAI2BB2XL U2723 ( .B0(n6850), .B1(n244), .A0N(\ram[119][5] ), .A1N(n6491), 
        .Y(n2491) );
  OAI2BB2XL U2724 ( .B0(n6827), .B1(n244), .A0N(\ram[119][6] ), .A1N(n6491), 
        .Y(n2492) );
  OAI2BB2XL U2725 ( .B0(n6804), .B1(n244), .A0N(\ram[119][7] ), .A1N(n6491), 
        .Y(n2493) );
  OAI2BB2XL U2726 ( .B0(n6781), .B1(n244), .A0N(\ram[119][8] ), .A1N(n6491), 
        .Y(n2494) );
  OAI2BB2XL U2727 ( .B0(n6758), .B1(n244), .A0N(\ram[119][9] ), .A1N(n6491), 
        .Y(n2495) );
  OAI2BB2XL U2728 ( .B0(n6735), .B1(n244), .A0N(\ram[119][10] ), .A1N(n6491), 
        .Y(n2496) );
  OAI2BB2XL U2729 ( .B0(n6712), .B1(n244), .A0N(\ram[119][11] ), .A1N(n6491), 
        .Y(n2497) );
  OAI2BB2XL U2730 ( .B0(n6689), .B1(n244), .A0N(\ram[119][12] ), .A1N(n6491), 
        .Y(n2498) );
  OAI2BB2XL U2731 ( .B0(n6666), .B1(n244), .A0N(\ram[119][13] ), .A1N(n6491), 
        .Y(n2499) );
  OAI2BB2XL U2732 ( .B0(n6643), .B1(n244), .A0N(\ram[119][14] ), .A1N(n6491), 
        .Y(n2500) );
  OAI2BB2XL U2733 ( .B0(n6620), .B1(n244), .A0N(\ram[119][15] ), .A1N(n6491), 
        .Y(n2501) );
  OAI2BB2XL U2734 ( .B0(n6970), .B1(n245), .A0N(\ram[120][0] ), .A1N(n6490), 
        .Y(n2502) );
  OAI2BB2XL U2735 ( .B0(n6947), .B1(n245), .A0N(\ram[120][1] ), .A1N(n6490), 
        .Y(n2503) );
  OAI2BB2XL U2736 ( .B0(n6924), .B1(n245), .A0N(\ram[120][2] ), .A1N(n6490), 
        .Y(n2504) );
  OAI2BB2XL U2737 ( .B0(n6901), .B1(n245), .A0N(\ram[120][3] ), .A1N(n6490), 
        .Y(n2505) );
  OAI2BB2XL U2738 ( .B0(n6873), .B1(n245), .A0N(\ram[120][4] ), .A1N(n6490), 
        .Y(n2506) );
  OAI2BB2XL U2739 ( .B0(n6850), .B1(n245), .A0N(\ram[120][5] ), .A1N(n6490), 
        .Y(n2507) );
  OAI2BB2XL U2740 ( .B0(n6827), .B1(n245), .A0N(\ram[120][6] ), .A1N(n6490), 
        .Y(n2508) );
  OAI2BB2XL U2741 ( .B0(n6804), .B1(n245), .A0N(\ram[120][7] ), .A1N(n6490), 
        .Y(n2509) );
  OAI2BB2XL U2742 ( .B0(n6781), .B1(n245), .A0N(\ram[120][8] ), .A1N(n6490), 
        .Y(n2510) );
  OAI2BB2XL U2743 ( .B0(n6758), .B1(n245), .A0N(\ram[120][9] ), .A1N(n6490), 
        .Y(n2511) );
  OAI2BB2XL U2744 ( .B0(n6735), .B1(n245), .A0N(\ram[120][10] ), .A1N(n6490), 
        .Y(n2512) );
  OAI2BB2XL U2745 ( .B0(n6712), .B1(n245), .A0N(\ram[120][11] ), .A1N(n6490), 
        .Y(n2513) );
  OAI2BB2XL U2746 ( .B0(n6689), .B1(n245), .A0N(\ram[120][12] ), .A1N(n6490), 
        .Y(n2514) );
  OAI2BB2XL U2747 ( .B0(n6666), .B1(n245), .A0N(\ram[120][13] ), .A1N(n6490), 
        .Y(n2515) );
  OAI2BB2XL U2748 ( .B0(n6643), .B1(n245), .A0N(\ram[120][14] ), .A1N(n6490), 
        .Y(n2516) );
  OAI2BB2XL U2749 ( .B0(n6620), .B1(n245), .A0N(\ram[120][15] ), .A1N(n6490), 
        .Y(n2517) );
  OAI2BB2XL U2750 ( .B0(n6970), .B1(n247), .A0N(\ram[121][0] ), .A1N(n6489), 
        .Y(n2518) );
  OAI2BB2XL U2751 ( .B0(n6947), .B1(n247), .A0N(\ram[121][1] ), .A1N(n6489), 
        .Y(n2519) );
  OAI2BB2XL U2752 ( .B0(n6924), .B1(n247), .A0N(\ram[121][2] ), .A1N(n6489), 
        .Y(n2520) );
  OAI2BB2XL U2753 ( .B0(n6901), .B1(n247), .A0N(\ram[121][3] ), .A1N(n6489), 
        .Y(n2521) );
  OAI2BB2XL U2754 ( .B0(n6873), .B1(n247), .A0N(\ram[121][4] ), .A1N(n6489), 
        .Y(n2522) );
  OAI2BB2XL U2755 ( .B0(n6850), .B1(n247), .A0N(\ram[121][5] ), .A1N(n6489), 
        .Y(n2523) );
  OAI2BB2XL U2756 ( .B0(n6827), .B1(n247), .A0N(\ram[121][6] ), .A1N(n6489), 
        .Y(n2524) );
  OAI2BB2XL U2757 ( .B0(n6804), .B1(n247), .A0N(\ram[121][7] ), .A1N(n6489), 
        .Y(n2525) );
  OAI2BB2XL U2758 ( .B0(n6781), .B1(n247), .A0N(\ram[121][8] ), .A1N(n6489), 
        .Y(n2526) );
  OAI2BB2XL U2759 ( .B0(n6758), .B1(n247), .A0N(\ram[121][9] ), .A1N(n6489), 
        .Y(n2527) );
  OAI2BB2XL U2760 ( .B0(n6735), .B1(n247), .A0N(\ram[121][10] ), .A1N(n6489), 
        .Y(n2528) );
  OAI2BB2XL U2761 ( .B0(n6712), .B1(n247), .A0N(\ram[121][11] ), .A1N(n6489), 
        .Y(n2529) );
  OAI2BB2XL U2762 ( .B0(n6689), .B1(n247), .A0N(\ram[121][12] ), .A1N(n6489), 
        .Y(n2530) );
  OAI2BB2XL U2763 ( .B0(n6666), .B1(n247), .A0N(\ram[121][13] ), .A1N(n6489), 
        .Y(n2531) );
  OAI2BB2XL U2764 ( .B0(n6643), .B1(n247), .A0N(\ram[121][14] ), .A1N(n6489), 
        .Y(n2532) );
  OAI2BB2XL U2765 ( .B0(n6620), .B1(n247), .A0N(\ram[121][15] ), .A1N(n6489), 
        .Y(n2533) );
  OAI2BB2XL U2766 ( .B0(n6970), .B1(n249), .A0N(\ram[122][0] ), .A1N(n6488), 
        .Y(n2534) );
  OAI2BB2XL U2767 ( .B0(n6947), .B1(n249), .A0N(\ram[122][1] ), .A1N(n6488), 
        .Y(n2535) );
  OAI2BB2XL U2768 ( .B0(n6924), .B1(n249), .A0N(\ram[122][2] ), .A1N(n6488), 
        .Y(n2536) );
  OAI2BB2XL U2769 ( .B0(n6901), .B1(n249), .A0N(\ram[122][3] ), .A1N(n6488), 
        .Y(n2537) );
  OAI2BB2XL U2770 ( .B0(n6873), .B1(n249), .A0N(\ram[122][4] ), .A1N(n6488), 
        .Y(n2538) );
  OAI2BB2XL U2771 ( .B0(n6850), .B1(n249), .A0N(\ram[122][5] ), .A1N(n6488), 
        .Y(n2539) );
  OAI2BB2XL U2772 ( .B0(n6827), .B1(n249), .A0N(\ram[122][6] ), .A1N(n6488), 
        .Y(n2540) );
  OAI2BB2XL U2773 ( .B0(n6804), .B1(n249), .A0N(\ram[122][7] ), .A1N(n6488), 
        .Y(n2541) );
  OAI2BB2XL U2774 ( .B0(n6781), .B1(n249), .A0N(\ram[122][8] ), .A1N(n6488), 
        .Y(n2542) );
  OAI2BB2XL U2775 ( .B0(n6758), .B1(n249), .A0N(\ram[122][9] ), .A1N(n6488), 
        .Y(n2543) );
  OAI2BB2XL U2776 ( .B0(n6735), .B1(n249), .A0N(\ram[122][10] ), .A1N(n6488), 
        .Y(n2544) );
  OAI2BB2XL U2777 ( .B0(n6712), .B1(n249), .A0N(\ram[122][11] ), .A1N(n6488), 
        .Y(n2545) );
  OAI2BB2XL U2778 ( .B0(n6689), .B1(n249), .A0N(\ram[122][12] ), .A1N(n6488), 
        .Y(n2546) );
  OAI2BB2XL U2779 ( .B0(n6666), .B1(n249), .A0N(\ram[122][13] ), .A1N(n6488), 
        .Y(n2547) );
  OAI2BB2XL U2780 ( .B0(n6643), .B1(n249), .A0N(\ram[122][14] ), .A1N(n6488), 
        .Y(n2548) );
  OAI2BB2XL U2781 ( .B0(n6620), .B1(n249), .A0N(\ram[122][15] ), .A1N(n6488), 
        .Y(n2549) );
  OAI2BB2XL U2782 ( .B0(n6970), .B1(n251), .A0N(\ram[123][0] ), .A1N(n6487), 
        .Y(n2550) );
  OAI2BB2XL U2783 ( .B0(n6947), .B1(n251), .A0N(\ram[123][1] ), .A1N(n6487), 
        .Y(n2551) );
  OAI2BB2XL U2784 ( .B0(n6924), .B1(n251), .A0N(\ram[123][2] ), .A1N(n6487), 
        .Y(n2552) );
  OAI2BB2XL U2785 ( .B0(n6901), .B1(n251), .A0N(\ram[123][3] ), .A1N(n6487), 
        .Y(n2553) );
  OAI2BB2XL U2786 ( .B0(n6873), .B1(n251), .A0N(\ram[123][4] ), .A1N(n6487), 
        .Y(n2554) );
  OAI2BB2XL U2787 ( .B0(n6850), .B1(n251), .A0N(\ram[123][5] ), .A1N(n6487), 
        .Y(n2555) );
  OAI2BB2XL U2788 ( .B0(n6827), .B1(n251), .A0N(\ram[123][6] ), .A1N(n6487), 
        .Y(n2556) );
  OAI2BB2XL U2789 ( .B0(n6804), .B1(n251), .A0N(\ram[123][7] ), .A1N(n6487), 
        .Y(n2557) );
  OAI2BB2XL U2790 ( .B0(n6781), .B1(n251), .A0N(\ram[123][8] ), .A1N(n6487), 
        .Y(n2558) );
  OAI2BB2XL U2791 ( .B0(n6758), .B1(n251), .A0N(\ram[123][9] ), .A1N(n6487), 
        .Y(n2559) );
  OAI2BB2XL U2792 ( .B0(n6735), .B1(n251), .A0N(\ram[123][10] ), .A1N(n6487), 
        .Y(n2560) );
  OAI2BB2XL U2793 ( .B0(n6712), .B1(n251), .A0N(\ram[123][11] ), .A1N(n6487), 
        .Y(n2561) );
  OAI2BB2XL U2794 ( .B0(n6689), .B1(n251), .A0N(\ram[123][12] ), .A1N(n6487), 
        .Y(n2562) );
  OAI2BB2XL U2795 ( .B0(n6666), .B1(n251), .A0N(\ram[123][13] ), .A1N(n6487), 
        .Y(n2563) );
  OAI2BB2XL U2796 ( .B0(n6643), .B1(n251), .A0N(\ram[123][14] ), .A1N(n6487), 
        .Y(n2564) );
  OAI2BB2XL U2797 ( .B0(n6620), .B1(n251), .A0N(\ram[123][15] ), .A1N(n6487), 
        .Y(n2565) );
  OAI2BB2XL U2798 ( .B0(n6969), .B1(n253), .A0N(\ram[124][0] ), .A1N(n6486), 
        .Y(n2566) );
  OAI2BB2XL U2799 ( .B0(n6946), .B1(n253), .A0N(\ram[124][1] ), .A1N(n6486), 
        .Y(n2567) );
  OAI2BB2XL U2800 ( .B0(n6923), .B1(n253), .A0N(\ram[124][2] ), .A1N(n6486), 
        .Y(n2568) );
  OAI2BB2XL U2801 ( .B0(n6900), .B1(n253), .A0N(\ram[124][3] ), .A1N(n6486), 
        .Y(n2569) );
  OAI2BB2XL U2802 ( .B0(n6872), .B1(n253), .A0N(\ram[124][4] ), .A1N(n6486), 
        .Y(n2570) );
  OAI2BB2XL U2803 ( .B0(n6849), .B1(n253), .A0N(\ram[124][5] ), .A1N(n6486), 
        .Y(n2571) );
  OAI2BB2XL U2804 ( .B0(n6826), .B1(n253), .A0N(\ram[124][6] ), .A1N(n6486), 
        .Y(n2572) );
  OAI2BB2XL U2805 ( .B0(n6803), .B1(n253), .A0N(\ram[124][7] ), .A1N(n6486), 
        .Y(n2573) );
  OAI2BB2XL U2806 ( .B0(n6780), .B1(n253), .A0N(\ram[124][8] ), .A1N(n6486), 
        .Y(n2574) );
  OAI2BB2XL U2807 ( .B0(n6757), .B1(n253), .A0N(\ram[124][9] ), .A1N(n6486), 
        .Y(n2575) );
  OAI2BB2XL U2808 ( .B0(n6734), .B1(n253), .A0N(\ram[124][10] ), .A1N(n6486), 
        .Y(n2576) );
  OAI2BB2XL U2809 ( .B0(n6711), .B1(n253), .A0N(\ram[124][11] ), .A1N(n6486), 
        .Y(n2577) );
  OAI2BB2XL U2810 ( .B0(n6688), .B1(n253), .A0N(\ram[124][12] ), .A1N(n6486), 
        .Y(n2578) );
  OAI2BB2XL U2811 ( .B0(n6665), .B1(n253), .A0N(\ram[124][13] ), .A1N(n6486), 
        .Y(n2579) );
  OAI2BB2XL U2812 ( .B0(n6642), .B1(n253), .A0N(\ram[124][14] ), .A1N(n6486), 
        .Y(n2580) );
  OAI2BB2XL U2813 ( .B0(n6619), .B1(n253), .A0N(\ram[124][15] ), .A1N(n6486), 
        .Y(n2581) );
  OAI2BB2XL U2814 ( .B0(n6969), .B1(n255), .A0N(\ram[125][0] ), .A1N(n6485), 
        .Y(n2582) );
  OAI2BB2XL U2815 ( .B0(n6946), .B1(n255), .A0N(\ram[125][1] ), .A1N(n6485), 
        .Y(n2583) );
  OAI2BB2XL U2816 ( .B0(n6923), .B1(n255), .A0N(\ram[125][2] ), .A1N(n6485), 
        .Y(n2584) );
  OAI2BB2XL U2817 ( .B0(n6900), .B1(n255), .A0N(\ram[125][3] ), .A1N(n6485), 
        .Y(n2585) );
  OAI2BB2XL U2818 ( .B0(n6872), .B1(n255), .A0N(\ram[125][4] ), .A1N(n6485), 
        .Y(n2586) );
  OAI2BB2XL U2819 ( .B0(n6849), .B1(n255), .A0N(\ram[125][5] ), .A1N(n6485), 
        .Y(n2587) );
  OAI2BB2XL U2820 ( .B0(n6826), .B1(n255), .A0N(\ram[125][6] ), .A1N(n6485), 
        .Y(n2588) );
  OAI2BB2XL U2821 ( .B0(n6803), .B1(n255), .A0N(\ram[125][7] ), .A1N(n6485), 
        .Y(n2589) );
  OAI2BB2XL U2822 ( .B0(n6780), .B1(n255), .A0N(\ram[125][8] ), .A1N(n6485), 
        .Y(n2590) );
  OAI2BB2XL U2823 ( .B0(n6757), .B1(n255), .A0N(\ram[125][9] ), .A1N(n6485), 
        .Y(n2591) );
  OAI2BB2XL U2824 ( .B0(n6734), .B1(n255), .A0N(\ram[125][10] ), .A1N(n6485), 
        .Y(n2592) );
  OAI2BB2XL U2825 ( .B0(n6711), .B1(n255), .A0N(\ram[125][11] ), .A1N(n6485), 
        .Y(n2593) );
  OAI2BB2XL U2826 ( .B0(n6688), .B1(n255), .A0N(\ram[125][12] ), .A1N(n6485), 
        .Y(n2594) );
  OAI2BB2XL U2827 ( .B0(n6665), .B1(n255), .A0N(\ram[125][13] ), .A1N(n6485), 
        .Y(n2595) );
  OAI2BB2XL U2828 ( .B0(n6642), .B1(n255), .A0N(\ram[125][14] ), .A1N(n6485), 
        .Y(n2596) );
  OAI2BB2XL U2829 ( .B0(n6619), .B1(n255), .A0N(\ram[125][15] ), .A1N(n6485), 
        .Y(n2597) );
  OAI2BB2XL U2830 ( .B0(n6969), .B1(n257), .A0N(\ram[126][0] ), .A1N(n6484), 
        .Y(n2598) );
  OAI2BB2XL U2831 ( .B0(n6946), .B1(n257), .A0N(\ram[126][1] ), .A1N(n6484), 
        .Y(n2599) );
  OAI2BB2XL U2832 ( .B0(n6923), .B1(n257), .A0N(\ram[126][2] ), .A1N(n6484), 
        .Y(n2600) );
  OAI2BB2XL U2833 ( .B0(n6900), .B1(n257), .A0N(\ram[126][3] ), .A1N(n6484), 
        .Y(n2601) );
  OAI2BB2XL U2834 ( .B0(n6872), .B1(n257), .A0N(\ram[126][4] ), .A1N(n6484), 
        .Y(n2602) );
  OAI2BB2XL U2835 ( .B0(n6849), .B1(n257), .A0N(\ram[126][5] ), .A1N(n6484), 
        .Y(n2603) );
  OAI2BB2XL U2836 ( .B0(n6826), .B1(n257), .A0N(\ram[126][6] ), .A1N(n6484), 
        .Y(n2604) );
  OAI2BB2XL U2837 ( .B0(n6803), .B1(n257), .A0N(\ram[126][7] ), .A1N(n6484), 
        .Y(n2605) );
  OAI2BB2XL U2838 ( .B0(n6780), .B1(n257), .A0N(\ram[126][8] ), .A1N(n6484), 
        .Y(n2606) );
  OAI2BB2XL U2839 ( .B0(n6757), .B1(n257), .A0N(\ram[126][9] ), .A1N(n6484), 
        .Y(n2607) );
  OAI2BB2XL U2840 ( .B0(n6734), .B1(n257), .A0N(\ram[126][10] ), .A1N(n6484), 
        .Y(n2608) );
  OAI2BB2XL U2841 ( .B0(n6711), .B1(n257), .A0N(\ram[126][11] ), .A1N(n6484), 
        .Y(n2609) );
  OAI2BB2XL U2842 ( .B0(n6688), .B1(n257), .A0N(\ram[126][12] ), .A1N(n6484), 
        .Y(n2610) );
  OAI2BB2XL U2843 ( .B0(n6665), .B1(n257), .A0N(\ram[126][13] ), .A1N(n6484), 
        .Y(n2611) );
  OAI2BB2XL U2844 ( .B0(n6642), .B1(n257), .A0N(\ram[126][14] ), .A1N(n6484), 
        .Y(n2612) );
  OAI2BB2XL U2845 ( .B0(n6619), .B1(n257), .A0N(\ram[126][15] ), .A1N(n6484), 
        .Y(n2613) );
  OAI2BB2XL U2846 ( .B0(n6969), .B1(n259), .A0N(\ram[127][0] ), .A1N(n6483), 
        .Y(n2614) );
  OAI2BB2XL U2847 ( .B0(n6946), .B1(n259), .A0N(\ram[127][1] ), .A1N(n6483), 
        .Y(n2615) );
  OAI2BB2XL U2848 ( .B0(n6923), .B1(n259), .A0N(\ram[127][2] ), .A1N(n6483), 
        .Y(n2616) );
  OAI2BB2XL U2849 ( .B0(n6900), .B1(n259), .A0N(\ram[127][3] ), .A1N(n6483), 
        .Y(n2617) );
  OAI2BB2XL U2850 ( .B0(n6872), .B1(n259), .A0N(\ram[127][4] ), .A1N(n6483), 
        .Y(n2618) );
  OAI2BB2XL U2851 ( .B0(n6849), .B1(n259), .A0N(\ram[127][5] ), .A1N(n6483), 
        .Y(n2619) );
  OAI2BB2XL U2852 ( .B0(n6826), .B1(n259), .A0N(\ram[127][6] ), .A1N(n6483), 
        .Y(n2620) );
  OAI2BB2XL U2853 ( .B0(n6803), .B1(n259), .A0N(\ram[127][7] ), .A1N(n6483), 
        .Y(n2621) );
  OAI2BB2XL U2854 ( .B0(n6780), .B1(n259), .A0N(\ram[127][8] ), .A1N(n6483), 
        .Y(n2622) );
  OAI2BB2XL U2855 ( .B0(n6757), .B1(n259), .A0N(\ram[127][9] ), .A1N(n6483), 
        .Y(n2623) );
  OAI2BB2XL U2856 ( .B0(n6734), .B1(n259), .A0N(\ram[127][10] ), .A1N(n6483), 
        .Y(n2624) );
  OAI2BB2XL U2857 ( .B0(n6711), .B1(n259), .A0N(\ram[127][11] ), .A1N(n6483), 
        .Y(n2625) );
  OAI2BB2XL U2858 ( .B0(n6688), .B1(n259), .A0N(\ram[127][12] ), .A1N(n6483), 
        .Y(n2626) );
  OAI2BB2XL U2859 ( .B0(n6665), .B1(n259), .A0N(\ram[127][13] ), .A1N(n6483), 
        .Y(n2627) );
  OAI2BB2XL U2860 ( .B0(n6642), .B1(n259), .A0N(\ram[127][14] ), .A1N(n6483), 
        .Y(n2628) );
  OAI2BB2XL U2861 ( .B0(n6619), .B1(n259), .A0N(\ram[127][15] ), .A1N(n6483), 
        .Y(n2629) );
  OAI2BB2XL U2862 ( .B0(n6968), .B1(n286), .A0N(\ram[144][0] ), .A1N(n6466), 
        .Y(n2886) );
  OAI2BB2XL U2863 ( .B0(n6945), .B1(n286), .A0N(\ram[144][1] ), .A1N(n6466), 
        .Y(n2887) );
  OAI2BB2XL U2864 ( .B0(n6922), .B1(n286), .A0N(\ram[144][2] ), .A1N(n6466), 
        .Y(n2888) );
  OAI2BB2XL U2865 ( .B0(n6899), .B1(n286), .A0N(\ram[144][3] ), .A1N(n6466), 
        .Y(n2889) );
  OAI2BB2XL U2866 ( .B0(n6871), .B1(n286), .A0N(\ram[144][4] ), .A1N(n6466), 
        .Y(n2890) );
  OAI2BB2XL U2867 ( .B0(n6848), .B1(n286), .A0N(\ram[144][5] ), .A1N(n6466), 
        .Y(n2891) );
  OAI2BB2XL U2868 ( .B0(n6825), .B1(n286), .A0N(\ram[144][6] ), .A1N(n6466), 
        .Y(n2892) );
  OAI2BB2XL U2869 ( .B0(n6802), .B1(n286), .A0N(\ram[144][7] ), .A1N(n6466), 
        .Y(n2893) );
  OAI2BB2XL U2870 ( .B0(n6779), .B1(n286), .A0N(\ram[144][8] ), .A1N(n6466), 
        .Y(n2894) );
  OAI2BB2XL U2871 ( .B0(n6756), .B1(n286), .A0N(\ram[144][9] ), .A1N(n6466), 
        .Y(n2895) );
  OAI2BB2XL U2872 ( .B0(n6733), .B1(n286), .A0N(\ram[144][10] ), .A1N(n6466), 
        .Y(n2896) );
  OAI2BB2XL U2873 ( .B0(n6710), .B1(n286), .A0N(\ram[144][11] ), .A1N(n6466), 
        .Y(n2897) );
  OAI2BB2XL U2874 ( .B0(n6687), .B1(n286), .A0N(\ram[144][12] ), .A1N(n6466), 
        .Y(n2898) );
  OAI2BB2XL U2875 ( .B0(n6664), .B1(n286), .A0N(\ram[144][13] ), .A1N(n6466), 
        .Y(n2899) );
  OAI2BB2XL U2876 ( .B0(n6641), .B1(n286), .A0N(\ram[144][14] ), .A1N(n6466), 
        .Y(n2900) );
  OAI2BB2XL U2877 ( .B0(n6618), .B1(n286), .A0N(\ram[144][15] ), .A1N(n6466), 
        .Y(n2901) );
  OAI2BB2XL U2878 ( .B0(n6968), .B1(n288), .A0N(\ram[145][0] ), .A1N(n6465), 
        .Y(n2902) );
  OAI2BB2XL U2879 ( .B0(n6945), .B1(n288), .A0N(\ram[145][1] ), .A1N(n6465), 
        .Y(n2903) );
  OAI2BB2XL U2880 ( .B0(n6922), .B1(n288), .A0N(\ram[145][2] ), .A1N(n6465), 
        .Y(n2904) );
  OAI2BB2XL U2881 ( .B0(n6899), .B1(n288), .A0N(\ram[145][3] ), .A1N(n6465), 
        .Y(n2905) );
  OAI2BB2XL U2882 ( .B0(n6871), .B1(n288), .A0N(\ram[145][4] ), .A1N(n6465), 
        .Y(n2906) );
  OAI2BB2XL U2883 ( .B0(n6848), .B1(n288), .A0N(\ram[145][5] ), .A1N(n6465), 
        .Y(n2907) );
  OAI2BB2XL U2884 ( .B0(n6825), .B1(n288), .A0N(\ram[145][6] ), .A1N(n6465), 
        .Y(n2908) );
  OAI2BB2XL U2885 ( .B0(n6802), .B1(n288), .A0N(\ram[145][7] ), .A1N(n6465), 
        .Y(n2909) );
  OAI2BB2XL U2886 ( .B0(n6779), .B1(n288), .A0N(\ram[145][8] ), .A1N(n6465), 
        .Y(n2910) );
  OAI2BB2XL U2887 ( .B0(n6756), .B1(n288), .A0N(\ram[145][9] ), .A1N(n6465), 
        .Y(n2911) );
  OAI2BB2XL U2888 ( .B0(n6733), .B1(n288), .A0N(\ram[145][10] ), .A1N(n6465), 
        .Y(n2912) );
  OAI2BB2XL U2889 ( .B0(n6710), .B1(n288), .A0N(\ram[145][11] ), .A1N(n6465), 
        .Y(n2913) );
  OAI2BB2XL U2890 ( .B0(n6687), .B1(n288), .A0N(\ram[145][12] ), .A1N(n6465), 
        .Y(n2914) );
  OAI2BB2XL U2891 ( .B0(n6664), .B1(n288), .A0N(\ram[145][13] ), .A1N(n6465), 
        .Y(n2915) );
  OAI2BB2XL U2892 ( .B0(n6641), .B1(n288), .A0N(\ram[145][14] ), .A1N(n6465), 
        .Y(n2916) );
  OAI2BB2XL U2893 ( .B0(n6618), .B1(n288), .A0N(\ram[145][15] ), .A1N(n6465), 
        .Y(n2917) );
  OAI2BB2XL U2894 ( .B0(n6968), .B1(n290), .A0N(\ram[146][0] ), .A1N(n6464), 
        .Y(n2918) );
  OAI2BB2XL U2895 ( .B0(n6945), .B1(n290), .A0N(\ram[146][1] ), .A1N(n6464), 
        .Y(n2919) );
  OAI2BB2XL U2896 ( .B0(n6922), .B1(n290), .A0N(\ram[146][2] ), .A1N(n6464), 
        .Y(n2920) );
  OAI2BB2XL U2897 ( .B0(n6899), .B1(n290), .A0N(\ram[146][3] ), .A1N(n6464), 
        .Y(n2921) );
  OAI2BB2XL U2898 ( .B0(n6871), .B1(n290), .A0N(\ram[146][4] ), .A1N(n6464), 
        .Y(n2922) );
  OAI2BB2XL U2899 ( .B0(n6848), .B1(n290), .A0N(\ram[146][5] ), .A1N(n6464), 
        .Y(n2923) );
  OAI2BB2XL U2900 ( .B0(n6825), .B1(n290), .A0N(\ram[146][6] ), .A1N(n6464), 
        .Y(n2924) );
  OAI2BB2XL U2901 ( .B0(n6802), .B1(n290), .A0N(\ram[146][7] ), .A1N(n6464), 
        .Y(n2925) );
  OAI2BB2XL U2902 ( .B0(n6779), .B1(n290), .A0N(\ram[146][8] ), .A1N(n6464), 
        .Y(n2926) );
  OAI2BB2XL U2903 ( .B0(n6756), .B1(n290), .A0N(\ram[146][9] ), .A1N(n6464), 
        .Y(n2927) );
  OAI2BB2XL U2904 ( .B0(n6733), .B1(n290), .A0N(\ram[146][10] ), .A1N(n6464), 
        .Y(n2928) );
  OAI2BB2XL U2905 ( .B0(n6710), .B1(n290), .A0N(\ram[146][11] ), .A1N(n6464), 
        .Y(n2929) );
  OAI2BB2XL U2906 ( .B0(n6687), .B1(n290), .A0N(\ram[146][12] ), .A1N(n6464), 
        .Y(n2930) );
  OAI2BB2XL U2907 ( .B0(n6664), .B1(n290), .A0N(\ram[146][13] ), .A1N(n6464), 
        .Y(n2931) );
  OAI2BB2XL U2908 ( .B0(n6641), .B1(n290), .A0N(\ram[146][14] ), .A1N(n6464), 
        .Y(n2932) );
  OAI2BB2XL U2909 ( .B0(n6618), .B1(n290), .A0N(\ram[146][15] ), .A1N(n6464), 
        .Y(n2933) );
  OAI2BB2XL U2910 ( .B0(n6968), .B1(n292), .A0N(\ram[147][0] ), .A1N(n6463), 
        .Y(n2934) );
  OAI2BB2XL U2911 ( .B0(n6945), .B1(n292), .A0N(\ram[147][1] ), .A1N(n6463), 
        .Y(n2935) );
  OAI2BB2XL U2912 ( .B0(n6922), .B1(n292), .A0N(\ram[147][2] ), .A1N(n6463), 
        .Y(n2936) );
  OAI2BB2XL U2913 ( .B0(n6899), .B1(n292), .A0N(\ram[147][3] ), .A1N(n6463), 
        .Y(n2937) );
  OAI2BB2XL U2914 ( .B0(n6871), .B1(n292), .A0N(\ram[147][4] ), .A1N(n6463), 
        .Y(n2938) );
  OAI2BB2XL U2915 ( .B0(n6848), .B1(n292), .A0N(\ram[147][5] ), .A1N(n6463), 
        .Y(n2939) );
  OAI2BB2XL U2916 ( .B0(n6825), .B1(n292), .A0N(\ram[147][6] ), .A1N(n6463), 
        .Y(n2940) );
  OAI2BB2XL U2917 ( .B0(n6802), .B1(n292), .A0N(\ram[147][7] ), .A1N(n6463), 
        .Y(n2941) );
  OAI2BB2XL U2918 ( .B0(n6779), .B1(n292), .A0N(\ram[147][8] ), .A1N(n6463), 
        .Y(n2942) );
  OAI2BB2XL U2919 ( .B0(n6756), .B1(n292), .A0N(\ram[147][9] ), .A1N(n6463), 
        .Y(n2943) );
  OAI2BB2XL U2920 ( .B0(n6733), .B1(n292), .A0N(\ram[147][10] ), .A1N(n6463), 
        .Y(n2944) );
  OAI2BB2XL U2921 ( .B0(n6710), .B1(n292), .A0N(\ram[147][11] ), .A1N(n6463), 
        .Y(n2945) );
  OAI2BB2XL U2922 ( .B0(n6687), .B1(n292), .A0N(\ram[147][12] ), .A1N(n6463), 
        .Y(n2946) );
  OAI2BB2XL U2923 ( .B0(n6664), .B1(n292), .A0N(\ram[147][13] ), .A1N(n6463), 
        .Y(n2947) );
  OAI2BB2XL U2924 ( .B0(n6641), .B1(n292), .A0N(\ram[147][14] ), .A1N(n6463), 
        .Y(n2948) );
  OAI2BB2XL U2925 ( .B0(n6618), .B1(n292), .A0N(\ram[147][15] ), .A1N(n6463), 
        .Y(n2949) );
  OAI2BB2XL U2926 ( .B0(n6967), .B1(n294), .A0N(\ram[148][0] ), .A1N(n6462), 
        .Y(n2950) );
  OAI2BB2XL U2927 ( .B0(n6944), .B1(n294), .A0N(\ram[148][1] ), .A1N(n6462), 
        .Y(n2951) );
  OAI2BB2XL U2928 ( .B0(n6921), .B1(n294), .A0N(\ram[148][2] ), .A1N(n6462), 
        .Y(n2952) );
  OAI2BB2XL U2929 ( .B0(n6898), .B1(n294), .A0N(\ram[148][3] ), .A1N(n6462), 
        .Y(n2953) );
  OAI2BB2XL U2930 ( .B0(n6870), .B1(n294), .A0N(\ram[148][4] ), .A1N(n6462), 
        .Y(n2954) );
  OAI2BB2XL U2931 ( .B0(n6847), .B1(n294), .A0N(\ram[148][5] ), .A1N(n6462), 
        .Y(n2955) );
  OAI2BB2XL U2932 ( .B0(n6824), .B1(n294), .A0N(\ram[148][6] ), .A1N(n6462), 
        .Y(n2956) );
  OAI2BB2XL U2933 ( .B0(n6801), .B1(n294), .A0N(\ram[148][7] ), .A1N(n6462), 
        .Y(n2957) );
  OAI2BB2XL U2934 ( .B0(n6778), .B1(n294), .A0N(\ram[148][8] ), .A1N(n6462), 
        .Y(n2958) );
  OAI2BB2XL U2935 ( .B0(n6755), .B1(n294), .A0N(\ram[148][9] ), .A1N(n6462), 
        .Y(n2959) );
  OAI2BB2XL U2936 ( .B0(n6732), .B1(n294), .A0N(\ram[148][10] ), .A1N(n6462), 
        .Y(n2960) );
  OAI2BB2XL U2937 ( .B0(n6709), .B1(n294), .A0N(\ram[148][11] ), .A1N(n6462), 
        .Y(n2961) );
  OAI2BB2XL U2938 ( .B0(n6686), .B1(n294), .A0N(\ram[148][12] ), .A1N(n6462), 
        .Y(n2962) );
  OAI2BB2XL U2939 ( .B0(n6663), .B1(n294), .A0N(\ram[148][13] ), .A1N(n6462), 
        .Y(n2963) );
  OAI2BB2XL U2940 ( .B0(n6640), .B1(n294), .A0N(\ram[148][14] ), .A1N(n6462), 
        .Y(n2964) );
  OAI2BB2XL U2941 ( .B0(n6617), .B1(n294), .A0N(\ram[148][15] ), .A1N(n6462), 
        .Y(n2965) );
  OAI2BB2XL U2942 ( .B0(n6967), .B1(n506), .A0N(\ram[149][0] ), .A1N(n6461), 
        .Y(n2966) );
  OAI2BB2XL U2943 ( .B0(n6944), .B1(n506), .A0N(\ram[149][1] ), .A1N(n6461), 
        .Y(n2967) );
  OAI2BB2XL U2944 ( .B0(n6921), .B1(n506), .A0N(\ram[149][2] ), .A1N(n6461), 
        .Y(n2968) );
  OAI2BB2XL U2945 ( .B0(n6898), .B1(n506), .A0N(\ram[149][3] ), .A1N(n6461), 
        .Y(n2969) );
  OAI2BB2XL U2946 ( .B0(n6870), .B1(n506), .A0N(\ram[149][4] ), .A1N(n6461), 
        .Y(n2970) );
  OAI2BB2XL U2947 ( .B0(n6847), .B1(n506), .A0N(\ram[149][5] ), .A1N(n6461), 
        .Y(n2971) );
  OAI2BB2XL U2948 ( .B0(n6824), .B1(n506), .A0N(\ram[149][6] ), .A1N(n6461), 
        .Y(n2972) );
  OAI2BB2XL U2949 ( .B0(n6801), .B1(n506), .A0N(\ram[149][7] ), .A1N(n6461), 
        .Y(n2973) );
  OAI2BB2XL U2950 ( .B0(n6778), .B1(n506), .A0N(\ram[149][8] ), .A1N(n6461), 
        .Y(n2974) );
  OAI2BB2XL U2951 ( .B0(n6755), .B1(n506), .A0N(\ram[149][9] ), .A1N(n6461), 
        .Y(n2975) );
  OAI2BB2XL U2952 ( .B0(n6732), .B1(n506), .A0N(\ram[149][10] ), .A1N(n6461), 
        .Y(n2976) );
  OAI2BB2XL U2953 ( .B0(n6709), .B1(n506), .A0N(\ram[149][11] ), .A1N(n6461), 
        .Y(n2977) );
  OAI2BB2XL U2954 ( .B0(n6686), .B1(n506), .A0N(\ram[149][12] ), .A1N(n6461), 
        .Y(n2978) );
  OAI2BB2XL U2955 ( .B0(n6663), .B1(n506), .A0N(\ram[149][13] ), .A1N(n6461), 
        .Y(n2979) );
  OAI2BB2XL U2956 ( .B0(n6640), .B1(n506), .A0N(\ram[149][14] ), .A1N(n6461), 
        .Y(n2980) );
  OAI2BB2XL U2957 ( .B0(n6617), .B1(n506), .A0N(\ram[149][15] ), .A1N(n6461), 
        .Y(n2981) );
  OAI2BB2XL U2958 ( .B0(n6967), .B1(n508), .A0N(\ram[150][0] ), .A1N(n6460), 
        .Y(n2982) );
  OAI2BB2XL U2959 ( .B0(n6944), .B1(n508), .A0N(\ram[150][1] ), .A1N(n6460), 
        .Y(n2983) );
  OAI2BB2XL U2960 ( .B0(n6921), .B1(n508), .A0N(\ram[150][2] ), .A1N(n6460), 
        .Y(n2984) );
  OAI2BB2XL U2961 ( .B0(n6898), .B1(n508), .A0N(\ram[150][3] ), .A1N(n6460), 
        .Y(n2985) );
  OAI2BB2XL U2962 ( .B0(n6870), .B1(n508), .A0N(\ram[150][4] ), .A1N(n6460), 
        .Y(n2986) );
  OAI2BB2XL U2963 ( .B0(n6847), .B1(n508), .A0N(\ram[150][5] ), .A1N(n6460), 
        .Y(n2987) );
  OAI2BB2XL U2964 ( .B0(n6824), .B1(n508), .A0N(\ram[150][6] ), .A1N(n6460), 
        .Y(n2988) );
  OAI2BB2XL U2965 ( .B0(n6801), .B1(n508), .A0N(\ram[150][7] ), .A1N(n6460), 
        .Y(n2989) );
  OAI2BB2XL U2966 ( .B0(n6778), .B1(n508), .A0N(\ram[150][8] ), .A1N(n6460), 
        .Y(n2990) );
  OAI2BB2XL U2967 ( .B0(n6755), .B1(n508), .A0N(\ram[150][9] ), .A1N(n6460), 
        .Y(n2991) );
  OAI2BB2XL U2968 ( .B0(n6732), .B1(n508), .A0N(\ram[150][10] ), .A1N(n6460), 
        .Y(n2992) );
  OAI2BB2XL U2969 ( .B0(n6709), .B1(n508), .A0N(\ram[150][11] ), .A1N(n6460), 
        .Y(n2993) );
  OAI2BB2XL U2970 ( .B0(n6686), .B1(n508), .A0N(\ram[150][12] ), .A1N(n6460), 
        .Y(n2994) );
  OAI2BB2XL U2971 ( .B0(n6663), .B1(n508), .A0N(\ram[150][13] ), .A1N(n6460), 
        .Y(n2995) );
  OAI2BB2XL U2972 ( .B0(n6640), .B1(n508), .A0N(\ram[150][14] ), .A1N(n6460), 
        .Y(n2996) );
  OAI2BB2XL U2973 ( .B0(n6617), .B1(n508), .A0N(\ram[150][15] ), .A1N(n6460), 
        .Y(n2997) );
  OAI2BB2XL U2974 ( .B0(n6967), .B1(n510), .A0N(\ram[151][0] ), .A1N(n6459), 
        .Y(n2998) );
  OAI2BB2XL U2975 ( .B0(n6944), .B1(n510), .A0N(\ram[151][1] ), .A1N(n6459), 
        .Y(n2999) );
  OAI2BB2XL U2976 ( .B0(n6921), .B1(n510), .A0N(\ram[151][2] ), .A1N(n6459), 
        .Y(n3000) );
  OAI2BB2XL U2977 ( .B0(n6898), .B1(n510), .A0N(\ram[151][3] ), .A1N(n6459), 
        .Y(n3001) );
  OAI2BB2XL U2978 ( .B0(n6870), .B1(n510), .A0N(\ram[151][4] ), .A1N(n6459), 
        .Y(n3002) );
  OAI2BB2XL U2979 ( .B0(n6847), .B1(n510), .A0N(\ram[151][5] ), .A1N(n6459), 
        .Y(n3003) );
  OAI2BB2XL U2980 ( .B0(n6824), .B1(n510), .A0N(\ram[151][6] ), .A1N(n6459), 
        .Y(n3004) );
  OAI2BB2XL U2981 ( .B0(n6801), .B1(n510), .A0N(\ram[151][7] ), .A1N(n6459), 
        .Y(n3005) );
  OAI2BB2XL U2982 ( .B0(n6778), .B1(n510), .A0N(\ram[151][8] ), .A1N(n6459), 
        .Y(n3006) );
  OAI2BB2XL U2983 ( .B0(n6755), .B1(n510), .A0N(\ram[151][9] ), .A1N(n6459), 
        .Y(n3007) );
  OAI2BB2XL U2984 ( .B0(n6732), .B1(n510), .A0N(\ram[151][10] ), .A1N(n6459), 
        .Y(n3008) );
  OAI2BB2XL U2985 ( .B0(n6709), .B1(n510), .A0N(\ram[151][11] ), .A1N(n6459), 
        .Y(n3009) );
  OAI2BB2XL U2986 ( .B0(n6686), .B1(n510), .A0N(\ram[151][12] ), .A1N(n6459), 
        .Y(n3010) );
  OAI2BB2XL U2987 ( .B0(n6663), .B1(n510), .A0N(\ram[151][13] ), .A1N(n6459), 
        .Y(n3011) );
  OAI2BB2XL U2988 ( .B0(n6640), .B1(n510), .A0N(\ram[151][14] ), .A1N(n6459), 
        .Y(n3012) );
  OAI2BB2XL U2989 ( .B0(n6617), .B1(n510), .A0N(\ram[151][15] ), .A1N(n6459), 
        .Y(n3013) );
  OAI2BB2XL U2990 ( .B0(n6967), .B1(n296), .A0N(\ram[152][0] ), .A1N(n6458), 
        .Y(n3014) );
  OAI2BB2XL U2991 ( .B0(n6944), .B1(n296), .A0N(\ram[152][1] ), .A1N(n6458), 
        .Y(n3015) );
  OAI2BB2XL U2992 ( .B0(n6921), .B1(n296), .A0N(\ram[152][2] ), .A1N(n6458), 
        .Y(n3016) );
  OAI2BB2XL U2993 ( .B0(n6898), .B1(n296), .A0N(\ram[152][3] ), .A1N(n6458), 
        .Y(n3017) );
  OAI2BB2XL U2994 ( .B0(n6870), .B1(n296), .A0N(\ram[152][4] ), .A1N(n6458), 
        .Y(n3018) );
  OAI2BB2XL U2995 ( .B0(n6847), .B1(n296), .A0N(\ram[152][5] ), .A1N(n6458), 
        .Y(n3019) );
  OAI2BB2XL U2996 ( .B0(n6824), .B1(n296), .A0N(\ram[152][6] ), .A1N(n6458), 
        .Y(n3020) );
  OAI2BB2XL U2997 ( .B0(n6801), .B1(n296), .A0N(\ram[152][7] ), .A1N(n6458), 
        .Y(n3021) );
  OAI2BB2XL U2998 ( .B0(n6778), .B1(n296), .A0N(\ram[152][8] ), .A1N(n6458), 
        .Y(n3022) );
  OAI2BB2XL U2999 ( .B0(n6755), .B1(n296), .A0N(\ram[152][9] ), .A1N(n6458), 
        .Y(n3023) );
  OAI2BB2XL U3000 ( .B0(n6732), .B1(n296), .A0N(\ram[152][10] ), .A1N(n6458), 
        .Y(n3024) );
  OAI2BB2XL U3001 ( .B0(n6709), .B1(n296), .A0N(\ram[152][11] ), .A1N(n6458), 
        .Y(n3025) );
  OAI2BB2XL U3002 ( .B0(n6686), .B1(n296), .A0N(\ram[152][12] ), .A1N(n6458), 
        .Y(n3026) );
  OAI2BB2XL U3003 ( .B0(n6663), .B1(n296), .A0N(\ram[152][13] ), .A1N(n6458), 
        .Y(n3027) );
  OAI2BB2XL U3004 ( .B0(n6640), .B1(n296), .A0N(\ram[152][14] ), .A1N(n6458), 
        .Y(n3028) );
  OAI2BB2XL U3005 ( .B0(n6617), .B1(n296), .A0N(\ram[152][15] ), .A1N(n6458), 
        .Y(n3029) );
  OAI2BB2XL U3006 ( .B0(n6967), .B1(n298), .A0N(\ram[153][0] ), .A1N(n6457), 
        .Y(n3030) );
  OAI2BB2XL U3007 ( .B0(n6944), .B1(n298), .A0N(\ram[153][1] ), .A1N(n6457), 
        .Y(n3031) );
  OAI2BB2XL U3008 ( .B0(n6921), .B1(n298), .A0N(\ram[153][2] ), .A1N(n6457), 
        .Y(n3032) );
  OAI2BB2XL U3009 ( .B0(n6898), .B1(n298), .A0N(\ram[153][3] ), .A1N(n6457), 
        .Y(n3033) );
  OAI2BB2XL U3010 ( .B0(n6870), .B1(n298), .A0N(\ram[153][4] ), .A1N(n6457), 
        .Y(n3034) );
  OAI2BB2XL U3011 ( .B0(n6847), .B1(n298), .A0N(\ram[153][5] ), .A1N(n6457), 
        .Y(n3035) );
  OAI2BB2XL U3012 ( .B0(n6824), .B1(n298), .A0N(\ram[153][6] ), .A1N(n6457), 
        .Y(n3036) );
  OAI2BB2XL U3013 ( .B0(n6801), .B1(n298), .A0N(\ram[153][7] ), .A1N(n6457), 
        .Y(n3037) );
  OAI2BB2XL U3014 ( .B0(n6778), .B1(n298), .A0N(\ram[153][8] ), .A1N(n6457), 
        .Y(n3038) );
  OAI2BB2XL U3015 ( .B0(n6755), .B1(n298), .A0N(\ram[153][9] ), .A1N(n6457), 
        .Y(n3039) );
  OAI2BB2XL U3016 ( .B0(n6732), .B1(n298), .A0N(\ram[153][10] ), .A1N(n6457), 
        .Y(n3040) );
  OAI2BB2XL U3017 ( .B0(n6709), .B1(n298), .A0N(\ram[153][11] ), .A1N(n6457), 
        .Y(n3041) );
  OAI2BB2XL U3018 ( .B0(n6686), .B1(n298), .A0N(\ram[153][12] ), .A1N(n6457), 
        .Y(n3042) );
  OAI2BB2XL U3019 ( .B0(n6663), .B1(n298), .A0N(\ram[153][13] ), .A1N(n6457), 
        .Y(n3043) );
  OAI2BB2XL U3020 ( .B0(n6640), .B1(n298), .A0N(\ram[153][14] ), .A1N(n6457), 
        .Y(n3044) );
  OAI2BB2XL U3021 ( .B0(n6617), .B1(n298), .A0N(\ram[153][15] ), .A1N(n6457), 
        .Y(n3045) );
  OAI2BB2XL U3022 ( .B0(n6967), .B1(n300), .A0N(\ram[154][0] ), .A1N(n6456), 
        .Y(n3046) );
  OAI2BB2XL U3023 ( .B0(n6944), .B1(n300), .A0N(\ram[154][1] ), .A1N(n6456), 
        .Y(n3047) );
  OAI2BB2XL U3024 ( .B0(n6921), .B1(n300), .A0N(\ram[154][2] ), .A1N(n6456), 
        .Y(n3048) );
  OAI2BB2XL U3025 ( .B0(n6898), .B1(n300), .A0N(\ram[154][3] ), .A1N(n6456), 
        .Y(n3049) );
  OAI2BB2XL U3026 ( .B0(n6870), .B1(n300), .A0N(\ram[154][4] ), .A1N(n6456), 
        .Y(n3050) );
  OAI2BB2XL U3027 ( .B0(n6847), .B1(n300), .A0N(\ram[154][5] ), .A1N(n6456), 
        .Y(n3051) );
  OAI2BB2XL U3028 ( .B0(n6824), .B1(n300), .A0N(\ram[154][6] ), .A1N(n6456), 
        .Y(n3052) );
  OAI2BB2XL U3029 ( .B0(n6801), .B1(n300), .A0N(\ram[154][7] ), .A1N(n6456), 
        .Y(n3053) );
  OAI2BB2XL U3030 ( .B0(n6778), .B1(n300), .A0N(\ram[154][8] ), .A1N(n6456), 
        .Y(n3054) );
  OAI2BB2XL U3031 ( .B0(n6755), .B1(n300), .A0N(\ram[154][9] ), .A1N(n6456), 
        .Y(n3055) );
  OAI2BB2XL U3032 ( .B0(n6732), .B1(n300), .A0N(\ram[154][10] ), .A1N(n6456), 
        .Y(n3056) );
  OAI2BB2XL U3033 ( .B0(n6709), .B1(n300), .A0N(\ram[154][11] ), .A1N(n6456), 
        .Y(n3057) );
  OAI2BB2XL U3034 ( .B0(n6686), .B1(n300), .A0N(\ram[154][12] ), .A1N(n6456), 
        .Y(n3058) );
  OAI2BB2XL U3035 ( .B0(n6663), .B1(n300), .A0N(\ram[154][13] ), .A1N(n6456), 
        .Y(n3059) );
  OAI2BB2XL U3036 ( .B0(n6640), .B1(n300), .A0N(\ram[154][14] ), .A1N(n6456), 
        .Y(n3060) );
  OAI2BB2XL U3037 ( .B0(n6617), .B1(n300), .A0N(\ram[154][15] ), .A1N(n6456), 
        .Y(n3061) );
  OAI2BB2XL U3038 ( .B0(n6967), .B1(n302), .A0N(\ram[155][0] ), .A1N(n6455), 
        .Y(n3062) );
  OAI2BB2XL U3039 ( .B0(n6944), .B1(n302), .A0N(\ram[155][1] ), .A1N(n6455), 
        .Y(n3063) );
  OAI2BB2XL U3040 ( .B0(n6921), .B1(n302), .A0N(\ram[155][2] ), .A1N(n6455), 
        .Y(n3064) );
  OAI2BB2XL U3041 ( .B0(n6898), .B1(n302), .A0N(\ram[155][3] ), .A1N(n6455), 
        .Y(n3065) );
  OAI2BB2XL U3042 ( .B0(n6870), .B1(n302), .A0N(\ram[155][4] ), .A1N(n6455), 
        .Y(n3066) );
  OAI2BB2XL U3043 ( .B0(n6847), .B1(n302), .A0N(\ram[155][5] ), .A1N(n6455), 
        .Y(n3067) );
  OAI2BB2XL U3044 ( .B0(n6824), .B1(n302), .A0N(\ram[155][6] ), .A1N(n6455), 
        .Y(n3068) );
  OAI2BB2XL U3045 ( .B0(n6801), .B1(n302), .A0N(\ram[155][7] ), .A1N(n6455), 
        .Y(n3069) );
  OAI2BB2XL U3046 ( .B0(n6778), .B1(n302), .A0N(\ram[155][8] ), .A1N(n6455), 
        .Y(n3070) );
  OAI2BB2XL U3047 ( .B0(n6755), .B1(n302), .A0N(\ram[155][9] ), .A1N(n6455), 
        .Y(n3071) );
  OAI2BB2XL U3048 ( .B0(n6732), .B1(n302), .A0N(\ram[155][10] ), .A1N(n6455), 
        .Y(n3072) );
  OAI2BB2XL U3049 ( .B0(n6709), .B1(n302), .A0N(\ram[155][11] ), .A1N(n6455), 
        .Y(n3073) );
  OAI2BB2XL U3050 ( .B0(n6686), .B1(n302), .A0N(\ram[155][12] ), .A1N(n6455), 
        .Y(n3074) );
  OAI2BB2XL U3051 ( .B0(n6663), .B1(n302), .A0N(\ram[155][13] ), .A1N(n6455), 
        .Y(n3075) );
  OAI2BB2XL U3052 ( .B0(n6640), .B1(n302), .A0N(\ram[155][14] ), .A1N(n6455), 
        .Y(n3076) );
  OAI2BB2XL U3053 ( .B0(n6617), .B1(n302), .A0N(\ram[155][15] ), .A1N(n6455), 
        .Y(n3077) );
  OAI2BB2XL U3054 ( .B0(n6967), .B1(n304), .A0N(\ram[156][0] ), .A1N(n6454), 
        .Y(n3078) );
  OAI2BB2XL U3055 ( .B0(n6944), .B1(n304), .A0N(\ram[156][1] ), .A1N(n6454), 
        .Y(n3079) );
  OAI2BB2XL U3056 ( .B0(n6921), .B1(n304), .A0N(\ram[156][2] ), .A1N(n6454), 
        .Y(n3080) );
  OAI2BB2XL U3057 ( .B0(n6898), .B1(n304), .A0N(\ram[156][3] ), .A1N(n6454), 
        .Y(n3081) );
  OAI2BB2XL U3058 ( .B0(n6870), .B1(n304), .A0N(\ram[156][4] ), .A1N(n6454), 
        .Y(n3082) );
  OAI2BB2XL U3059 ( .B0(n6847), .B1(n304), .A0N(\ram[156][5] ), .A1N(n6454), 
        .Y(n3083) );
  OAI2BB2XL U3060 ( .B0(n6824), .B1(n304), .A0N(\ram[156][6] ), .A1N(n6454), 
        .Y(n3084) );
  OAI2BB2XL U3061 ( .B0(n6801), .B1(n304), .A0N(\ram[156][7] ), .A1N(n6454), 
        .Y(n3085) );
  OAI2BB2XL U3062 ( .B0(n6778), .B1(n304), .A0N(\ram[156][8] ), .A1N(n6454), 
        .Y(n3086) );
  OAI2BB2XL U3063 ( .B0(n6755), .B1(n304), .A0N(\ram[156][9] ), .A1N(n6454), 
        .Y(n3087) );
  OAI2BB2XL U3064 ( .B0(n6732), .B1(n304), .A0N(\ram[156][10] ), .A1N(n6454), 
        .Y(n3088) );
  OAI2BB2XL U3065 ( .B0(n6709), .B1(n304), .A0N(\ram[156][11] ), .A1N(n6454), 
        .Y(n3089) );
  OAI2BB2XL U3066 ( .B0(n6686), .B1(n304), .A0N(\ram[156][12] ), .A1N(n6454), 
        .Y(n3090) );
  OAI2BB2XL U3067 ( .B0(n6663), .B1(n304), .A0N(\ram[156][13] ), .A1N(n6454), 
        .Y(n3091) );
  OAI2BB2XL U3068 ( .B0(n6640), .B1(n304), .A0N(\ram[156][14] ), .A1N(n6454), 
        .Y(n3092) );
  OAI2BB2XL U3069 ( .B0(n6617), .B1(n304), .A0N(\ram[156][15] ), .A1N(n6454), 
        .Y(n3093) );
  OAI2BB2XL U3070 ( .B0(n6967), .B1(n306), .A0N(\ram[157][0] ), .A1N(n6453), 
        .Y(n3094) );
  OAI2BB2XL U3071 ( .B0(n6944), .B1(n306), .A0N(\ram[157][1] ), .A1N(n6453), 
        .Y(n3095) );
  OAI2BB2XL U3072 ( .B0(n6921), .B1(n306), .A0N(\ram[157][2] ), .A1N(n6453), 
        .Y(n3096) );
  OAI2BB2XL U3073 ( .B0(n6898), .B1(n306), .A0N(\ram[157][3] ), .A1N(n6453), 
        .Y(n3097) );
  OAI2BB2XL U3074 ( .B0(n6870), .B1(n306), .A0N(\ram[157][4] ), .A1N(n6453), 
        .Y(n3098) );
  OAI2BB2XL U3075 ( .B0(n6847), .B1(n306), .A0N(\ram[157][5] ), .A1N(n6453), 
        .Y(n3099) );
  OAI2BB2XL U3076 ( .B0(n6824), .B1(n306), .A0N(\ram[157][6] ), .A1N(n6453), 
        .Y(n3100) );
  OAI2BB2XL U3077 ( .B0(n6801), .B1(n306), .A0N(\ram[157][7] ), .A1N(n6453), 
        .Y(n3101) );
  OAI2BB2XL U3078 ( .B0(n6778), .B1(n306), .A0N(\ram[157][8] ), .A1N(n6453), 
        .Y(n3102) );
  OAI2BB2XL U3079 ( .B0(n6755), .B1(n306), .A0N(\ram[157][9] ), .A1N(n6453), 
        .Y(n3103) );
  OAI2BB2XL U3080 ( .B0(n6732), .B1(n306), .A0N(\ram[157][10] ), .A1N(n6453), 
        .Y(n3104) );
  OAI2BB2XL U3081 ( .B0(n6709), .B1(n306), .A0N(\ram[157][11] ), .A1N(n6453), 
        .Y(n3105) );
  OAI2BB2XL U3082 ( .B0(n6686), .B1(n306), .A0N(\ram[157][12] ), .A1N(n6453), 
        .Y(n3106) );
  OAI2BB2XL U3083 ( .B0(n6663), .B1(n306), .A0N(\ram[157][13] ), .A1N(n6453), 
        .Y(n3107) );
  OAI2BB2XL U3084 ( .B0(n6640), .B1(n306), .A0N(\ram[157][14] ), .A1N(n6453), 
        .Y(n3108) );
  OAI2BB2XL U3085 ( .B0(n6617), .B1(n306), .A0N(\ram[157][15] ), .A1N(n6453), 
        .Y(n3109) );
  OAI2BB2XL U3086 ( .B0(n6967), .B1(n308), .A0N(\ram[158][0] ), .A1N(n6452), 
        .Y(n3110) );
  OAI2BB2XL U3087 ( .B0(n6944), .B1(n308), .A0N(\ram[158][1] ), .A1N(n6452), 
        .Y(n3111) );
  OAI2BB2XL U3088 ( .B0(n6921), .B1(n308), .A0N(\ram[158][2] ), .A1N(n6452), 
        .Y(n3112) );
  OAI2BB2XL U3089 ( .B0(n6898), .B1(n308), .A0N(\ram[158][3] ), .A1N(n6452), 
        .Y(n3113) );
  OAI2BB2XL U3090 ( .B0(n6870), .B1(n308), .A0N(\ram[158][4] ), .A1N(n6452), 
        .Y(n3114) );
  OAI2BB2XL U3091 ( .B0(n6847), .B1(n308), .A0N(\ram[158][5] ), .A1N(n6452), 
        .Y(n3115) );
  OAI2BB2XL U3092 ( .B0(n6824), .B1(n308), .A0N(\ram[158][6] ), .A1N(n6452), 
        .Y(n3116) );
  OAI2BB2XL U3093 ( .B0(n6801), .B1(n308), .A0N(\ram[158][7] ), .A1N(n6452), 
        .Y(n3117) );
  OAI2BB2XL U3094 ( .B0(n6778), .B1(n308), .A0N(\ram[158][8] ), .A1N(n6452), 
        .Y(n3118) );
  OAI2BB2XL U3095 ( .B0(n6755), .B1(n308), .A0N(\ram[158][9] ), .A1N(n6452), 
        .Y(n3119) );
  OAI2BB2XL U3096 ( .B0(n6732), .B1(n308), .A0N(\ram[158][10] ), .A1N(n6452), 
        .Y(n3120) );
  OAI2BB2XL U3097 ( .B0(n6709), .B1(n308), .A0N(\ram[158][11] ), .A1N(n6452), 
        .Y(n3121) );
  OAI2BB2XL U3098 ( .B0(n6686), .B1(n308), .A0N(\ram[158][12] ), .A1N(n6452), 
        .Y(n3122) );
  OAI2BB2XL U3099 ( .B0(n6663), .B1(n308), .A0N(\ram[158][13] ), .A1N(n6452), 
        .Y(n3123) );
  OAI2BB2XL U3100 ( .B0(n6640), .B1(n308), .A0N(\ram[158][14] ), .A1N(n6452), 
        .Y(n3124) );
  OAI2BB2XL U3101 ( .B0(n6617), .B1(n308), .A0N(\ram[158][15] ), .A1N(n6452), 
        .Y(n3125) );
  OAI2BB2XL U3102 ( .B0(n6967), .B1(n310), .A0N(\ram[159][0] ), .A1N(n6451), 
        .Y(n3126) );
  OAI2BB2XL U3103 ( .B0(n6944), .B1(n310), .A0N(\ram[159][1] ), .A1N(n6451), 
        .Y(n3127) );
  OAI2BB2XL U3104 ( .B0(n6921), .B1(n310), .A0N(\ram[159][2] ), .A1N(n6451), 
        .Y(n3128) );
  OAI2BB2XL U3105 ( .B0(n6898), .B1(n310), .A0N(\ram[159][3] ), .A1N(n6451), 
        .Y(n3129) );
  OAI2BB2XL U3106 ( .B0(n6870), .B1(n310), .A0N(\ram[159][4] ), .A1N(n6451), 
        .Y(n3130) );
  OAI2BB2XL U3107 ( .B0(n6847), .B1(n310), .A0N(\ram[159][5] ), .A1N(n6451), 
        .Y(n3131) );
  OAI2BB2XL U3108 ( .B0(n6824), .B1(n310), .A0N(\ram[159][6] ), .A1N(n6451), 
        .Y(n3132) );
  OAI2BB2XL U3109 ( .B0(n6801), .B1(n310), .A0N(\ram[159][7] ), .A1N(n6451), 
        .Y(n3133) );
  OAI2BB2XL U3110 ( .B0(n6778), .B1(n310), .A0N(\ram[159][8] ), .A1N(n6451), 
        .Y(n3134) );
  OAI2BB2XL U3111 ( .B0(n6755), .B1(n310), .A0N(\ram[159][9] ), .A1N(n6451), 
        .Y(n3135) );
  OAI2BB2XL U3112 ( .B0(n6732), .B1(n310), .A0N(\ram[159][10] ), .A1N(n6451), 
        .Y(n3136) );
  OAI2BB2XL U3113 ( .B0(n6709), .B1(n310), .A0N(\ram[159][11] ), .A1N(n6451), 
        .Y(n3137) );
  OAI2BB2XL U3114 ( .B0(n6686), .B1(n310), .A0N(\ram[159][12] ), .A1N(n6451), 
        .Y(n3138) );
  OAI2BB2XL U3115 ( .B0(n6663), .B1(n310), .A0N(\ram[159][13] ), .A1N(n6451), 
        .Y(n3139) );
  OAI2BB2XL U3116 ( .B0(n6640), .B1(n310), .A0N(\ram[159][14] ), .A1N(n6451), 
        .Y(n3140) );
  OAI2BB2XL U3117 ( .B0(n6617), .B1(n310), .A0N(\ram[159][15] ), .A1N(n6451), 
        .Y(n3141) );
  OAI2BB2XL U3118 ( .B0(n6966), .B1(n311), .A0N(\ram[160][0] ), .A1N(n6450), 
        .Y(n3142) );
  OAI2BB2XL U3119 ( .B0(n6943), .B1(n311), .A0N(\ram[160][1] ), .A1N(n6450), 
        .Y(n3143) );
  OAI2BB2XL U3120 ( .B0(n6920), .B1(n311), .A0N(\ram[160][2] ), .A1N(n6450), 
        .Y(n3144) );
  OAI2BB2XL U3121 ( .B0(n6897), .B1(n311), .A0N(\ram[160][3] ), .A1N(n6450), 
        .Y(n3145) );
  OAI2BB2XL U3122 ( .B0(n6869), .B1(n311), .A0N(\ram[160][4] ), .A1N(n6450), 
        .Y(n3146) );
  OAI2BB2XL U3123 ( .B0(n6846), .B1(n311), .A0N(\ram[160][5] ), .A1N(n6450), 
        .Y(n3147) );
  OAI2BB2XL U3124 ( .B0(n6823), .B1(n311), .A0N(\ram[160][6] ), .A1N(n6450), 
        .Y(n3148) );
  OAI2BB2XL U3125 ( .B0(n6800), .B1(n311), .A0N(\ram[160][7] ), .A1N(n6450), 
        .Y(n3149) );
  OAI2BB2XL U3126 ( .B0(n6777), .B1(n311), .A0N(\ram[160][8] ), .A1N(n6450), 
        .Y(n3150) );
  OAI2BB2XL U3127 ( .B0(n6754), .B1(n311), .A0N(\ram[160][9] ), .A1N(n6450), 
        .Y(n3151) );
  OAI2BB2XL U3128 ( .B0(n6731), .B1(n311), .A0N(\ram[160][10] ), .A1N(n6450), 
        .Y(n3152) );
  OAI2BB2XL U3129 ( .B0(n6708), .B1(n311), .A0N(\ram[160][11] ), .A1N(n6450), 
        .Y(n3153) );
  OAI2BB2XL U3130 ( .B0(n6685), .B1(n311), .A0N(\ram[160][12] ), .A1N(n6450), 
        .Y(n3154) );
  OAI2BB2XL U3131 ( .B0(n6662), .B1(n311), .A0N(\ram[160][13] ), .A1N(n6450), 
        .Y(n3155) );
  OAI2BB2XL U3132 ( .B0(n6639), .B1(n311), .A0N(\ram[160][14] ), .A1N(n6450), 
        .Y(n3156) );
  OAI2BB2XL U3133 ( .B0(n6616), .B1(n311), .A0N(\ram[160][15] ), .A1N(n6450), 
        .Y(n3157) );
  OAI2BB2XL U3134 ( .B0(n6966), .B1(n313), .A0N(\ram[161][0] ), .A1N(n6449), 
        .Y(n3158) );
  OAI2BB2XL U3135 ( .B0(n6943), .B1(n313), .A0N(\ram[161][1] ), .A1N(n6449), 
        .Y(n3159) );
  OAI2BB2XL U3136 ( .B0(n6920), .B1(n313), .A0N(\ram[161][2] ), .A1N(n6449), 
        .Y(n3160) );
  OAI2BB2XL U3137 ( .B0(n6897), .B1(n313), .A0N(\ram[161][3] ), .A1N(n6449), 
        .Y(n3161) );
  OAI2BB2XL U3138 ( .B0(n6869), .B1(n313), .A0N(\ram[161][4] ), .A1N(n6449), 
        .Y(n3162) );
  OAI2BB2XL U3139 ( .B0(n6846), .B1(n313), .A0N(\ram[161][5] ), .A1N(n6449), 
        .Y(n3163) );
  OAI2BB2XL U3140 ( .B0(n6823), .B1(n313), .A0N(\ram[161][6] ), .A1N(n6449), 
        .Y(n3164) );
  OAI2BB2XL U3141 ( .B0(n6800), .B1(n313), .A0N(\ram[161][7] ), .A1N(n6449), 
        .Y(n3165) );
  OAI2BB2XL U3142 ( .B0(n6777), .B1(n313), .A0N(\ram[161][8] ), .A1N(n6449), 
        .Y(n3166) );
  OAI2BB2XL U3143 ( .B0(n6754), .B1(n313), .A0N(\ram[161][9] ), .A1N(n6449), 
        .Y(n3167) );
  OAI2BB2XL U3144 ( .B0(n6731), .B1(n313), .A0N(\ram[161][10] ), .A1N(n6449), 
        .Y(n3168) );
  OAI2BB2XL U3145 ( .B0(n6708), .B1(n313), .A0N(\ram[161][11] ), .A1N(n6449), 
        .Y(n3169) );
  OAI2BB2XL U3146 ( .B0(n6685), .B1(n313), .A0N(\ram[161][12] ), .A1N(n6449), 
        .Y(n3170) );
  OAI2BB2XL U3147 ( .B0(n6662), .B1(n313), .A0N(\ram[161][13] ), .A1N(n6449), 
        .Y(n3171) );
  OAI2BB2XL U3148 ( .B0(n6639), .B1(n313), .A0N(\ram[161][14] ), .A1N(n6449), 
        .Y(n3172) );
  OAI2BB2XL U3149 ( .B0(n6616), .B1(n313), .A0N(\ram[161][15] ), .A1N(n6449), 
        .Y(n3173) );
  OAI2BB2XL U3150 ( .B0(n6966), .B1(n315), .A0N(\ram[162][0] ), .A1N(n6448), 
        .Y(n3174) );
  OAI2BB2XL U3151 ( .B0(n6943), .B1(n315), .A0N(\ram[162][1] ), .A1N(n6448), 
        .Y(n3175) );
  OAI2BB2XL U3152 ( .B0(n6920), .B1(n315), .A0N(\ram[162][2] ), .A1N(n6448), 
        .Y(n3176) );
  OAI2BB2XL U3153 ( .B0(n6897), .B1(n315), .A0N(\ram[162][3] ), .A1N(n6448), 
        .Y(n3177) );
  OAI2BB2XL U3154 ( .B0(n6869), .B1(n315), .A0N(\ram[162][4] ), .A1N(n6448), 
        .Y(n3178) );
  OAI2BB2XL U3155 ( .B0(n6846), .B1(n315), .A0N(\ram[162][5] ), .A1N(n6448), 
        .Y(n3179) );
  OAI2BB2XL U3156 ( .B0(n6823), .B1(n315), .A0N(\ram[162][6] ), .A1N(n6448), 
        .Y(n3180) );
  OAI2BB2XL U3157 ( .B0(n6800), .B1(n315), .A0N(\ram[162][7] ), .A1N(n6448), 
        .Y(n3181) );
  OAI2BB2XL U3158 ( .B0(n6777), .B1(n315), .A0N(\ram[162][8] ), .A1N(n6448), 
        .Y(n3182) );
  OAI2BB2XL U3159 ( .B0(n6754), .B1(n315), .A0N(\ram[162][9] ), .A1N(n6448), 
        .Y(n3183) );
  OAI2BB2XL U3160 ( .B0(n6731), .B1(n315), .A0N(\ram[162][10] ), .A1N(n6448), 
        .Y(n3184) );
  OAI2BB2XL U3161 ( .B0(n6708), .B1(n315), .A0N(\ram[162][11] ), .A1N(n6448), 
        .Y(n3185) );
  OAI2BB2XL U3162 ( .B0(n6685), .B1(n315), .A0N(\ram[162][12] ), .A1N(n6448), 
        .Y(n3186) );
  OAI2BB2XL U3163 ( .B0(n6662), .B1(n315), .A0N(\ram[162][13] ), .A1N(n6448), 
        .Y(n3187) );
  OAI2BB2XL U3164 ( .B0(n6639), .B1(n315), .A0N(\ram[162][14] ), .A1N(n6448), 
        .Y(n3188) );
  OAI2BB2XL U3165 ( .B0(n6616), .B1(n315), .A0N(\ram[162][15] ), .A1N(n6448), 
        .Y(n3189) );
  OAI2BB2XL U3166 ( .B0(n6966), .B1(n317), .A0N(\ram[163][0] ), .A1N(n6447), 
        .Y(n3190) );
  OAI2BB2XL U3167 ( .B0(n6943), .B1(n317), .A0N(\ram[163][1] ), .A1N(n6447), 
        .Y(n3191) );
  OAI2BB2XL U3168 ( .B0(n6920), .B1(n317), .A0N(\ram[163][2] ), .A1N(n6447), 
        .Y(n3192) );
  OAI2BB2XL U3169 ( .B0(n6897), .B1(n317), .A0N(\ram[163][3] ), .A1N(n6447), 
        .Y(n3193) );
  OAI2BB2XL U3170 ( .B0(n6869), .B1(n317), .A0N(\ram[163][4] ), .A1N(n6447), 
        .Y(n3194) );
  OAI2BB2XL U3171 ( .B0(n6846), .B1(n317), .A0N(\ram[163][5] ), .A1N(n6447), 
        .Y(n3195) );
  OAI2BB2XL U3172 ( .B0(n6823), .B1(n317), .A0N(\ram[163][6] ), .A1N(n6447), 
        .Y(n3196) );
  OAI2BB2XL U3173 ( .B0(n6800), .B1(n317), .A0N(\ram[163][7] ), .A1N(n6447), 
        .Y(n3197) );
  OAI2BB2XL U3174 ( .B0(n6777), .B1(n317), .A0N(\ram[163][8] ), .A1N(n6447), 
        .Y(n3198) );
  OAI2BB2XL U3175 ( .B0(n6754), .B1(n317), .A0N(\ram[163][9] ), .A1N(n6447), 
        .Y(n3199) );
  OAI2BB2XL U3176 ( .B0(n6731), .B1(n317), .A0N(\ram[163][10] ), .A1N(n6447), 
        .Y(n3200) );
  OAI2BB2XL U3177 ( .B0(n6708), .B1(n317), .A0N(\ram[163][11] ), .A1N(n6447), 
        .Y(n3201) );
  OAI2BB2XL U3178 ( .B0(n6685), .B1(n317), .A0N(\ram[163][12] ), .A1N(n6447), 
        .Y(n3202) );
  OAI2BB2XL U3179 ( .B0(n6662), .B1(n317), .A0N(\ram[163][13] ), .A1N(n6447), 
        .Y(n3203) );
  OAI2BB2XL U3180 ( .B0(n6639), .B1(n317), .A0N(\ram[163][14] ), .A1N(n6447), 
        .Y(n3204) );
  OAI2BB2XL U3181 ( .B0(n6616), .B1(n317), .A0N(\ram[163][15] ), .A1N(n6447), 
        .Y(n3205) );
  OAI2BB2XL U3182 ( .B0(n6966), .B1(n319), .A0N(\ram[164][0] ), .A1N(n6446), 
        .Y(n3206) );
  OAI2BB2XL U3183 ( .B0(n6943), .B1(n319), .A0N(\ram[164][1] ), .A1N(n6446), 
        .Y(n3207) );
  OAI2BB2XL U3184 ( .B0(n6920), .B1(n319), .A0N(\ram[164][2] ), .A1N(n6446), 
        .Y(n3208) );
  OAI2BB2XL U3185 ( .B0(n6897), .B1(n319), .A0N(\ram[164][3] ), .A1N(n6446), 
        .Y(n3209) );
  OAI2BB2XL U3186 ( .B0(n6869), .B1(n319), .A0N(\ram[164][4] ), .A1N(n6446), 
        .Y(n3210) );
  OAI2BB2XL U3187 ( .B0(n6846), .B1(n319), .A0N(\ram[164][5] ), .A1N(n6446), 
        .Y(n3211) );
  OAI2BB2XL U3188 ( .B0(n6823), .B1(n319), .A0N(\ram[164][6] ), .A1N(n6446), 
        .Y(n3212) );
  OAI2BB2XL U3189 ( .B0(n6800), .B1(n319), .A0N(\ram[164][7] ), .A1N(n6446), 
        .Y(n3213) );
  OAI2BB2XL U3190 ( .B0(n6777), .B1(n319), .A0N(\ram[164][8] ), .A1N(n6446), 
        .Y(n3214) );
  OAI2BB2XL U3191 ( .B0(n6754), .B1(n319), .A0N(\ram[164][9] ), .A1N(n6446), 
        .Y(n3215) );
  OAI2BB2XL U3192 ( .B0(n6731), .B1(n319), .A0N(\ram[164][10] ), .A1N(n6446), 
        .Y(n3216) );
  OAI2BB2XL U3193 ( .B0(n6708), .B1(n319), .A0N(\ram[164][11] ), .A1N(n6446), 
        .Y(n3217) );
  OAI2BB2XL U3194 ( .B0(n6685), .B1(n319), .A0N(\ram[164][12] ), .A1N(n6446), 
        .Y(n3218) );
  OAI2BB2XL U3195 ( .B0(n6662), .B1(n319), .A0N(\ram[164][13] ), .A1N(n6446), 
        .Y(n3219) );
  OAI2BB2XL U3196 ( .B0(n6639), .B1(n319), .A0N(\ram[164][14] ), .A1N(n6446), 
        .Y(n3220) );
  OAI2BB2XL U3197 ( .B0(n6616), .B1(n319), .A0N(\ram[164][15] ), .A1N(n6446), 
        .Y(n3221) );
  OAI2BB2XL U3198 ( .B0(n6966), .B1(n549), .A0N(\ram[165][0] ), .A1N(n6445), 
        .Y(n3222) );
  OAI2BB2XL U3199 ( .B0(n6943), .B1(n549), .A0N(\ram[165][1] ), .A1N(n6445), 
        .Y(n3223) );
  OAI2BB2XL U3200 ( .B0(n6920), .B1(n549), .A0N(\ram[165][2] ), .A1N(n6445), 
        .Y(n3224) );
  OAI2BB2XL U3201 ( .B0(n6897), .B1(n549), .A0N(\ram[165][3] ), .A1N(n6445), 
        .Y(n3225) );
  OAI2BB2XL U3202 ( .B0(n6869), .B1(n549), .A0N(\ram[165][4] ), .A1N(n6445), 
        .Y(n3226) );
  OAI2BB2XL U3203 ( .B0(n6846), .B1(n549), .A0N(\ram[165][5] ), .A1N(n6445), 
        .Y(n3227) );
  OAI2BB2XL U3204 ( .B0(n6823), .B1(n549), .A0N(\ram[165][6] ), .A1N(n6445), 
        .Y(n3228) );
  OAI2BB2XL U3205 ( .B0(n6800), .B1(n549), .A0N(\ram[165][7] ), .A1N(n6445), 
        .Y(n3229) );
  OAI2BB2XL U3206 ( .B0(n6777), .B1(n549), .A0N(\ram[165][8] ), .A1N(n6445), 
        .Y(n3230) );
  OAI2BB2XL U3207 ( .B0(n6754), .B1(n549), .A0N(\ram[165][9] ), .A1N(n6445), 
        .Y(n3231) );
  OAI2BB2XL U3208 ( .B0(n6731), .B1(n549), .A0N(\ram[165][10] ), .A1N(n6445), 
        .Y(n3232) );
  OAI2BB2XL U3209 ( .B0(n6708), .B1(n549), .A0N(\ram[165][11] ), .A1N(n6445), 
        .Y(n3233) );
  OAI2BB2XL U3210 ( .B0(n6685), .B1(n549), .A0N(\ram[165][12] ), .A1N(n6445), 
        .Y(n3234) );
  OAI2BB2XL U3211 ( .B0(n6662), .B1(n549), .A0N(\ram[165][13] ), .A1N(n6445), 
        .Y(n3235) );
  OAI2BB2XL U3212 ( .B0(n6639), .B1(n549), .A0N(\ram[165][14] ), .A1N(n6445), 
        .Y(n3236) );
  OAI2BB2XL U3213 ( .B0(n6616), .B1(n549), .A0N(\ram[165][15] ), .A1N(n6445), 
        .Y(n3237) );
  OAI2BB2XL U3214 ( .B0(n6966), .B1(n552), .A0N(\ram[166][0] ), .A1N(n6444), 
        .Y(n3238) );
  OAI2BB2XL U3215 ( .B0(n6943), .B1(n552), .A0N(\ram[166][1] ), .A1N(n6444), 
        .Y(n3239) );
  OAI2BB2XL U3216 ( .B0(n6920), .B1(n552), .A0N(\ram[166][2] ), .A1N(n6444), 
        .Y(n3240) );
  OAI2BB2XL U3217 ( .B0(n6897), .B1(n552), .A0N(\ram[166][3] ), .A1N(n6444), 
        .Y(n3241) );
  OAI2BB2XL U3218 ( .B0(n6869), .B1(n552), .A0N(\ram[166][4] ), .A1N(n6444), 
        .Y(n3242) );
  OAI2BB2XL U3219 ( .B0(n6846), .B1(n552), .A0N(\ram[166][5] ), .A1N(n6444), 
        .Y(n3243) );
  OAI2BB2XL U3220 ( .B0(n6823), .B1(n552), .A0N(\ram[166][6] ), .A1N(n6444), 
        .Y(n3244) );
  OAI2BB2XL U3221 ( .B0(n6800), .B1(n552), .A0N(\ram[166][7] ), .A1N(n6444), 
        .Y(n3245) );
  OAI2BB2XL U3222 ( .B0(n6777), .B1(n552), .A0N(\ram[166][8] ), .A1N(n6444), 
        .Y(n3246) );
  OAI2BB2XL U3223 ( .B0(n6754), .B1(n552), .A0N(\ram[166][9] ), .A1N(n6444), 
        .Y(n3247) );
  OAI2BB2XL U3224 ( .B0(n6731), .B1(n552), .A0N(\ram[166][10] ), .A1N(n6444), 
        .Y(n3248) );
  OAI2BB2XL U3225 ( .B0(n6708), .B1(n552), .A0N(\ram[166][11] ), .A1N(n6444), 
        .Y(n3249) );
  OAI2BB2XL U3226 ( .B0(n6685), .B1(n552), .A0N(\ram[166][12] ), .A1N(n6444), 
        .Y(n3250) );
  OAI2BB2XL U3227 ( .B0(n6662), .B1(n552), .A0N(\ram[166][13] ), .A1N(n6444), 
        .Y(n3251) );
  OAI2BB2XL U3228 ( .B0(n6639), .B1(n552), .A0N(\ram[166][14] ), .A1N(n6444), 
        .Y(n3252) );
  OAI2BB2XL U3229 ( .B0(n6616), .B1(n552), .A0N(\ram[166][15] ), .A1N(n6444), 
        .Y(n3253) );
  OAI2BB2XL U3230 ( .B0(n6966), .B1(n555), .A0N(\ram[167][0] ), .A1N(n6443), 
        .Y(n3254) );
  OAI2BB2XL U3231 ( .B0(n6943), .B1(n555), .A0N(\ram[167][1] ), .A1N(n6443), 
        .Y(n3255) );
  OAI2BB2XL U3232 ( .B0(n6920), .B1(n555), .A0N(\ram[167][2] ), .A1N(n6443), 
        .Y(n3256) );
  OAI2BB2XL U3233 ( .B0(n6897), .B1(n555), .A0N(\ram[167][3] ), .A1N(n6443), 
        .Y(n3257) );
  OAI2BB2XL U3234 ( .B0(n6869), .B1(n555), .A0N(\ram[167][4] ), .A1N(n6443), 
        .Y(n3258) );
  OAI2BB2XL U3235 ( .B0(n6846), .B1(n555), .A0N(\ram[167][5] ), .A1N(n6443), 
        .Y(n3259) );
  OAI2BB2XL U3236 ( .B0(n6823), .B1(n555), .A0N(\ram[167][6] ), .A1N(n6443), 
        .Y(n3260) );
  OAI2BB2XL U3237 ( .B0(n6800), .B1(n555), .A0N(\ram[167][7] ), .A1N(n6443), 
        .Y(n3261) );
  OAI2BB2XL U3238 ( .B0(n6777), .B1(n555), .A0N(\ram[167][8] ), .A1N(n6443), 
        .Y(n3262) );
  OAI2BB2XL U3239 ( .B0(n6754), .B1(n555), .A0N(\ram[167][9] ), .A1N(n6443), 
        .Y(n3263) );
  OAI2BB2XL U3240 ( .B0(n6731), .B1(n555), .A0N(\ram[167][10] ), .A1N(n6443), 
        .Y(n3264) );
  OAI2BB2XL U3241 ( .B0(n6708), .B1(n555), .A0N(\ram[167][11] ), .A1N(n6443), 
        .Y(n3265) );
  OAI2BB2XL U3242 ( .B0(n6685), .B1(n555), .A0N(\ram[167][12] ), .A1N(n6443), 
        .Y(n3266) );
  OAI2BB2XL U3243 ( .B0(n6662), .B1(n555), .A0N(\ram[167][13] ), .A1N(n6443), 
        .Y(n3267) );
  OAI2BB2XL U3244 ( .B0(n6639), .B1(n555), .A0N(\ram[167][14] ), .A1N(n6443), 
        .Y(n3268) );
  OAI2BB2XL U3245 ( .B0(n6616), .B1(n555), .A0N(\ram[167][15] ), .A1N(n6443), 
        .Y(n3269) );
  OAI2BB2XL U3246 ( .B0(n6966), .B1(n321), .A0N(\ram[168][0] ), .A1N(n6442), 
        .Y(n3270) );
  OAI2BB2XL U3247 ( .B0(n6943), .B1(n321), .A0N(\ram[168][1] ), .A1N(n6442), 
        .Y(n3271) );
  OAI2BB2XL U3248 ( .B0(n6920), .B1(n321), .A0N(\ram[168][2] ), .A1N(n6442), 
        .Y(n3272) );
  OAI2BB2XL U3249 ( .B0(n6897), .B1(n321), .A0N(\ram[168][3] ), .A1N(n6442), 
        .Y(n3273) );
  OAI2BB2XL U3250 ( .B0(n6869), .B1(n321), .A0N(\ram[168][4] ), .A1N(n6442), 
        .Y(n3274) );
  OAI2BB2XL U3251 ( .B0(n6846), .B1(n321), .A0N(\ram[168][5] ), .A1N(n6442), 
        .Y(n3275) );
  OAI2BB2XL U3252 ( .B0(n6823), .B1(n321), .A0N(\ram[168][6] ), .A1N(n6442), 
        .Y(n3276) );
  OAI2BB2XL U3253 ( .B0(n6800), .B1(n321), .A0N(\ram[168][7] ), .A1N(n6442), 
        .Y(n3277) );
  OAI2BB2XL U3254 ( .B0(n6777), .B1(n321), .A0N(\ram[168][8] ), .A1N(n6442), 
        .Y(n3278) );
  OAI2BB2XL U3255 ( .B0(n6754), .B1(n321), .A0N(\ram[168][9] ), .A1N(n6442), 
        .Y(n3279) );
  OAI2BB2XL U3256 ( .B0(n6731), .B1(n321), .A0N(\ram[168][10] ), .A1N(n6442), 
        .Y(n3280) );
  OAI2BB2XL U3257 ( .B0(n6708), .B1(n321), .A0N(\ram[168][11] ), .A1N(n6442), 
        .Y(n3281) );
  OAI2BB2XL U3258 ( .B0(n6685), .B1(n321), .A0N(\ram[168][12] ), .A1N(n6442), 
        .Y(n3282) );
  OAI2BB2XL U3259 ( .B0(n6662), .B1(n321), .A0N(\ram[168][13] ), .A1N(n6442), 
        .Y(n3283) );
  OAI2BB2XL U3260 ( .B0(n6639), .B1(n321), .A0N(\ram[168][14] ), .A1N(n6442), 
        .Y(n3284) );
  OAI2BB2XL U3261 ( .B0(n6616), .B1(n321), .A0N(\ram[168][15] ), .A1N(n6442), 
        .Y(n3285) );
  OAI2BB2XL U3262 ( .B0(n6966), .B1(n323), .A0N(\ram[169][0] ), .A1N(n6441), 
        .Y(n3286) );
  OAI2BB2XL U3263 ( .B0(n6943), .B1(n323), .A0N(\ram[169][1] ), .A1N(n6441), 
        .Y(n3287) );
  OAI2BB2XL U3264 ( .B0(n6920), .B1(n323), .A0N(\ram[169][2] ), .A1N(n6441), 
        .Y(n3288) );
  OAI2BB2XL U3265 ( .B0(n6897), .B1(n323), .A0N(\ram[169][3] ), .A1N(n6441), 
        .Y(n3289) );
  OAI2BB2XL U3266 ( .B0(n6869), .B1(n323), .A0N(\ram[169][4] ), .A1N(n6441), 
        .Y(n3290) );
  OAI2BB2XL U3267 ( .B0(n6846), .B1(n323), .A0N(\ram[169][5] ), .A1N(n6441), 
        .Y(n3291) );
  OAI2BB2XL U3268 ( .B0(n6823), .B1(n323), .A0N(\ram[169][6] ), .A1N(n6441), 
        .Y(n3292) );
  OAI2BB2XL U3269 ( .B0(n6800), .B1(n323), .A0N(\ram[169][7] ), .A1N(n6441), 
        .Y(n3293) );
  OAI2BB2XL U3270 ( .B0(n6777), .B1(n323), .A0N(\ram[169][8] ), .A1N(n6441), 
        .Y(n3294) );
  OAI2BB2XL U3271 ( .B0(n6754), .B1(n323), .A0N(\ram[169][9] ), .A1N(n6441), 
        .Y(n3295) );
  OAI2BB2XL U3272 ( .B0(n6731), .B1(n323), .A0N(\ram[169][10] ), .A1N(n6441), 
        .Y(n3296) );
  OAI2BB2XL U3273 ( .B0(n6708), .B1(n323), .A0N(\ram[169][11] ), .A1N(n6441), 
        .Y(n3297) );
  OAI2BB2XL U3274 ( .B0(n6685), .B1(n323), .A0N(\ram[169][12] ), .A1N(n6441), 
        .Y(n3298) );
  OAI2BB2XL U3275 ( .B0(n6662), .B1(n323), .A0N(\ram[169][13] ), .A1N(n6441), 
        .Y(n3299) );
  OAI2BB2XL U3276 ( .B0(n6639), .B1(n323), .A0N(\ram[169][14] ), .A1N(n6441), 
        .Y(n3300) );
  OAI2BB2XL U3277 ( .B0(n6616), .B1(n323), .A0N(\ram[169][15] ), .A1N(n6441), 
        .Y(n3301) );
  OAI2BB2XL U3278 ( .B0(n6966), .B1(n464), .A0N(\ram[170][0] ), .A1N(n6440), 
        .Y(n3302) );
  OAI2BB2XL U3279 ( .B0(n6943), .B1(n464), .A0N(\ram[170][1] ), .A1N(n6440), 
        .Y(n3303) );
  OAI2BB2XL U3280 ( .B0(n6920), .B1(n464), .A0N(\ram[170][2] ), .A1N(n6440), 
        .Y(n3304) );
  OAI2BB2XL U3281 ( .B0(n6897), .B1(n464), .A0N(\ram[170][3] ), .A1N(n6440), 
        .Y(n3305) );
  OAI2BB2XL U3282 ( .B0(n6869), .B1(n464), .A0N(\ram[170][4] ), .A1N(n6440), 
        .Y(n3306) );
  OAI2BB2XL U3283 ( .B0(n6846), .B1(n464), .A0N(\ram[170][5] ), .A1N(n6440), 
        .Y(n3307) );
  OAI2BB2XL U3284 ( .B0(n6823), .B1(n464), .A0N(\ram[170][6] ), .A1N(n6440), 
        .Y(n3308) );
  OAI2BB2XL U3285 ( .B0(n6800), .B1(n464), .A0N(\ram[170][7] ), .A1N(n6440), 
        .Y(n3309) );
  OAI2BB2XL U3286 ( .B0(n6777), .B1(n464), .A0N(\ram[170][8] ), .A1N(n6440), 
        .Y(n3310) );
  OAI2BB2XL U3287 ( .B0(n6754), .B1(n464), .A0N(\ram[170][9] ), .A1N(n6440), 
        .Y(n3311) );
  OAI2BB2XL U3288 ( .B0(n6731), .B1(n464), .A0N(\ram[170][10] ), .A1N(n6440), 
        .Y(n3312) );
  OAI2BB2XL U3289 ( .B0(n6708), .B1(n464), .A0N(\ram[170][11] ), .A1N(n6440), 
        .Y(n3313) );
  OAI2BB2XL U3290 ( .B0(n6685), .B1(n464), .A0N(\ram[170][12] ), .A1N(n6440), 
        .Y(n3314) );
  OAI2BB2XL U3291 ( .B0(n6662), .B1(n464), .A0N(\ram[170][13] ), .A1N(n6440), 
        .Y(n3315) );
  OAI2BB2XL U3292 ( .B0(n6639), .B1(n464), .A0N(\ram[170][14] ), .A1N(n6440), 
        .Y(n3316) );
  OAI2BB2XL U3293 ( .B0(n6616), .B1(n464), .A0N(\ram[170][15] ), .A1N(n6440), 
        .Y(n3317) );
  OAI2BB2XL U3294 ( .B0(n6966), .B1(n325), .A0N(\ram[171][0] ), .A1N(n6439), 
        .Y(n3318) );
  OAI2BB2XL U3295 ( .B0(n6943), .B1(n325), .A0N(\ram[171][1] ), .A1N(n6439), 
        .Y(n3319) );
  OAI2BB2XL U3296 ( .B0(n6920), .B1(n325), .A0N(\ram[171][2] ), .A1N(n6439), 
        .Y(n3320) );
  OAI2BB2XL U3297 ( .B0(n6897), .B1(n325), .A0N(\ram[171][3] ), .A1N(n6439), 
        .Y(n3321) );
  OAI2BB2XL U3298 ( .B0(n6869), .B1(n325), .A0N(\ram[171][4] ), .A1N(n6439), 
        .Y(n3322) );
  OAI2BB2XL U3299 ( .B0(n6846), .B1(n325), .A0N(\ram[171][5] ), .A1N(n6439), 
        .Y(n3323) );
  OAI2BB2XL U3300 ( .B0(n6823), .B1(n325), .A0N(\ram[171][6] ), .A1N(n6439), 
        .Y(n3324) );
  OAI2BB2XL U3301 ( .B0(n6800), .B1(n325), .A0N(\ram[171][7] ), .A1N(n6439), 
        .Y(n3325) );
  OAI2BB2XL U3302 ( .B0(n6777), .B1(n325), .A0N(\ram[171][8] ), .A1N(n6439), 
        .Y(n3326) );
  OAI2BB2XL U3303 ( .B0(n6754), .B1(n325), .A0N(\ram[171][9] ), .A1N(n6439), 
        .Y(n3327) );
  OAI2BB2XL U3304 ( .B0(n6731), .B1(n325), .A0N(\ram[171][10] ), .A1N(n6439), 
        .Y(n3328) );
  OAI2BB2XL U3305 ( .B0(n6708), .B1(n325), .A0N(\ram[171][11] ), .A1N(n6439), 
        .Y(n3329) );
  OAI2BB2XL U3306 ( .B0(n6685), .B1(n325), .A0N(\ram[171][12] ), .A1N(n6439), 
        .Y(n3330) );
  OAI2BB2XL U3307 ( .B0(n6662), .B1(n325), .A0N(\ram[171][13] ), .A1N(n6439), 
        .Y(n3331) );
  OAI2BB2XL U3308 ( .B0(n6639), .B1(n325), .A0N(\ram[171][14] ), .A1N(n6439), 
        .Y(n3332) );
  OAI2BB2XL U3309 ( .B0(n6616), .B1(n325), .A0N(\ram[171][15] ), .A1N(n6439), 
        .Y(n3333) );
  OAI2BB2XL U3310 ( .B0(n6965), .B1(n327), .A0N(\ram[172][0] ), .A1N(n6438), 
        .Y(n3334) );
  OAI2BB2XL U3311 ( .B0(n6942), .B1(n327), .A0N(\ram[172][1] ), .A1N(n6438), 
        .Y(n3335) );
  OAI2BB2XL U3312 ( .B0(n6919), .B1(n327), .A0N(\ram[172][2] ), .A1N(n6438), 
        .Y(n3336) );
  OAI2BB2XL U3313 ( .B0(n6896), .B1(n327), .A0N(\ram[172][3] ), .A1N(n6438), 
        .Y(n3337) );
  OAI2BB2XL U3314 ( .B0(n6868), .B1(n327), .A0N(\ram[172][4] ), .A1N(n6438), 
        .Y(n3338) );
  OAI2BB2XL U3315 ( .B0(n6845), .B1(n327), .A0N(\ram[172][5] ), .A1N(n6438), 
        .Y(n3339) );
  OAI2BB2XL U3316 ( .B0(n6822), .B1(n327), .A0N(\ram[172][6] ), .A1N(n6438), 
        .Y(n3340) );
  OAI2BB2XL U3317 ( .B0(n6799), .B1(n327), .A0N(\ram[172][7] ), .A1N(n6438), 
        .Y(n3341) );
  OAI2BB2XL U3318 ( .B0(n6776), .B1(n327), .A0N(\ram[172][8] ), .A1N(n6438), 
        .Y(n3342) );
  OAI2BB2XL U3319 ( .B0(n6753), .B1(n327), .A0N(\ram[172][9] ), .A1N(n6438), 
        .Y(n3343) );
  OAI2BB2XL U3320 ( .B0(n6730), .B1(n327), .A0N(\ram[172][10] ), .A1N(n6438), 
        .Y(n3344) );
  OAI2BB2XL U3321 ( .B0(n6707), .B1(n327), .A0N(\ram[172][11] ), .A1N(n6438), 
        .Y(n3345) );
  OAI2BB2XL U3322 ( .B0(n6684), .B1(n327), .A0N(\ram[172][12] ), .A1N(n6438), 
        .Y(n3346) );
  OAI2BB2XL U3323 ( .B0(n6661), .B1(n327), .A0N(\ram[172][13] ), .A1N(n6438), 
        .Y(n3347) );
  OAI2BB2XL U3324 ( .B0(n6638), .B1(n327), .A0N(\ram[172][14] ), .A1N(n6438), 
        .Y(n3348) );
  OAI2BB2XL U3325 ( .B0(n6615), .B1(n327), .A0N(\ram[172][15] ), .A1N(n6438), 
        .Y(n3349) );
  OAI2BB2XL U3326 ( .B0(n6965), .B1(n329), .A0N(\ram[173][0] ), .A1N(n6437), 
        .Y(n3350) );
  OAI2BB2XL U3327 ( .B0(n6942), .B1(n329), .A0N(\ram[173][1] ), .A1N(n6437), 
        .Y(n3351) );
  OAI2BB2XL U3328 ( .B0(n6919), .B1(n329), .A0N(\ram[173][2] ), .A1N(n6437), 
        .Y(n3352) );
  OAI2BB2XL U3329 ( .B0(n6896), .B1(n329), .A0N(\ram[173][3] ), .A1N(n6437), 
        .Y(n3353) );
  OAI2BB2XL U3330 ( .B0(n6867), .B1(n329), .A0N(\ram[173][4] ), .A1N(n6437), 
        .Y(n3354) );
  OAI2BB2XL U3331 ( .B0(n6844), .B1(n329), .A0N(\ram[173][5] ), .A1N(n6437), 
        .Y(n3355) );
  OAI2BB2XL U3332 ( .B0(n6821), .B1(n329), .A0N(\ram[173][6] ), .A1N(n6437), 
        .Y(n3356) );
  OAI2BB2XL U3333 ( .B0(n6798), .B1(n329), .A0N(\ram[173][7] ), .A1N(n6437), 
        .Y(n3357) );
  OAI2BB2XL U3334 ( .B0(n6775), .B1(n329), .A0N(\ram[173][8] ), .A1N(n6437), 
        .Y(n3358) );
  OAI2BB2XL U3335 ( .B0(n6752), .B1(n329), .A0N(\ram[173][9] ), .A1N(n6437), 
        .Y(n3359) );
  OAI2BB2XL U3336 ( .B0(n6729), .B1(n329), .A0N(\ram[173][10] ), .A1N(n6437), 
        .Y(n3360) );
  OAI2BB2XL U3337 ( .B0(n6706), .B1(n329), .A0N(\ram[173][11] ), .A1N(n6437), 
        .Y(n3361) );
  OAI2BB2XL U3338 ( .B0(n6683), .B1(n329), .A0N(\ram[173][12] ), .A1N(n6437), 
        .Y(n3362) );
  OAI2BB2XL U3339 ( .B0(n6660), .B1(n329), .A0N(\ram[173][13] ), .A1N(n6437), 
        .Y(n3363) );
  OAI2BB2XL U3340 ( .B0(n6637), .B1(n329), .A0N(\ram[173][14] ), .A1N(n6437), 
        .Y(n3364) );
  OAI2BB2XL U3341 ( .B0(n6614), .B1(n329), .A0N(\ram[173][15] ), .A1N(n6437), 
        .Y(n3365) );
  OAI2BB2XL U3342 ( .B0(n6965), .B1(n331), .A0N(\ram[174][0] ), .A1N(n6436), 
        .Y(n3366) );
  OAI2BB2XL U3343 ( .B0(n6942), .B1(n331), .A0N(\ram[174][1] ), .A1N(n6436), 
        .Y(n3367) );
  OAI2BB2XL U3344 ( .B0(n6919), .B1(n331), .A0N(\ram[174][2] ), .A1N(n6436), 
        .Y(n3368) );
  OAI2BB2XL U3345 ( .B0(n6896), .B1(n331), .A0N(\ram[174][3] ), .A1N(n6436), 
        .Y(n3369) );
  OAI2BB2XL U3346 ( .B0(n6869), .B1(n331), .A0N(\ram[174][4] ), .A1N(n6436), 
        .Y(n3370) );
  OAI2BB2XL U3347 ( .B0(n6846), .B1(n331), .A0N(\ram[174][5] ), .A1N(n6436), 
        .Y(n3371) );
  OAI2BB2XL U3348 ( .B0(n6823), .B1(n331), .A0N(\ram[174][6] ), .A1N(n6436), 
        .Y(n3372) );
  OAI2BB2XL U3349 ( .B0(n6800), .B1(n331), .A0N(\ram[174][7] ), .A1N(n6436), 
        .Y(n3373) );
  OAI2BB2XL U3350 ( .B0(n6777), .B1(n331), .A0N(\ram[174][8] ), .A1N(n6436), 
        .Y(n3374) );
  OAI2BB2XL U3351 ( .B0(n6754), .B1(n331), .A0N(\ram[174][9] ), .A1N(n6436), 
        .Y(n3375) );
  OAI2BB2XL U3352 ( .B0(n6731), .B1(n331), .A0N(\ram[174][10] ), .A1N(n6436), 
        .Y(n3376) );
  OAI2BB2XL U3353 ( .B0(n6708), .B1(n331), .A0N(\ram[174][11] ), .A1N(n6436), 
        .Y(n3377) );
  OAI2BB2XL U3354 ( .B0(n6685), .B1(n331), .A0N(\ram[174][12] ), .A1N(n6436), 
        .Y(n3378) );
  OAI2BB2XL U3355 ( .B0(n6662), .B1(n331), .A0N(\ram[174][13] ), .A1N(n6436), 
        .Y(n3379) );
  OAI2BB2XL U3356 ( .B0(n6639), .B1(n331), .A0N(\ram[174][14] ), .A1N(n6436), 
        .Y(n3380) );
  OAI2BB2XL U3357 ( .B0(n6616), .B1(n331), .A0N(\ram[174][15] ), .A1N(n6436), 
        .Y(n3381) );
  OAI2BB2XL U3358 ( .B0(n6965), .B1(n333), .A0N(\ram[175][0] ), .A1N(n6435), 
        .Y(n3382) );
  OAI2BB2XL U3359 ( .B0(n6942), .B1(n333), .A0N(\ram[175][1] ), .A1N(n6435), 
        .Y(n3383) );
  OAI2BB2XL U3360 ( .B0(n6919), .B1(n333), .A0N(\ram[175][2] ), .A1N(n6435), 
        .Y(n3384) );
  OAI2BB2XL U3361 ( .B0(n6896), .B1(n333), .A0N(\ram[175][3] ), .A1N(n6435), 
        .Y(n3385) );
  OAI2BB2XL U3362 ( .B0(n6868), .B1(n333), .A0N(\ram[175][4] ), .A1N(n6435), 
        .Y(n3386) );
  OAI2BB2XL U3363 ( .B0(n6845), .B1(n333), .A0N(\ram[175][5] ), .A1N(n6435), 
        .Y(n3387) );
  OAI2BB2XL U3364 ( .B0(n6822), .B1(n333), .A0N(\ram[175][6] ), .A1N(n6435), 
        .Y(n3388) );
  OAI2BB2XL U3365 ( .B0(n6799), .B1(n333), .A0N(\ram[175][7] ), .A1N(n6435), 
        .Y(n3389) );
  OAI2BB2XL U3366 ( .B0(n6776), .B1(n333), .A0N(\ram[175][8] ), .A1N(n6435), 
        .Y(n3390) );
  OAI2BB2XL U3367 ( .B0(n6753), .B1(n333), .A0N(\ram[175][9] ), .A1N(n6435), 
        .Y(n3391) );
  OAI2BB2XL U3368 ( .B0(n6730), .B1(n333), .A0N(\ram[175][10] ), .A1N(n6435), 
        .Y(n3392) );
  OAI2BB2XL U3369 ( .B0(n6707), .B1(n333), .A0N(\ram[175][11] ), .A1N(n6435), 
        .Y(n3393) );
  OAI2BB2XL U3370 ( .B0(n6684), .B1(n333), .A0N(\ram[175][12] ), .A1N(n6435), 
        .Y(n3394) );
  OAI2BB2XL U3371 ( .B0(n6661), .B1(n333), .A0N(\ram[175][13] ), .A1N(n6435), 
        .Y(n3395) );
  OAI2BB2XL U3372 ( .B0(n6638), .B1(n333), .A0N(\ram[175][14] ), .A1N(n6435), 
        .Y(n3396) );
  OAI2BB2XL U3373 ( .B0(n6615), .B1(n333), .A0N(\ram[175][15] ), .A1N(n6435), 
        .Y(n3397) );
  OAI2BB2XL U3374 ( .B0(n6965), .B1(n335), .A0N(\ram[176][0] ), .A1N(n6434), 
        .Y(n3398) );
  OAI2BB2XL U3375 ( .B0(n6942), .B1(n335), .A0N(\ram[176][1] ), .A1N(n6434), 
        .Y(n3399) );
  OAI2BB2XL U3376 ( .B0(n6919), .B1(n335), .A0N(\ram[176][2] ), .A1N(n6434), 
        .Y(n3400) );
  OAI2BB2XL U3377 ( .B0(n6896), .B1(n335), .A0N(\ram[176][3] ), .A1N(n6434), 
        .Y(n3401) );
  OAI2BB2XL U3378 ( .B0(n6867), .B1(n335), .A0N(\ram[176][4] ), .A1N(n6434), 
        .Y(n3402) );
  OAI2BB2XL U3379 ( .B0(n6844), .B1(n335), .A0N(\ram[176][5] ), .A1N(n6434), 
        .Y(n3403) );
  OAI2BB2XL U3380 ( .B0(n6821), .B1(n335), .A0N(\ram[176][6] ), .A1N(n6434), 
        .Y(n3404) );
  OAI2BB2XL U3381 ( .B0(n6798), .B1(n335), .A0N(\ram[176][7] ), .A1N(n6434), 
        .Y(n3405) );
  OAI2BB2XL U3382 ( .B0(n6775), .B1(n335), .A0N(\ram[176][8] ), .A1N(n6434), 
        .Y(n3406) );
  OAI2BB2XL U3383 ( .B0(n6752), .B1(n335), .A0N(\ram[176][9] ), .A1N(n6434), 
        .Y(n3407) );
  OAI2BB2XL U3384 ( .B0(n6729), .B1(n335), .A0N(\ram[176][10] ), .A1N(n6434), 
        .Y(n3408) );
  OAI2BB2XL U3385 ( .B0(n6706), .B1(n335), .A0N(\ram[176][11] ), .A1N(n6434), 
        .Y(n3409) );
  OAI2BB2XL U3386 ( .B0(n6683), .B1(n335), .A0N(\ram[176][12] ), .A1N(n6434), 
        .Y(n3410) );
  OAI2BB2XL U3387 ( .B0(n6660), .B1(n335), .A0N(\ram[176][13] ), .A1N(n6434), 
        .Y(n3411) );
  OAI2BB2XL U3388 ( .B0(n6637), .B1(n335), .A0N(\ram[176][14] ), .A1N(n6434), 
        .Y(n3412) );
  OAI2BB2XL U3389 ( .B0(n6614), .B1(n335), .A0N(\ram[176][15] ), .A1N(n6434), 
        .Y(n3413) );
  OAI2BB2XL U3390 ( .B0(n6965), .B1(n337), .A0N(\ram[177][0] ), .A1N(n6433), 
        .Y(n3414) );
  OAI2BB2XL U3391 ( .B0(n6942), .B1(n337), .A0N(\ram[177][1] ), .A1N(n6433), 
        .Y(n3415) );
  OAI2BB2XL U3392 ( .B0(n6919), .B1(n337), .A0N(\ram[177][2] ), .A1N(n6433), 
        .Y(n3416) );
  OAI2BB2XL U3393 ( .B0(n6896), .B1(n337), .A0N(\ram[177][3] ), .A1N(n6433), 
        .Y(n3417) );
  OAI2BB2XL U3394 ( .B0(n6869), .B1(n337), .A0N(\ram[177][4] ), .A1N(n6433), 
        .Y(n3418) );
  OAI2BB2XL U3395 ( .B0(n6846), .B1(n337), .A0N(\ram[177][5] ), .A1N(n6433), 
        .Y(n3419) );
  OAI2BB2XL U3396 ( .B0(n6823), .B1(n337), .A0N(\ram[177][6] ), .A1N(n6433), 
        .Y(n3420) );
  OAI2BB2XL U3397 ( .B0(n6800), .B1(n337), .A0N(\ram[177][7] ), .A1N(n6433), 
        .Y(n3421) );
  OAI2BB2XL U3398 ( .B0(n6777), .B1(n337), .A0N(\ram[177][8] ), .A1N(n6433), 
        .Y(n3422) );
  OAI2BB2XL U3399 ( .B0(n6754), .B1(n337), .A0N(\ram[177][9] ), .A1N(n6433), 
        .Y(n3423) );
  OAI2BB2XL U3400 ( .B0(n6731), .B1(n337), .A0N(\ram[177][10] ), .A1N(n6433), 
        .Y(n3424) );
  OAI2BB2XL U3401 ( .B0(n6708), .B1(n337), .A0N(\ram[177][11] ), .A1N(n6433), 
        .Y(n3425) );
  OAI2BB2XL U3402 ( .B0(n6685), .B1(n337), .A0N(\ram[177][12] ), .A1N(n6433), 
        .Y(n3426) );
  OAI2BB2XL U3403 ( .B0(n6662), .B1(n337), .A0N(\ram[177][13] ), .A1N(n6433), 
        .Y(n3427) );
  OAI2BB2XL U3404 ( .B0(n6639), .B1(n337), .A0N(\ram[177][14] ), .A1N(n6433), 
        .Y(n3428) );
  OAI2BB2XL U3405 ( .B0(n6616), .B1(n337), .A0N(\ram[177][15] ), .A1N(n6433), 
        .Y(n3429) );
  OAI2BB2XL U3406 ( .B0(n6965), .B1(n339), .A0N(\ram[178][0] ), .A1N(n6432), 
        .Y(n3430) );
  OAI2BB2XL U3407 ( .B0(n6942), .B1(n339), .A0N(\ram[178][1] ), .A1N(n6432), 
        .Y(n3431) );
  OAI2BB2XL U3408 ( .B0(n6919), .B1(n339), .A0N(\ram[178][2] ), .A1N(n6432), 
        .Y(n3432) );
  OAI2BB2XL U3409 ( .B0(n6896), .B1(n339), .A0N(\ram[178][3] ), .A1N(n6432), 
        .Y(n3433) );
  OAI2BB2XL U3410 ( .B0(n6868), .B1(n339), .A0N(\ram[178][4] ), .A1N(n6432), 
        .Y(n3434) );
  OAI2BB2XL U3411 ( .B0(n6845), .B1(n339), .A0N(\ram[178][5] ), .A1N(n6432), 
        .Y(n3435) );
  OAI2BB2XL U3412 ( .B0(n6822), .B1(n339), .A0N(\ram[178][6] ), .A1N(n6432), 
        .Y(n3436) );
  OAI2BB2XL U3413 ( .B0(n6799), .B1(n339), .A0N(\ram[178][7] ), .A1N(n6432), 
        .Y(n3437) );
  OAI2BB2XL U3414 ( .B0(n6776), .B1(n339), .A0N(\ram[178][8] ), .A1N(n6432), 
        .Y(n3438) );
  OAI2BB2XL U3415 ( .B0(n6753), .B1(n339), .A0N(\ram[178][9] ), .A1N(n6432), 
        .Y(n3439) );
  OAI2BB2XL U3416 ( .B0(n6730), .B1(n339), .A0N(\ram[178][10] ), .A1N(n6432), 
        .Y(n3440) );
  OAI2BB2XL U3417 ( .B0(n6707), .B1(n339), .A0N(\ram[178][11] ), .A1N(n6432), 
        .Y(n3441) );
  OAI2BB2XL U3418 ( .B0(n6684), .B1(n339), .A0N(\ram[178][12] ), .A1N(n6432), 
        .Y(n3442) );
  OAI2BB2XL U3419 ( .B0(n6661), .B1(n339), .A0N(\ram[178][13] ), .A1N(n6432), 
        .Y(n3443) );
  OAI2BB2XL U3420 ( .B0(n6638), .B1(n339), .A0N(\ram[178][14] ), .A1N(n6432), 
        .Y(n3444) );
  OAI2BB2XL U3421 ( .B0(n6615), .B1(n339), .A0N(\ram[178][15] ), .A1N(n6432), 
        .Y(n3445) );
  OAI2BB2XL U3422 ( .B0(n6965), .B1(n342), .A0N(\ram[179][0] ), .A1N(n6431), 
        .Y(n3446) );
  OAI2BB2XL U3423 ( .B0(n6942), .B1(n342), .A0N(\ram[179][1] ), .A1N(n6431), 
        .Y(n3447) );
  OAI2BB2XL U3424 ( .B0(n6919), .B1(n342), .A0N(\ram[179][2] ), .A1N(n6431), 
        .Y(n3448) );
  OAI2BB2XL U3425 ( .B0(n6896), .B1(n342), .A0N(\ram[179][3] ), .A1N(n6431), 
        .Y(n3449) );
  OAI2BB2XL U3426 ( .B0(n6867), .B1(n342), .A0N(\ram[179][4] ), .A1N(n6431), 
        .Y(n3450) );
  OAI2BB2XL U3427 ( .B0(n6844), .B1(n342), .A0N(\ram[179][5] ), .A1N(n6431), 
        .Y(n3451) );
  OAI2BB2XL U3428 ( .B0(n6821), .B1(n342), .A0N(\ram[179][6] ), .A1N(n6431), 
        .Y(n3452) );
  OAI2BB2XL U3429 ( .B0(n6798), .B1(n342), .A0N(\ram[179][7] ), .A1N(n6431), 
        .Y(n3453) );
  OAI2BB2XL U3430 ( .B0(n6775), .B1(n342), .A0N(\ram[179][8] ), .A1N(n6431), 
        .Y(n3454) );
  OAI2BB2XL U3431 ( .B0(n6752), .B1(n342), .A0N(\ram[179][9] ), .A1N(n6431), 
        .Y(n3455) );
  OAI2BB2XL U3432 ( .B0(n6729), .B1(n342), .A0N(\ram[179][10] ), .A1N(n6431), 
        .Y(n3456) );
  OAI2BB2XL U3433 ( .B0(n6706), .B1(n342), .A0N(\ram[179][11] ), .A1N(n6431), 
        .Y(n3457) );
  OAI2BB2XL U3434 ( .B0(n6683), .B1(n342), .A0N(\ram[179][12] ), .A1N(n6431), 
        .Y(n3458) );
  OAI2BB2XL U3435 ( .B0(n6660), .B1(n342), .A0N(\ram[179][13] ), .A1N(n6431), 
        .Y(n3459) );
  OAI2BB2XL U3436 ( .B0(n6637), .B1(n342), .A0N(\ram[179][14] ), .A1N(n6431), 
        .Y(n3460) );
  OAI2BB2XL U3437 ( .B0(n6614), .B1(n342), .A0N(\ram[179][15] ), .A1N(n6431), 
        .Y(n3461) );
  OAI2BB2XL U3438 ( .B0(n6965), .B1(n344), .A0N(\ram[180][0] ), .A1N(n6430), 
        .Y(n3462) );
  OAI2BB2XL U3439 ( .B0(n6942), .B1(n344), .A0N(\ram[180][1] ), .A1N(n6430), 
        .Y(n3463) );
  OAI2BB2XL U3440 ( .B0(n6919), .B1(n344), .A0N(\ram[180][2] ), .A1N(n6430), 
        .Y(n3464) );
  OAI2BB2XL U3441 ( .B0(n6896), .B1(n344), .A0N(\ram[180][3] ), .A1N(n6430), 
        .Y(n3465) );
  OAI2BB2XL U3442 ( .B0(n6869), .B1(n344), .A0N(\ram[180][4] ), .A1N(n6430), 
        .Y(n3466) );
  OAI2BB2XL U3443 ( .B0(n6846), .B1(n344), .A0N(\ram[180][5] ), .A1N(n6430), 
        .Y(n3467) );
  OAI2BB2XL U3444 ( .B0(n6823), .B1(n344), .A0N(\ram[180][6] ), .A1N(n6430), 
        .Y(n3468) );
  OAI2BB2XL U3445 ( .B0(n6800), .B1(n344), .A0N(\ram[180][7] ), .A1N(n6430), 
        .Y(n3469) );
  OAI2BB2XL U3446 ( .B0(n6777), .B1(n344), .A0N(\ram[180][8] ), .A1N(n6430), 
        .Y(n3470) );
  OAI2BB2XL U3447 ( .B0(n6754), .B1(n344), .A0N(\ram[180][9] ), .A1N(n6430), 
        .Y(n3471) );
  OAI2BB2XL U3448 ( .B0(n6731), .B1(n344), .A0N(\ram[180][10] ), .A1N(n6430), 
        .Y(n3472) );
  OAI2BB2XL U3449 ( .B0(n6708), .B1(n344), .A0N(\ram[180][11] ), .A1N(n6430), 
        .Y(n3473) );
  OAI2BB2XL U3450 ( .B0(n6685), .B1(n344), .A0N(\ram[180][12] ), .A1N(n6430), 
        .Y(n3474) );
  OAI2BB2XL U3451 ( .B0(n6662), .B1(n344), .A0N(\ram[180][13] ), .A1N(n6430), 
        .Y(n3475) );
  OAI2BB2XL U3452 ( .B0(n6639), .B1(n344), .A0N(\ram[180][14] ), .A1N(n6430), 
        .Y(n3476) );
  OAI2BB2XL U3453 ( .B0(n6616), .B1(n344), .A0N(\ram[180][15] ), .A1N(n6430), 
        .Y(n3477) );
  OAI2BB2XL U3454 ( .B0(n6965), .B1(n511), .A0N(\ram[181][0] ), .A1N(n6429), 
        .Y(n3478) );
  OAI2BB2XL U3455 ( .B0(n6942), .B1(n511), .A0N(\ram[181][1] ), .A1N(n6429), 
        .Y(n3479) );
  OAI2BB2XL U3456 ( .B0(n6919), .B1(n511), .A0N(\ram[181][2] ), .A1N(n6429), 
        .Y(n3480) );
  OAI2BB2XL U3457 ( .B0(n6896), .B1(n511), .A0N(\ram[181][3] ), .A1N(n6429), 
        .Y(n3481) );
  OAI2BB2XL U3458 ( .B0(n6865), .B1(n511), .A0N(\ram[181][4] ), .A1N(n6429), 
        .Y(n3482) );
  OAI2BB2XL U3459 ( .B0(n6842), .B1(n511), .A0N(\ram[181][5] ), .A1N(n6429), 
        .Y(n3483) );
  OAI2BB2XL U3460 ( .B0(n6819), .B1(n511), .A0N(\ram[181][6] ), .A1N(n6429), 
        .Y(n3484) );
  OAI2BB2XL U3461 ( .B0(n6796), .B1(n511), .A0N(\ram[181][7] ), .A1N(n6429), 
        .Y(n3485) );
  OAI2BB2XL U3462 ( .B0(n6773), .B1(n511), .A0N(\ram[181][8] ), .A1N(n6429), 
        .Y(n3486) );
  OAI2BB2XL U3463 ( .B0(n6750), .B1(n511), .A0N(\ram[181][9] ), .A1N(n6429), 
        .Y(n3487) );
  OAI2BB2XL U3464 ( .B0(n6727), .B1(n511), .A0N(\ram[181][10] ), .A1N(n6429), 
        .Y(n3488) );
  OAI2BB2XL U3465 ( .B0(n6704), .B1(n511), .A0N(\ram[181][11] ), .A1N(n6429), 
        .Y(n3489) );
  OAI2BB2XL U3466 ( .B0(n6681), .B1(n511), .A0N(\ram[181][12] ), .A1N(n6429), 
        .Y(n3490) );
  OAI2BB2XL U3467 ( .B0(n6658), .B1(n511), .A0N(\ram[181][13] ), .A1N(n6429), 
        .Y(n3491) );
  OAI2BB2XL U3468 ( .B0(n6635), .B1(n511), .A0N(\ram[181][14] ), .A1N(n6429), 
        .Y(n3492) );
  OAI2BB2XL U3469 ( .B0(n6612), .B1(n511), .A0N(\ram[181][15] ), .A1N(n6429), 
        .Y(n3493) );
  OAI2BB2XL U3470 ( .B0(n6965), .B1(n513), .A0N(\ram[182][0] ), .A1N(n6428), 
        .Y(n3494) );
  OAI2BB2XL U3471 ( .B0(n6942), .B1(n513), .A0N(\ram[182][1] ), .A1N(n6428), 
        .Y(n3495) );
  OAI2BB2XL U3472 ( .B0(n6919), .B1(n513), .A0N(\ram[182][2] ), .A1N(n6428), 
        .Y(n3496) );
  OAI2BB2XL U3473 ( .B0(n6896), .B1(n513), .A0N(\ram[182][3] ), .A1N(n6428), 
        .Y(n3497) );
  OAI2BB2XL U3474 ( .B0(n6866), .B1(n513), .A0N(\ram[182][4] ), .A1N(n6428), 
        .Y(n3498) );
  OAI2BB2XL U3475 ( .B0(n6843), .B1(n513), .A0N(\ram[182][5] ), .A1N(n6428), 
        .Y(n3499) );
  OAI2BB2XL U3476 ( .B0(n6820), .B1(n513), .A0N(\ram[182][6] ), .A1N(n6428), 
        .Y(n3500) );
  OAI2BB2XL U3477 ( .B0(n6797), .B1(n513), .A0N(\ram[182][7] ), .A1N(n6428), 
        .Y(n3501) );
  OAI2BB2XL U3478 ( .B0(n6774), .B1(n513), .A0N(\ram[182][8] ), .A1N(n6428), 
        .Y(n3502) );
  OAI2BB2XL U3479 ( .B0(n6751), .B1(n513), .A0N(\ram[182][9] ), .A1N(n6428), 
        .Y(n3503) );
  OAI2BB2XL U3480 ( .B0(n6728), .B1(n513), .A0N(\ram[182][10] ), .A1N(n6428), 
        .Y(n3504) );
  OAI2BB2XL U3481 ( .B0(n6705), .B1(n513), .A0N(\ram[182][11] ), .A1N(n6428), 
        .Y(n3505) );
  OAI2BB2XL U3482 ( .B0(n6682), .B1(n513), .A0N(\ram[182][12] ), .A1N(n6428), 
        .Y(n3506) );
  OAI2BB2XL U3483 ( .B0(n6659), .B1(n513), .A0N(\ram[182][13] ), .A1N(n6428), 
        .Y(n3507) );
  OAI2BB2XL U3484 ( .B0(n6636), .B1(n513), .A0N(\ram[182][14] ), .A1N(n6428), 
        .Y(n3508) );
  OAI2BB2XL U3485 ( .B0(n6613), .B1(n513), .A0N(\ram[182][15] ), .A1N(n6428), 
        .Y(n3509) );
  OAI2BB2XL U3486 ( .B0(n6965), .B1(n515), .A0N(\ram[183][0] ), .A1N(n6427), 
        .Y(n3510) );
  OAI2BB2XL U3487 ( .B0(n6942), .B1(n515), .A0N(\ram[183][1] ), .A1N(n6427), 
        .Y(n3511) );
  OAI2BB2XL U3488 ( .B0(n6919), .B1(n515), .A0N(\ram[183][2] ), .A1N(n6427), 
        .Y(n3512) );
  OAI2BB2XL U3489 ( .B0(n6896), .B1(n515), .A0N(\ram[183][3] ), .A1N(n6427), 
        .Y(n3513) );
  OAI2BB2XL U3490 ( .B0(n6871), .B1(n515), .A0N(\ram[183][4] ), .A1N(n6427), 
        .Y(n3514) );
  OAI2BB2XL U3491 ( .B0(n6848), .B1(n515), .A0N(\ram[183][5] ), .A1N(n6427), 
        .Y(n3515) );
  OAI2BB2XL U3492 ( .B0(n6825), .B1(n515), .A0N(\ram[183][6] ), .A1N(n6427), 
        .Y(n3516) );
  OAI2BB2XL U3493 ( .B0(n6802), .B1(n515), .A0N(\ram[183][7] ), .A1N(n6427), 
        .Y(n3517) );
  OAI2BB2XL U3494 ( .B0(n6779), .B1(n515), .A0N(\ram[183][8] ), .A1N(n6427), 
        .Y(n3518) );
  OAI2BB2XL U3495 ( .B0(n6756), .B1(n515), .A0N(\ram[183][9] ), .A1N(n6427), 
        .Y(n3519) );
  OAI2BB2XL U3496 ( .B0(n6733), .B1(n515), .A0N(\ram[183][10] ), .A1N(n6427), 
        .Y(n3520) );
  OAI2BB2XL U3497 ( .B0(n6710), .B1(n515), .A0N(\ram[183][11] ), .A1N(n6427), 
        .Y(n3521) );
  OAI2BB2XL U3498 ( .B0(n6687), .B1(n515), .A0N(\ram[183][12] ), .A1N(n6427), 
        .Y(n3522) );
  OAI2BB2XL U3499 ( .B0(n6664), .B1(n515), .A0N(\ram[183][13] ), .A1N(n6427), 
        .Y(n3523) );
  OAI2BB2XL U3500 ( .B0(n6641), .B1(n515), .A0N(\ram[183][14] ), .A1N(n6427), 
        .Y(n3524) );
  OAI2BB2XL U3501 ( .B0(n6618), .B1(n515), .A0N(\ram[183][15] ), .A1N(n6427), 
        .Y(n3525) );
  OAI2BB2XL U3502 ( .B0(n6964), .B1(n345), .A0N(\ram[184][0] ), .A1N(n6426), 
        .Y(n3526) );
  OAI2BB2XL U3503 ( .B0(n6941), .B1(n345), .A0N(\ram[184][1] ), .A1N(n6426), 
        .Y(n3527) );
  OAI2BB2XL U3504 ( .B0(n6918), .B1(n345), .A0N(\ram[184][2] ), .A1N(n6426), 
        .Y(n3528) );
  OAI2BB2XL U3505 ( .B0(n6895), .B1(n345), .A0N(\ram[184][3] ), .A1N(n6426), 
        .Y(n3529) );
  OAI2BB2XL U3506 ( .B0(n6868), .B1(n345), .A0N(\ram[184][4] ), .A1N(n6426), 
        .Y(n3530) );
  OAI2BB2XL U3507 ( .B0(n6845), .B1(n345), .A0N(\ram[184][5] ), .A1N(n6426), 
        .Y(n3531) );
  OAI2BB2XL U3508 ( .B0(n6822), .B1(n345), .A0N(\ram[184][6] ), .A1N(n6426), 
        .Y(n3532) );
  OAI2BB2XL U3509 ( .B0(n6799), .B1(n345), .A0N(\ram[184][7] ), .A1N(n6426), 
        .Y(n3533) );
  OAI2BB2XL U3510 ( .B0(n6776), .B1(n345), .A0N(\ram[184][8] ), .A1N(n6426), 
        .Y(n3534) );
  OAI2BB2XL U3511 ( .B0(n6753), .B1(n345), .A0N(\ram[184][9] ), .A1N(n6426), 
        .Y(n3535) );
  OAI2BB2XL U3512 ( .B0(n6730), .B1(n345), .A0N(\ram[184][10] ), .A1N(n6426), 
        .Y(n3536) );
  OAI2BB2XL U3513 ( .B0(n6707), .B1(n345), .A0N(\ram[184][11] ), .A1N(n6426), 
        .Y(n3537) );
  OAI2BB2XL U3514 ( .B0(n6684), .B1(n345), .A0N(\ram[184][12] ), .A1N(n6426), 
        .Y(n3538) );
  OAI2BB2XL U3515 ( .B0(n6661), .B1(n345), .A0N(\ram[184][13] ), .A1N(n6426), 
        .Y(n3539) );
  OAI2BB2XL U3516 ( .B0(n6638), .B1(n345), .A0N(\ram[184][14] ), .A1N(n6426), 
        .Y(n3540) );
  OAI2BB2XL U3517 ( .B0(n6615), .B1(n345), .A0N(\ram[184][15] ), .A1N(n6426), 
        .Y(n3541) );
  OAI2BB2XL U3518 ( .B0(n6964), .B1(n347), .A0N(\ram[185][0] ), .A1N(n6425), 
        .Y(n3542) );
  OAI2BB2XL U3519 ( .B0(n6941), .B1(n347), .A0N(\ram[185][1] ), .A1N(n6425), 
        .Y(n3543) );
  OAI2BB2XL U3520 ( .B0(n6918), .B1(n347), .A0N(\ram[185][2] ), .A1N(n6425), 
        .Y(n3544) );
  OAI2BB2XL U3521 ( .B0(n6895), .B1(n347), .A0N(\ram[185][3] ), .A1N(n6425), 
        .Y(n3545) );
  OAI2BB2XL U3522 ( .B0(n6868), .B1(n347), .A0N(\ram[185][4] ), .A1N(n6425), 
        .Y(n3546) );
  OAI2BB2XL U3523 ( .B0(n6845), .B1(n347), .A0N(\ram[185][5] ), .A1N(n6425), 
        .Y(n3547) );
  OAI2BB2XL U3524 ( .B0(n6822), .B1(n347), .A0N(\ram[185][6] ), .A1N(n6425), 
        .Y(n3548) );
  OAI2BB2XL U3525 ( .B0(n6799), .B1(n347), .A0N(\ram[185][7] ), .A1N(n6425), 
        .Y(n3549) );
  OAI2BB2XL U3526 ( .B0(n6776), .B1(n347), .A0N(\ram[185][8] ), .A1N(n6425), 
        .Y(n3550) );
  OAI2BB2XL U3527 ( .B0(n6753), .B1(n347), .A0N(\ram[185][9] ), .A1N(n6425), 
        .Y(n3551) );
  OAI2BB2XL U3528 ( .B0(n6730), .B1(n347), .A0N(\ram[185][10] ), .A1N(n6425), 
        .Y(n3552) );
  OAI2BB2XL U3529 ( .B0(n6707), .B1(n347), .A0N(\ram[185][11] ), .A1N(n6425), 
        .Y(n3553) );
  OAI2BB2XL U3530 ( .B0(n6684), .B1(n347), .A0N(\ram[185][12] ), .A1N(n6425), 
        .Y(n3554) );
  OAI2BB2XL U3531 ( .B0(n6661), .B1(n347), .A0N(\ram[185][13] ), .A1N(n6425), 
        .Y(n3555) );
  OAI2BB2XL U3532 ( .B0(n6638), .B1(n347), .A0N(\ram[185][14] ), .A1N(n6425), 
        .Y(n3556) );
  OAI2BB2XL U3533 ( .B0(n6615), .B1(n347), .A0N(\ram[185][15] ), .A1N(n6425), 
        .Y(n3557) );
  OAI2BB2XL U3534 ( .B0(n6964), .B1(n349), .A0N(\ram[186][0] ), .A1N(n6424), 
        .Y(n3558) );
  OAI2BB2XL U3535 ( .B0(n6941), .B1(n349), .A0N(\ram[186][1] ), .A1N(n6424), 
        .Y(n3559) );
  OAI2BB2XL U3536 ( .B0(n6918), .B1(n349), .A0N(\ram[186][2] ), .A1N(n6424), 
        .Y(n3560) );
  OAI2BB2XL U3537 ( .B0(n6895), .B1(n349), .A0N(\ram[186][3] ), .A1N(n6424), 
        .Y(n3561) );
  OAI2BB2XL U3538 ( .B0(n6868), .B1(n349), .A0N(\ram[186][4] ), .A1N(n6424), 
        .Y(n3562) );
  OAI2BB2XL U3539 ( .B0(n6845), .B1(n349), .A0N(\ram[186][5] ), .A1N(n6424), 
        .Y(n3563) );
  OAI2BB2XL U3540 ( .B0(n6822), .B1(n349), .A0N(\ram[186][6] ), .A1N(n6424), 
        .Y(n3564) );
  OAI2BB2XL U3541 ( .B0(n6799), .B1(n349), .A0N(\ram[186][7] ), .A1N(n6424), 
        .Y(n3565) );
  OAI2BB2XL U3542 ( .B0(n6776), .B1(n349), .A0N(\ram[186][8] ), .A1N(n6424), 
        .Y(n3566) );
  OAI2BB2XL U3543 ( .B0(n6753), .B1(n349), .A0N(\ram[186][9] ), .A1N(n6424), 
        .Y(n3567) );
  OAI2BB2XL U3544 ( .B0(n6730), .B1(n349), .A0N(\ram[186][10] ), .A1N(n6424), 
        .Y(n3568) );
  OAI2BB2XL U3545 ( .B0(n6707), .B1(n349), .A0N(\ram[186][11] ), .A1N(n6424), 
        .Y(n3569) );
  OAI2BB2XL U3546 ( .B0(n6684), .B1(n349), .A0N(\ram[186][12] ), .A1N(n6424), 
        .Y(n3570) );
  OAI2BB2XL U3547 ( .B0(n6661), .B1(n349), .A0N(\ram[186][13] ), .A1N(n6424), 
        .Y(n3571) );
  OAI2BB2XL U3548 ( .B0(n6638), .B1(n349), .A0N(\ram[186][14] ), .A1N(n6424), 
        .Y(n3572) );
  OAI2BB2XL U3549 ( .B0(n6615), .B1(n349), .A0N(\ram[186][15] ), .A1N(n6424), 
        .Y(n3573) );
  OAI2BB2XL U3550 ( .B0(n6964), .B1(n351), .A0N(\ram[187][0] ), .A1N(n6423), 
        .Y(n3574) );
  OAI2BB2XL U3551 ( .B0(n6941), .B1(n351), .A0N(\ram[187][1] ), .A1N(n6423), 
        .Y(n3575) );
  OAI2BB2XL U3552 ( .B0(n6918), .B1(n351), .A0N(\ram[187][2] ), .A1N(n6423), 
        .Y(n3576) );
  OAI2BB2XL U3553 ( .B0(n6895), .B1(n351), .A0N(\ram[187][3] ), .A1N(n6423), 
        .Y(n3577) );
  OAI2BB2XL U3554 ( .B0(n6868), .B1(n351), .A0N(\ram[187][4] ), .A1N(n6423), 
        .Y(n3578) );
  OAI2BB2XL U3555 ( .B0(n6845), .B1(n351), .A0N(\ram[187][5] ), .A1N(n6423), 
        .Y(n3579) );
  OAI2BB2XL U3556 ( .B0(n6822), .B1(n351), .A0N(\ram[187][6] ), .A1N(n6423), 
        .Y(n3580) );
  OAI2BB2XL U3557 ( .B0(n6799), .B1(n351), .A0N(\ram[187][7] ), .A1N(n6423), 
        .Y(n3581) );
  OAI2BB2XL U3558 ( .B0(n6776), .B1(n351), .A0N(\ram[187][8] ), .A1N(n6423), 
        .Y(n3582) );
  OAI2BB2XL U3559 ( .B0(n6753), .B1(n351), .A0N(\ram[187][9] ), .A1N(n6423), 
        .Y(n3583) );
  OAI2BB2XL U3560 ( .B0(n6730), .B1(n351), .A0N(\ram[187][10] ), .A1N(n6423), 
        .Y(n3584) );
  OAI2BB2XL U3561 ( .B0(n6707), .B1(n351), .A0N(\ram[187][11] ), .A1N(n6423), 
        .Y(n3585) );
  OAI2BB2XL U3562 ( .B0(n6684), .B1(n351), .A0N(\ram[187][12] ), .A1N(n6423), 
        .Y(n3586) );
  OAI2BB2XL U3563 ( .B0(n6661), .B1(n351), .A0N(\ram[187][13] ), .A1N(n6423), 
        .Y(n3587) );
  OAI2BB2XL U3564 ( .B0(n6638), .B1(n351), .A0N(\ram[187][14] ), .A1N(n6423), 
        .Y(n3588) );
  OAI2BB2XL U3565 ( .B0(n6615), .B1(n351), .A0N(\ram[187][15] ), .A1N(n6423), 
        .Y(n3589) );
  OAI2BB2XL U3566 ( .B0(n6964), .B1(n353), .A0N(\ram[188][0] ), .A1N(n6422), 
        .Y(n3590) );
  OAI2BB2XL U3567 ( .B0(n6941), .B1(n353), .A0N(\ram[188][1] ), .A1N(n6422), 
        .Y(n3591) );
  OAI2BB2XL U3568 ( .B0(n6918), .B1(n353), .A0N(\ram[188][2] ), .A1N(n6422), 
        .Y(n3592) );
  OAI2BB2XL U3569 ( .B0(n6895), .B1(n353), .A0N(\ram[188][3] ), .A1N(n6422), 
        .Y(n3593) );
  OAI2BB2XL U3570 ( .B0(n6868), .B1(n353), .A0N(\ram[188][4] ), .A1N(n6422), 
        .Y(n3594) );
  OAI2BB2XL U3571 ( .B0(n6845), .B1(n353), .A0N(\ram[188][5] ), .A1N(n6422), 
        .Y(n3595) );
  OAI2BB2XL U3572 ( .B0(n6822), .B1(n353), .A0N(\ram[188][6] ), .A1N(n6422), 
        .Y(n3596) );
  OAI2BB2XL U3573 ( .B0(n6799), .B1(n353), .A0N(\ram[188][7] ), .A1N(n6422), 
        .Y(n3597) );
  OAI2BB2XL U3574 ( .B0(n6776), .B1(n353), .A0N(\ram[188][8] ), .A1N(n6422), 
        .Y(n3598) );
  OAI2BB2XL U3575 ( .B0(n6753), .B1(n353), .A0N(\ram[188][9] ), .A1N(n6422), 
        .Y(n3599) );
  OAI2BB2XL U3576 ( .B0(n6730), .B1(n353), .A0N(\ram[188][10] ), .A1N(n6422), 
        .Y(n3600) );
  OAI2BB2XL U3577 ( .B0(n6707), .B1(n353), .A0N(\ram[188][11] ), .A1N(n6422), 
        .Y(n3601) );
  OAI2BB2XL U3578 ( .B0(n6684), .B1(n353), .A0N(\ram[188][12] ), .A1N(n6422), 
        .Y(n3602) );
  OAI2BB2XL U3579 ( .B0(n6661), .B1(n353), .A0N(\ram[188][13] ), .A1N(n6422), 
        .Y(n3603) );
  OAI2BB2XL U3580 ( .B0(n6638), .B1(n353), .A0N(\ram[188][14] ), .A1N(n6422), 
        .Y(n3604) );
  OAI2BB2XL U3581 ( .B0(n6615), .B1(n353), .A0N(\ram[188][15] ), .A1N(n6422), 
        .Y(n3605) );
  OAI2BB2XL U3582 ( .B0(n6964), .B1(n355), .A0N(\ram[189][0] ), .A1N(n6421), 
        .Y(n3606) );
  OAI2BB2XL U3583 ( .B0(n6941), .B1(n355), .A0N(\ram[189][1] ), .A1N(n6421), 
        .Y(n3607) );
  OAI2BB2XL U3584 ( .B0(n6918), .B1(n355), .A0N(\ram[189][2] ), .A1N(n6421), 
        .Y(n3608) );
  OAI2BB2XL U3585 ( .B0(n6895), .B1(n355), .A0N(\ram[189][3] ), .A1N(n6421), 
        .Y(n3609) );
  OAI2BB2XL U3586 ( .B0(n6868), .B1(n355), .A0N(\ram[189][4] ), .A1N(n6421), 
        .Y(n3610) );
  OAI2BB2XL U3587 ( .B0(n6845), .B1(n355), .A0N(\ram[189][5] ), .A1N(n6421), 
        .Y(n3611) );
  OAI2BB2XL U3588 ( .B0(n6822), .B1(n355), .A0N(\ram[189][6] ), .A1N(n6421), 
        .Y(n3612) );
  OAI2BB2XL U3589 ( .B0(n6799), .B1(n355), .A0N(\ram[189][7] ), .A1N(n6421), 
        .Y(n3613) );
  OAI2BB2XL U3590 ( .B0(n6776), .B1(n355), .A0N(\ram[189][8] ), .A1N(n6421), 
        .Y(n3614) );
  OAI2BB2XL U3591 ( .B0(n6753), .B1(n355), .A0N(\ram[189][9] ), .A1N(n6421), 
        .Y(n3615) );
  OAI2BB2XL U3592 ( .B0(n6730), .B1(n355), .A0N(\ram[189][10] ), .A1N(n6421), 
        .Y(n3616) );
  OAI2BB2XL U3593 ( .B0(n6707), .B1(n355), .A0N(\ram[189][11] ), .A1N(n6421), 
        .Y(n3617) );
  OAI2BB2XL U3594 ( .B0(n6684), .B1(n355), .A0N(\ram[189][12] ), .A1N(n6421), 
        .Y(n3618) );
  OAI2BB2XL U3595 ( .B0(n6661), .B1(n355), .A0N(\ram[189][13] ), .A1N(n6421), 
        .Y(n3619) );
  OAI2BB2XL U3596 ( .B0(n6638), .B1(n355), .A0N(\ram[189][14] ), .A1N(n6421), 
        .Y(n3620) );
  OAI2BB2XL U3597 ( .B0(n6615), .B1(n355), .A0N(\ram[189][15] ), .A1N(n6421), 
        .Y(n3621) );
  OAI2BB2XL U3598 ( .B0(n6964), .B1(n357), .A0N(\ram[190][0] ), .A1N(n6420), 
        .Y(n3622) );
  OAI2BB2XL U3599 ( .B0(n6941), .B1(n357), .A0N(\ram[190][1] ), .A1N(n6420), 
        .Y(n3623) );
  OAI2BB2XL U3600 ( .B0(n6918), .B1(n357), .A0N(\ram[190][2] ), .A1N(n6420), 
        .Y(n3624) );
  OAI2BB2XL U3601 ( .B0(n6895), .B1(n357), .A0N(\ram[190][3] ), .A1N(n6420), 
        .Y(n3625) );
  OAI2BB2XL U3602 ( .B0(n6868), .B1(n357), .A0N(\ram[190][4] ), .A1N(n6420), 
        .Y(n3626) );
  OAI2BB2XL U3603 ( .B0(n6845), .B1(n357), .A0N(\ram[190][5] ), .A1N(n6420), 
        .Y(n3627) );
  OAI2BB2XL U3604 ( .B0(n6822), .B1(n357), .A0N(\ram[190][6] ), .A1N(n6420), 
        .Y(n3628) );
  OAI2BB2XL U3605 ( .B0(n6799), .B1(n357), .A0N(\ram[190][7] ), .A1N(n6420), 
        .Y(n3629) );
  OAI2BB2XL U3606 ( .B0(n6776), .B1(n357), .A0N(\ram[190][8] ), .A1N(n6420), 
        .Y(n3630) );
  OAI2BB2XL U3607 ( .B0(n6753), .B1(n357), .A0N(\ram[190][9] ), .A1N(n6420), 
        .Y(n3631) );
  OAI2BB2XL U3608 ( .B0(n6730), .B1(n357), .A0N(\ram[190][10] ), .A1N(n6420), 
        .Y(n3632) );
  OAI2BB2XL U3609 ( .B0(n6707), .B1(n357), .A0N(\ram[190][11] ), .A1N(n6420), 
        .Y(n3633) );
  OAI2BB2XL U3610 ( .B0(n6684), .B1(n357), .A0N(\ram[190][12] ), .A1N(n6420), 
        .Y(n3634) );
  OAI2BB2XL U3611 ( .B0(n6661), .B1(n357), .A0N(\ram[190][13] ), .A1N(n6420), 
        .Y(n3635) );
  OAI2BB2XL U3612 ( .B0(n6638), .B1(n357), .A0N(\ram[190][14] ), .A1N(n6420), 
        .Y(n3636) );
  OAI2BB2XL U3613 ( .B0(n6615), .B1(n357), .A0N(\ram[190][15] ), .A1N(n6420), 
        .Y(n3637) );
  OAI2BB2XL U3614 ( .B0(n6964), .B1(n359), .A0N(\ram[191][0] ), .A1N(n6419), 
        .Y(n3638) );
  OAI2BB2XL U3615 ( .B0(n6941), .B1(n359), .A0N(\ram[191][1] ), .A1N(n6419), 
        .Y(n3639) );
  OAI2BB2XL U3616 ( .B0(n6918), .B1(n359), .A0N(\ram[191][2] ), .A1N(n6419), 
        .Y(n3640) );
  OAI2BB2XL U3617 ( .B0(n6895), .B1(n359), .A0N(\ram[191][3] ), .A1N(n6419), 
        .Y(n3641) );
  OAI2BB2XL U3618 ( .B0(n6868), .B1(n359), .A0N(\ram[191][4] ), .A1N(n6419), 
        .Y(n3642) );
  OAI2BB2XL U3619 ( .B0(n6845), .B1(n359), .A0N(\ram[191][5] ), .A1N(n6419), 
        .Y(n3643) );
  OAI2BB2XL U3620 ( .B0(n6822), .B1(n359), .A0N(\ram[191][6] ), .A1N(n6419), 
        .Y(n3644) );
  OAI2BB2XL U3621 ( .B0(n6799), .B1(n359), .A0N(\ram[191][7] ), .A1N(n6419), 
        .Y(n3645) );
  OAI2BB2XL U3622 ( .B0(n6776), .B1(n359), .A0N(\ram[191][8] ), .A1N(n6419), 
        .Y(n3646) );
  OAI2BB2XL U3623 ( .B0(n6753), .B1(n359), .A0N(\ram[191][9] ), .A1N(n6419), 
        .Y(n3647) );
  OAI2BB2XL U3624 ( .B0(n6730), .B1(n359), .A0N(\ram[191][10] ), .A1N(n6419), 
        .Y(n3648) );
  OAI2BB2XL U3625 ( .B0(n6707), .B1(n359), .A0N(\ram[191][11] ), .A1N(n6419), 
        .Y(n3649) );
  OAI2BB2XL U3626 ( .B0(n6684), .B1(n359), .A0N(\ram[191][12] ), .A1N(n6419), 
        .Y(n3650) );
  OAI2BB2XL U3627 ( .B0(n6661), .B1(n359), .A0N(\ram[191][13] ), .A1N(n6419), 
        .Y(n3651) );
  OAI2BB2XL U3628 ( .B0(n6638), .B1(n359), .A0N(\ram[191][14] ), .A1N(n6419), 
        .Y(n3652) );
  OAI2BB2XL U3629 ( .B0(n6615), .B1(n359), .A0N(\ram[191][15] ), .A1N(n6419), 
        .Y(n3653) );
  OAI2BB2XL U3630 ( .B0(n6962), .B1(n392), .A0N(\ram[208][0] ), .A1N(n6402), 
        .Y(n3910) );
  OAI2BB2XL U3631 ( .B0(n6939), .B1(n392), .A0N(\ram[208][1] ), .A1N(n6402), 
        .Y(n3911) );
  OAI2BB2XL U3632 ( .B0(n6916), .B1(n392), .A0N(\ram[208][2] ), .A1N(n6402), 
        .Y(n3912) );
  OAI2BB2XL U3633 ( .B0(n6893), .B1(n392), .A0N(\ram[208][3] ), .A1N(n6402), 
        .Y(n3913) );
  OAI2BB2XL U3634 ( .B0(n6872), .B1(n392), .A0N(\ram[208][4] ), .A1N(n6402), 
        .Y(n3914) );
  OAI2BB2XL U3635 ( .B0(n6849), .B1(n392), .A0N(\ram[208][5] ), .A1N(n6402), 
        .Y(n3915) );
  OAI2BB2XL U3636 ( .B0(n6826), .B1(n392), .A0N(\ram[208][6] ), .A1N(n6402), 
        .Y(n3916) );
  OAI2BB2XL U3637 ( .B0(n6803), .B1(n392), .A0N(\ram[208][7] ), .A1N(n6402), 
        .Y(n3917) );
  OAI2BB2XL U3638 ( .B0(n6780), .B1(n392), .A0N(\ram[208][8] ), .A1N(n6402), 
        .Y(n3918) );
  OAI2BB2XL U3639 ( .B0(n6757), .B1(n392), .A0N(\ram[208][9] ), .A1N(n6402), 
        .Y(n3919) );
  OAI2BB2XL U3640 ( .B0(n6734), .B1(n392), .A0N(\ram[208][10] ), .A1N(n6402), 
        .Y(n3920) );
  OAI2BB2XL U3641 ( .B0(n6711), .B1(n392), .A0N(\ram[208][11] ), .A1N(n6402), 
        .Y(n3921) );
  OAI2BB2XL U3642 ( .B0(n6688), .B1(n392), .A0N(\ram[208][12] ), .A1N(n6402), 
        .Y(n3922) );
  OAI2BB2XL U3643 ( .B0(n6665), .B1(n392), .A0N(\ram[208][13] ), .A1N(n6402), 
        .Y(n3923) );
  OAI2BB2XL U3644 ( .B0(n6642), .B1(n392), .A0N(\ram[208][14] ), .A1N(n6402), 
        .Y(n3924) );
  OAI2BB2XL U3645 ( .B0(n6619), .B1(n392), .A0N(\ram[208][15] ), .A1N(n6402), 
        .Y(n3925) );
  OAI2BB2XL U3646 ( .B0(n6962), .B1(n394), .A0N(\ram[209][0] ), .A1N(n6401), 
        .Y(n3926) );
  OAI2BB2XL U3647 ( .B0(n6939), .B1(n394), .A0N(\ram[209][1] ), .A1N(n6401), 
        .Y(n3927) );
  OAI2BB2XL U3648 ( .B0(n6916), .B1(n394), .A0N(\ram[209][2] ), .A1N(n6401), 
        .Y(n3928) );
  OAI2BB2XL U3649 ( .B0(n6893), .B1(n394), .A0N(\ram[209][3] ), .A1N(n6401), 
        .Y(n3929) );
  OAI2BB2XL U3650 ( .B0(n6875), .B1(n394), .A0N(\ram[209][4] ), .A1N(n6401), 
        .Y(n3930) );
  OAI2BB2XL U3651 ( .B0(n6852), .B1(n394), .A0N(\ram[209][5] ), .A1N(n6401), 
        .Y(n3931) );
  OAI2BB2XL U3652 ( .B0(n6829), .B1(n394), .A0N(\ram[209][6] ), .A1N(n6401), 
        .Y(n3932) );
  OAI2BB2XL U3653 ( .B0(n6806), .B1(n394), .A0N(\ram[209][7] ), .A1N(n6401), 
        .Y(n3933) );
  OAI2BB2XL U3654 ( .B0(n6783), .B1(n394), .A0N(\ram[209][8] ), .A1N(n6401), 
        .Y(n3934) );
  OAI2BB2XL U3655 ( .B0(n6760), .B1(n394), .A0N(\ram[209][9] ), .A1N(n6401), 
        .Y(n3935) );
  OAI2BB2XL U3656 ( .B0(n6737), .B1(n394), .A0N(\ram[209][10] ), .A1N(n6401), 
        .Y(n3936) );
  OAI2BB2XL U3657 ( .B0(n6714), .B1(n394), .A0N(\ram[209][11] ), .A1N(n6401), 
        .Y(n3937) );
  OAI2BB2XL U3658 ( .B0(n6691), .B1(n394), .A0N(\ram[209][12] ), .A1N(n6401), 
        .Y(n3938) );
  OAI2BB2XL U3659 ( .B0(n6668), .B1(n394), .A0N(\ram[209][13] ), .A1N(n6401), 
        .Y(n3939) );
  OAI2BB2XL U3660 ( .B0(n6645), .B1(n394), .A0N(\ram[209][14] ), .A1N(n6401), 
        .Y(n3940) );
  OAI2BB2XL U3661 ( .B0(n6622), .B1(n394), .A0N(\ram[209][15] ), .A1N(n6401), 
        .Y(n3941) );
  OAI2BB2XL U3662 ( .B0(n6962), .B1(n396), .A0N(\ram[210][0] ), .A1N(n6400), 
        .Y(n3942) );
  OAI2BB2XL U3663 ( .B0(n6939), .B1(n396), .A0N(\ram[210][1] ), .A1N(n6400), 
        .Y(n3943) );
  OAI2BB2XL U3664 ( .B0(n6916), .B1(n396), .A0N(\ram[210][2] ), .A1N(n6400), 
        .Y(n3944) );
  OAI2BB2XL U3665 ( .B0(n6893), .B1(n396), .A0N(\ram[210][3] ), .A1N(n6400), 
        .Y(n3945) );
  OAI2BB2XL U3666 ( .B0(n6874), .B1(n396), .A0N(\ram[210][4] ), .A1N(n6400), 
        .Y(n3946) );
  OAI2BB2XL U3667 ( .B0(n6851), .B1(n396), .A0N(\ram[210][5] ), .A1N(n6400), 
        .Y(n3947) );
  OAI2BB2XL U3668 ( .B0(n6828), .B1(n396), .A0N(\ram[210][6] ), .A1N(n6400), 
        .Y(n3948) );
  OAI2BB2XL U3669 ( .B0(n6805), .B1(n396), .A0N(\ram[210][7] ), .A1N(n6400), 
        .Y(n3949) );
  OAI2BB2XL U3670 ( .B0(n6782), .B1(n396), .A0N(\ram[210][8] ), .A1N(n6400), 
        .Y(n3950) );
  OAI2BB2XL U3671 ( .B0(n6759), .B1(n396), .A0N(\ram[210][9] ), .A1N(n6400), 
        .Y(n3951) );
  OAI2BB2XL U3672 ( .B0(n6736), .B1(n396), .A0N(\ram[210][10] ), .A1N(n6400), 
        .Y(n3952) );
  OAI2BB2XL U3673 ( .B0(n6713), .B1(n396), .A0N(\ram[210][11] ), .A1N(n6400), 
        .Y(n3953) );
  OAI2BB2XL U3674 ( .B0(n6690), .B1(n396), .A0N(\ram[210][12] ), .A1N(n6400), 
        .Y(n3954) );
  OAI2BB2XL U3675 ( .B0(n6667), .B1(n396), .A0N(\ram[210][13] ), .A1N(n6400), 
        .Y(n3955) );
  OAI2BB2XL U3676 ( .B0(n6644), .B1(n396), .A0N(\ram[210][14] ), .A1N(n6400), 
        .Y(n3956) );
  OAI2BB2XL U3677 ( .B0(n6621), .B1(n396), .A0N(\ram[210][15] ), .A1N(n6400), 
        .Y(n3957) );
  OAI2BB2XL U3678 ( .B0(n6962), .B1(n398), .A0N(\ram[211][0] ), .A1N(n6399), 
        .Y(n3958) );
  OAI2BB2XL U3679 ( .B0(n6939), .B1(n398), .A0N(\ram[211][1] ), .A1N(n6399), 
        .Y(n3959) );
  OAI2BB2XL U3680 ( .B0(n6916), .B1(n398), .A0N(\ram[211][2] ), .A1N(n6399), 
        .Y(n3960) );
  OAI2BB2XL U3681 ( .B0(n6893), .B1(n398), .A0N(\ram[211][3] ), .A1N(n6399), 
        .Y(n3961) );
  OAI2BB2XL U3682 ( .B0(n6872), .B1(n398), .A0N(\ram[211][4] ), .A1N(n6399), 
        .Y(n3962) );
  OAI2BB2XL U3683 ( .B0(n6849), .B1(n398), .A0N(\ram[211][5] ), .A1N(n6399), 
        .Y(n3963) );
  OAI2BB2XL U3684 ( .B0(n6826), .B1(n398), .A0N(\ram[211][6] ), .A1N(n6399), 
        .Y(n3964) );
  OAI2BB2XL U3685 ( .B0(n6803), .B1(n398), .A0N(\ram[211][7] ), .A1N(n6399), 
        .Y(n3965) );
  OAI2BB2XL U3686 ( .B0(n6780), .B1(n398), .A0N(\ram[211][8] ), .A1N(n6399), 
        .Y(n3966) );
  OAI2BB2XL U3687 ( .B0(n6757), .B1(n398), .A0N(\ram[211][9] ), .A1N(n6399), 
        .Y(n3967) );
  OAI2BB2XL U3688 ( .B0(n6734), .B1(n398), .A0N(\ram[211][10] ), .A1N(n6399), 
        .Y(n3968) );
  OAI2BB2XL U3689 ( .B0(n6711), .B1(n398), .A0N(\ram[211][11] ), .A1N(n6399), 
        .Y(n3969) );
  OAI2BB2XL U3690 ( .B0(n6688), .B1(n398), .A0N(\ram[211][12] ), .A1N(n6399), 
        .Y(n3970) );
  OAI2BB2XL U3691 ( .B0(n6665), .B1(n398), .A0N(\ram[211][13] ), .A1N(n6399), 
        .Y(n3971) );
  OAI2BB2XL U3692 ( .B0(n6642), .B1(n398), .A0N(\ram[211][14] ), .A1N(n6399), 
        .Y(n3972) );
  OAI2BB2XL U3693 ( .B0(n6619), .B1(n398), .A0N(\ram[211][15] ), .A1N(n6399), 
        .Y(n3973) );
  OAI2BB2XL U3694 ( .B0(n6962), .B1(n400), .A0N(\ram[212][0] ), .A1N(n6398), 
        .Y(n3974) );
  OAI2BB2XL U3695 ( .B0(n6939), .B1(n400), .A0N(\ram[212][1] ), .A1N(n6398), 
        .Y(n3975) );
  OAI2BB2XL U3696 ( .B0(n6916), .B1(n400), .A0N(\ram[212][2] ), .A1N(n6398), 
        .Y(n3976) );
  OAI2BB2XL U3697 ( .B0(n6893), .B1(n400), .A0N(\ram[212][3] ), .A1N(n6398), 
        .Y(n3977) );
  OAI2BB2XL U3698 ( .B0(n6875), .B1(n400), .A0N(\ram[212][4] ), .A1N(n6398), 
        .Y(n3978) );
  OAI2BB2XL U3699 ( .B0(n6852), .B1(n400), .A0N(\ram[212][5] ), .A1N(n6398), 
        .Y(n3979) );
  OAI2BB2XL U3700 ( .B0(n6829), .B1(n400), .A0N(\ram[212][6] ), .A1N(n6398), 
        .Y(n3980) );
  OAI2BB2XL U3701 ( .B0(n6806), .B1(n400), .A0N(\ram[212][7] ), .A1N(n6398), 
        .Y(n3981) );
  OAI2BB2XL U3702 ( .B0(n6783), .B1(n400), .A0N(\ram[212][8] ), .A1N(n6398), 
        .Y(n3982) );
  OAI2BB2XL U3703 ( .B0(n6760), .B1(n400), .A0N(\ram[212][9] ), .A1N(n6398), 
        .Y(n3983) );
  OAI2BB2XL U3704 ( .B0(n6737), .B1(n400), .A0N(\ram[212][10] ), .A1N(n6398), 
        .Y(n3984) );
  OAI2BB2XL U3705 ( .B0(n6714), .B1(n400), .A0N(\ram[212][11] ), .A1N(n6398), 
        .Y(n3985) );
  OAI2BB2XL U3706 ( .B0(n6691), .B1(n400), .A0N(\ram[212][12] ), .A1N(n6398), 
        .Y(n3986) );
  OAI2BB2XL U3707 ( .B0(n6668), .B1(n400), .A0N(\ram[212][13] ), .A1N(n6398), 
        .Y(n3987) );
  OAI2BB2XL U3708 ( .B0(n6645), .B1(n400), .A0N(\ram[212][14] ), .A1N(n6398), 
        .Y(n3988) );
  OAI2BB2XL U3709 ( .B0(n6622), .B1(n400), .A0N(\ram[212][15] ), .A1N(n6398), 
        .Y(n3989) );
  OAI2BB2XL U3710 ( .B0(n6962), .B1(n402), .A0N(\ram[213][0] ), .A1N(n6397), 
        .Y(n3990) );
  OAI2BB2XL U3711 ( .B0(n6939), .B1(n402), .A0N(\ram[213][1] ), .A1N(n6397), 
        .Y(n3991) );
  OAI2BB2XL U3712 ( .B0(n6916), .B1(n402), .A0N(\ram[213][2] ), .A1N(n6397), 
        .Y(n3992) );
  OAI2BB2XL U3713 ( .B0(n6893), .B1(n402), .A0N(\ram[213][3] ), .A1N(n6397), 
        .Y(n3993) );
  OAI2BB2XL U3714 ( .B0(n6874), .B1(n402), .A0N(\ram[213][4] ), .A1N(n6397), 
        .Y(n3994) );
  OAI2BB2XL U3715 ( .B0(n6851), .B1(n402), .A0N(\ram[213][5] ), .A1N(n6397), 
        .Y(n3995) );
  OAI2BB2XL U3716 ( .B0(n6828), .B1(n402), .A0N(\ram[213][6] ), .A1N(n6397), 
        .Y(n3996) );
  OAI2BB2XL U3717 ( .B0(n6805), .B1(n402), .A0N(\ram[213][7] ), .A1N(n6397), 
        .Y(n3997) );
  OAI2BB2XL U3718 ( .B0(n6782), .B1(n402), .A0N(\ram[213][8] ), .A1N(n6397), 
        .Y(n3998) );
  OAI2BB2XL U3719 ( .B0(n6759), .B1(n402), .A0N(\ram[213][9] ), .A1N(n6397), 
        .Y(n3999) );
  OAI2BB2XL U3720 ( .B0(n6736), .B1(n402), .A0N(\ram[213][10] ), .A1N(n6397), 
        .Y(n4000) );
  OAI2BB2XL U3721 ( .B0(n6713), .B1(n402), .A0N(\ram[213][11] ), .A1N(n6397), 
        .Y(n4001) );
  OAI2BB2XL U3722 ( .B0(n6690), .B1(n402), .A0N(\ram[213][12] ), .A1N(n6397), 
        .Y(n4002) );
  OAI2BB2XL U3723 ( .B0(n6667), .B1(n402), .A0N(\ram[213][13] ), .A1N(n6397), 
        .Y(n4003) );
  OAI2BB2XL U3724 ( .B0(n6644), .B1(n402), .A0N(\ram[213][14] ), .A1N(n6397), 
        .Y(n4004) );
  OAI2BB2XL U3725 ( .B0(n6621), .B1(n402), .A0N(\ram[213][15] ), .A1N(n6397), 
        .Y(n4005) );
  OAI2BB2XL U3726 ( .B0(n6962), .B1(n404), .A0N(\ram[214][0] ), .A1N(n6396), 
        .Y(n4006) );
  OAI2BB2XL U3727 ( .B0(n6939), .B1(n404), .A0N(\ram[214][1] ), .A1N(n6396), 
        .Y(n4007) );
  OAI2BB2XL U3728 ( .B0(n6916), .B1(n404), .A0N(\ram[214][2] ), .A1N(n6396), 
        .Y(n4008) );
  OAI2BB2XL U3729 ( .B0(n6893), .B1(n404), .A0N(\ram[214][3] ), .A1N(n6396), 
        .Y(n4009) );
  OAI2BB2XL U3730 ( .B0(n6872), .B1(n404), .A0N(\ram[214][4] ), .A1N(n6396), 
        .Y(n4010) );
  OAI2BB2XL U3731 ( .B0(n6849), .B1(n404), .A0N(\ram[214][5] ), .A1N(n6396), 
        .Y(n4011) );
  OAI2BB2XL U3732 ( .B0(n6826), .B1(n404), .A0N(\ram[214][6] ), .A1N(n6396), 
        .Y(n4012) );
  OAI2BB2XL U3733 ( .B0(n6803), .B1(n404), .A0N(\ram[214][7] ), .A1N(n6396), 
        .Y(n4013) );
  OAI2BB2XL U3734 ( .B0(n6780), .B1(n404), .A0N(\ram[214][8] ), .A1N(n6396), 
        .Y(n4014) );
  OAI2BB2XL U3735 ( .B0(n6757), .B1(n404), .A0N(\ram[214][9] ), .A1N(n6396), 
        .Y(n4015) );
  OAI2BB2XL U3736 ( .B0(n6734), .B1(n404), .A0N(\ram[214][10] ), .A1N(n6396), 
        .Y(n4016) );
  OAI2BB2XL U3737 ( .B0(n6711), .B1(n404), .A0N(\ram[214][11] ), .A1N(n6396), 
        .Y(n4017) );
  OAI2BB2XL U3738 ( .B0(n6688), .B1(n404), .A0N(\ram[214][12] ), .A1N(n6396), 
        .Y(n4018) );
  OAI2BB2XL U3739 ( .B0(n6665), .B1(n404), .A0N(\ram[214][13] ), .A1N(n6396), 
        .Y(n4019) );
  OAI2BB2XL U3740 ( .B0(n6642), .B1(n404), .A0N(\ram[214][14] ), .A1N(n6396), 
        .Y(n4020) );
  OAI2BB2XL U3741 ( .B0(n6619), .B1(n404), .A0N(\ram[214][15] ), .A1N(n6396), 
        .Y(n4021) );
  OAI2BB2XL U3742 ( .B0(n6962), .B1(n406), .A0N(\ram[215][0] ), .A1N(n6395), 
        .Y(n4022) );
  OAI2BB2XL U3743 ( .B0(n6939), .B1(n406), .A0N(\ram[215][1] ), .A1N(n6395), 
        .Y(n4023) );
  OAI2BB2XL U3744 ( .B0(n6916), .B1(n406), .A0N(\ram[215][2] ), .A1N(n6395), 
        .Y(n4024) );
  OAI2BB2XL U3745 ( .B0(n6893), .B1(n406), .A0N(\ram[215][3] ), .A1N(n6395), 
        .Y(n4025) );
  OAI2BB2XL U3746 ( .B0(n6875), .B1(n406), .A0N(\ram[215][4] ), .A1N(n6395), 
        .Y(n4026) );
  OAI2BB2XL U3747 ( .B0(n6852), .B1(n406), .A0N(\ram[215][5] ), .A1N(n6395), 
        .Y(n4027) );
  OAI2BB2XL U3748 ( .B0(n6829), .B1(n406), .A0N(\ram[215][6] ), .A1N(n6395), 
        .Y(n4028) );
  OAI2BB2XL U3749 ( .B0(n6806), .B1(n406), .A0N(\ram[215][7] ), .A1N(n6395), 
        .Y(n4029) );
  OAI2BB2XL U3750 ( .B0(n6783), .B1(n406), .A0N(\ram[215][8] ), .A1N(n6395), 
        .Y(n4030) );
  OAI2BB2XL U3751 ( .B0(n6760), .B1(n406), .A0N(\ram[215][9] ), .A1N(n6395), 
        .Y(n4031) );
  OAI2BB2XL U3752 ( .B0(n6737), .B1(n406), .A0N(\ram[215][10] ), .A1N(n6395), 
        .Y(n4032) );
  OAI2BB2XL U3753 ( .B0(n6714), .B1(n406), .A0N(\ram[215][11] ), .A1N(n6395), 
        .Y(n4033) );
  OAI2BB2XL U3754 ( .B0(n6691), .B1(n406), .A0N(\ram[215][12] ), .A1N(n6395), 
        .Y(n4034) );
  OAI2BB2XL U3755 ( .B0(n6668), .B1(n406), .A0N(\ram[215][13] ), .A1N(n6395), 
        .Y(n4035) );
  OAI2BB2XL U3756 ( .B0(n6645), .B1(n406), .A0N(\ram[215][14] ), .A1N(n6395), 
        .Y(n4036) );
  OAI2BB2XL U3757 ( .B0(n6622), .B1(n406), .A0N(\ram[215][15] ), .A1N(n6395), 
        .Y(n4037) );
  OAI2BB2XL U3758 ( .B0(n6962), .B1(n408), .A0N(\ram[216][0] ), .A1N(n6394), 
        .Y(n4038) );
  OAI2BB2XL U3759 ( .B0(n6939), .B1(n408), .A0N(\ram[216][1] ), .A1N(n6394), 
        .Y(n4039) );
  OAI2BB2XL U3760 ( .B0(n6916), .B1(n408), .A0N(\ram[216][2] ), .A1N(n6394), 
        .Y(n4040) );
  OAI2BB2XL U3761 ( .B0(n6893), .B1(n408), .A0N(\ram[216][3] ), .A1N(n6394), 
        .Y(n4041) );
  OAI2BB2XL U3762 ( .B0(n6874), .B1(n408), .A0N(\ram[216][4] ), .A1N(n6394), 
        .Y(n4042) );
  OAI2BB2XL U3763 ( .B0(n6851), .B1(n408), .A0N(\ram[216][5] ), .A1N(n6394), 
        .Y(n4043) );
  OAI2BB2XL U3764 ( .B0(n6828), .B1(n408), .A0N(\ram[216][6] ), .A1N(n6394), 
        .Y(n4044) );
  OAI2BB2XL U3765 ( .B0(n6805), .B1(n408), .A0N(\ram[216][7] ), .A1N(n6394), 
        .Y(n4045) );
  OAI2BB2XL U3766 ( .B0(n6782), .B1(n408), .A0N(\ram[216][8] ), .A1N(n6394), 
        .Y(n4046) );
  OAI2BB2XL U3767 ( .B0(n6759), .B1(n408), .A0N(\ram[216][9] ), .A1N(n6394), 
        .Y(n4047) );
  OAI2BB2XL U3768 ( .B0(n6736), .B1(n408), .A0N(\ram[216][10] ), .A1N(n6394), 
        .Y(n4048) );
  OAI2BB2XL U3769 ( .B0(n6713), .B1(n408), .A0N(\ram[216][11] ), .A1N(n6394), 
        .Y(n4049) );
  OAI2BB2XL U3770 ( .B0(n6690), .B1(n408), .A0N(\ram[216][12] ), .A1N(n6394), 
        .Y(n4050) );
  OAI2BB2XL U3771 ( .B0(n6667), .B1(n408), .A0N(\ram[216][13] ), .A1N(n6394), 
        .Y(n4051) );
  OAI2BB2XL U3772 ( .B0(n6644), .B1(n408), .A0N(\ram[216][14] ), .A1N(n6394), 
        .Y(n4052) );
  OAI2BB2XL U3773 ( .B0(n6621), .B1(n408), .A0N(\ram[216][15] ), .A1N(n6394), 
        .Y(n4053) );
  OAI2BB2XL U3774 ( .B0(n6962), .B1(n410), .A0N(\ram[217][0] ), .A1N(n6393), 
        .Y(n4054) );
  OAI2BB2XL U3775 ( .B0(n6939), .B1(n410), .A0N(\ram[217][1] ), .A1N(n6393), 
        .Y(n4055) );
  OAI2BB2XL U3776 ( .B0(n6916), .B1(n410), .A0N(\ram[217][2] ), .A1N(n6393), 
        .Y(n4056) );
  OAI2BB2XL U3777 ( .B0(n6893), .B1(n410), .A0N(\ram[217][3] ), .A1N(n6393), 
        .Y(n4057) );
  OAI2BB2XL U3778 ( .B0(n6868), .B1(n410), .A0N(\ram[217][4] ), .A1N(n6393), 
        .Y(n4058) );
  OAI2BB2XL U3779 ( .B0(n6845), .B1(n410), .A0N(\ram[217][5] ), .A1N(n6393), 
        .Y(n4059) );
  OAI2BB2XL U3780 ( .B0(n6822), .B1(n410), .A0N(\ram[217][6] ), .A1N(n6393), 
        .Y(n4060) );
  OAI2BB2XL U3781 ( .B0(n6799), .B1(n410), .A0N(\ram[217][7] ), .A1N(n6393), 
        .Y(n4061) );
  OAI2BB2XL U3782 ( .B0(n6776), .B1(n410), .A0N(\ram[217][8] ), .A1N(n6393), 
        .Y(n4062) );
  OAI2BB2XL U3783 ( .B0(n6753), .B1(n410), .A0N(\ram[217][9] ), .A1N(n6393), 
        .Y(n4063) );
  OAI2BB2XL U3784 ( .B0(n6730), .B1(n410), .A0N(\ram[217][10] ), .A1N(n6393), 
        .Y(n4064) );
  OAI2BB2XL U3785 ( .B0(n6707), .B1(n410), .A0N(\ram[217][11] ), .A1N(n6393), 
        .Y(n4065) );
  OAI2BB2XL U3786 ( .B0(n6684), .B1(n410), .A0N(\ram[217][12] ), .A1N(n6393), 
        .Y(n4066) );
  OAI2BB2XL U3787 ( .B0(n6661), .B1(n410), .A0N(\ram[217][13] ), .A1N(n6393), 
        .Y(n4067) );
  OAI2BB2XL U3788 ( .B0(n6638), .B1(n410), .A0N(\ram[217][14] ), .A1N(n6393), 
        .Y(n4068) );
  OAI2BB2XL U3789 ( .B0(n6615), .B1(n410), .A0N(\ram[217][15] ), .A1N(n6393), 
        .Y(n4069) );
  OAI2BB2XL U3790 ( .B0(n6962), .B1(n411), .A0N(\ram[218][0] ), .A1N(n6392), 
        .Y(n4070) );
  OAI2BB2XL U3791 ( .B0(n6939), .B1(n411), .A0N(\ram[218][1] ), .A1N(n6392), 
        .Y(n4071) );
  OAI2BB2XL U3792 ( .B0(n6916), .B1(n411), .A0N(\ram[218][2] ), .A1N(n6392), 
        .Y(n4072) );
  OAI2BB2XL U3793 ( .B0(n6893), .B1(n411), .A0N(\ram[218][3] ), .A1N(n6392), 
        .Y(n4073) );
  OAI2BB2XL U3794 ( .B0(n6867), .B1(n411), .A0N(\ram[218][4] ), .A1N(n6392), 
        .Y(n4074) );
  OAI2BB2XL U3795 ( .B0(n6844), .B1(n411), .A0N(\ram[218][5] ), .A1N(n6392), 
        .Y(n4075) );
  OAI2BB2XL U3796 ( .B0(n6821), .B1(n411), .A0N(\ram[218][6] ), .A1N(n6392), 
        .Y(n4076) );
  OAI2BB2XL U3797 ( .B0(n6798), .B1(n411), .A0N(\ram[218][7] ), .A1N(n6392), 
        .Y(n4077) );
  OAI2BB2XL U3798 ( .B0(n6775), .B1(n411), .A0N(\ram[218][8] ), .A1N(n6392), 
        .Y(n4078) );
  OAI2BB2XL U3799 ( .B0(n6752), .B1(n411), .A0N(\ram[218][9] ), .A1N(n6392), 
        .Y(n4079) );
  OAI2BB2XL U3800 ( .B0(n6729), .B1(n411), .A0N(\ram[218][10] ), .A1N(n6392), 
        .Y(n4080) );
  OAI2BB2XL U3801 ( .B0(n6706), .B1(n411), .A0N(\ram[218][11] ), .A1N(n6392), 
        .Y(n4081) );
  OAI2BB2XL U3802 ( .B0(n6683), .B1(n411), .A0N(\ram[218][12] ), .A1N(n6392), 
        .Y(n4082) );
  OAI2BB2XL U3803 ( .B0(n6660), .B1(n411), .A0N(\ram[218][13] ), .A1N(n6392), 
        .Y(n4083) );
  OAI2BB2XL U3804 ( .B0(n6637), .B1(n411), .A0N(\ram[218][14] ), .A1N(n6392), 
        .Y(n4084) );
  OAI2BB2XL U3805 ( .B0(n6614), .B1(n411), .A0N(\ram[218][15] ), .A1N(n6392), 
        .Y(n4085) );
  OAI2BB2XL U3806 ( .B0(n6962), .B1(n413), .A0N(\ram[219][0] ), .A1N(n6391), 
        .Y(n4086) );
  OAI2BB2XL U3807 ( .B0(n6939), .B1(n413), .A0N(\ram[219][1] ), .A1N(n6391), 
        .Y(n4087) );
  OAI2BB2XL U3808 ( .B0(n6916), .B1(n413), .A0N(\ram[219][2] ), .A1N(n6391), 
        .Y(n4088) );
  OAI2BB2XL U3809 ( .B0(n6893), .B1(n413), .A0N(\ram[219][3] ), .A1N(n6391), 
        .Y(n4089) );
  OAI2BB2XL U3810 ( .B0(n6869), .B1(n413), .A0N(\ram[219][4] ), .A1N(n6391), 
        .Y(n4090) );
  OAI2BB2XL U3811 ( .B0(n6846), .B1(n413), .A0N(\ram[219][5] ), .A1N(n6391), 
        .Y(n4091) );
  OAI2BB2XL U3812 ( .B0(n6823), .B1(n413), .A0N(\ram[219][6] ), .A1N(n6391), 
        .Y(n4092) );
  OAI2BB2XL U3813 ( .B0(n6800), .B1(n413), .A0N(\ram[219][7] ), .A1N(n6391), 
        .Y(n4093) );
  OAI2BB2XL U3814 ( .B0(n6777), .B1(n413), .A0N(\ram[219][8] ), .A1N(n6391), 
        .Y(n4094) );
  OAI2BB2XL U3815 ( .B0(n6754), .B1(n413), .A0N(\ram[219][9] ), .A1N(n6391), 
        .Y(n4095) );
  OAI2BB2XL U3816 ( .B0(n6731), .B1(n413), .A0N(\ram[219][10] ), .A1N(n6391), 
        .Y(n4096) );
  OAI2BB2XL U3817 ( .B0(n6708), .B1(n413), .A0N(\ram[219][11] ), .A1N(n6391), 
        .Y(n4097) );
  OAI2BB2XL U3818 ( .B0(n6685), .B1(n413), .A0N(\ram[219][12] ), .A1N(n6391), 
        .Y(n4098) );
  OAI2BB2XL U3819 ( .B0(n6662), .B1(n413), .A0N(\ram[219][13] ), .A1N(n6391), 
        .Y(n4099) );
  OAI2BB2XL U3820 ( .B0(n6639), .B1(n413), .A0N(\ram[219][14] ), .A1N(n6391), 
        .Y(n4100) );
  OAI2BB2XL U3821 ( .B0(n6616), .B1(n413), .A0N(\ram[219][15] ), .A1N(n6391), 
        .Y(n4101) );
  OAI2BB2XL U3822 ( .B0(n6961), .B1(n415), .A0N(\ram[220][0] ), .A1N(n6390), 
        .Y(n4102) );
  OAI2BB2XL U3823 ( .B0(n6938), .B1(n415), .A0N(\ram[220][1] ), .A1N(n6390), 
        .Y(n4103) );
  OAI2BB2XL U3824 ( .B0(n6915), .B1(n415), .A0N(\ram[220][2] ), .A1N(n6390), 
        .Y(n4104) );
  OAI2BB2XL U3825 ( .B0(n6892), .B1(n415), .A0N(\ram[220][3] ), .A1N(n6390), 
        .Y(n4105) );
  OAI2BB2XL U3826 ( .B0(n6866), .B1(n415), .A0N(\ram[220][4] ), .A1N(n6390), 
        .Y(n4106) );
  OAI2BB2XL U3827 ( .B0(n6843), .B1(n415), .A0N(\ram[220][5] ), .A1N(n6390), 
        .Y(n4107) );
  OAI2BB2XL U3828 ( .B0(n6820), .B1(n415), .A0N(\ram[220][6] ), .A1N(n6390), 
        .Y(n4108) );
  OAI2BB2XL U3829 ( .B0(n6797), .B1(n415), .A0N(\ram[220][7] ), .A1N(n6390), 
        .Y(n4109) );
  OAI2BB2XL U3830 ( .B0(n6774), .B1(n415), .A0N(\ram[220][8] ), .A1N(n6390), 
        .Y(n4110) );
  OAI2BB2XL U3831 ( .B0(n6751), .B1(n415), .A0N(\ram[220][9] ), .A1N(n6390), 
        .Y(n4111) );
  OAI2BB2XL U3832 ( .B0(n6728), .B1(n415), .A0N(\ram[220][10] ), .A1N(n6390), 
        .Y(n4112) );
  OAI2BB2XL U3833 ( .B0(n6705), .B1(n415), .A0N(\ram[220][11] ), .A1N(n6390), 
        .Y(n4113) );
  OAI2BB2XL U3834 ( .B0(n6682), .B1(n415), .A0N(\ram[220][12] ), .A1N(n6390), 
        .Y(n4114) );
  OAI2BB2XL U3835 ( .B0(n6659), .B1(n415), .A0N(\ram[220][13] ), .A1N(n6390), 
        .Y(n4115) );
  OAI2BB2XL U3836 ( .B0(n6636), .B1(n415), .A0N(\ram[220][14] ), .A1N(n6390), 
        .Y(n4116) );
  OAI2BB2XL U3837 ( .B0(n6613), .B1(n415), .A0N(\ram[220][15] ), .A1N(n6390), 
        .Y(n4117) );
  OAI2BB2XL U3838 ( .B0(n6961), .B1(n417), .A0N(\ram[221][0] ), .A1N(n6389), 
        .Y(n4118) );
  OAI2BB2XL U3839 ( .B0(n6938), .B1(n417), .A0N(\ram[221][1] ), .A1N(n6389), 
        .Y(n4119) );
  OAI2BB2XL U3840 ( .B0(n6915), .B1(n417), .A0N(\ram[221][2] ), .A1N(n6389), 
        .Y(n4120) );
  OAI2BB2XL U3841 ( .B0(n6892), .B1(n417), .A0N(\ram[221][3] ), .A1N(n6389), 
        .Y(n4121) );
  OAI2BB2XL U3842 ( .B0(n6866), .B1(n417), .A0N(\ram[221][4] ), .A1N(n6389), 
        .Y(n4122) );
  OAI2BB2XL U3843 ( .B0(n6843), .B1(n417), .A0N(\ram[221][5] ), .A1N(n6389), 
        .Y(n4123) );
  OAI2BB2XL U3844 ( .B0(n6820), .B1(n417), .A0N(\ram[221][6] ), .A1N(n6389), 
        .Y(n4124) );
  OAI2BB2XL U3845 ( .B0(n6797), .B1(n417), .A0N(\ram[221][7] ), .A1N(n6389), 
        .Y(n4125) );
  OAI2BB2XL U3846 ( .B0(n6774), .B1(n417), .A0N(\ram[221][8] ), .A1N(n6389), 
        .Y(n4126) );
  OAI2BB2XL U3847 ( .B0(n6751), .B1(n417), .A0N(\ram[221][9] ), .A1N(n6389), 
        .Y(n4127) );
  OAI2BB2XL U3848 ( .B0(n6728), .B1(n417), .A0N(\ram[221][10] ), .A1N(n6389), 
        .Y(n4128) );
  OAI2BB2XL U3849 ( .B0(n6705), .B1(n417), .A0N(\ram[221][11] ), .A1N(n6389), 
        .Y(n4129) );
  OAI2BB2XL U3850 ( .B0(n6682), .B1(n417), .A0N(\ram[221][12] ), .A1N(n6389), 
        .Y(n4130) );
  OAI2BB2XL U3851 ( .B0(n6659), .B1(n417), .A0N(\ram[221][13] ), .A1N(n6389), 
        .Y(n4131) );
  OAI2BB2XL U3852 ( .B0(n6636), .B1(n417), .A0N(\ram[221][14] ), .A1N(n6389), 
        .Y(n4132) );
  OAI2BB2XL U3853 ( .B0(n6613), .B1(n417), .A0N(\ram[221][15] ), .A1N(n6389), 
        .Y(n4133) );
  OAI2BB2XL U3854 ( .B0(n6961), .B1(n22), .A0N(\ram[222][0] ), .A1N(n6388), 
        .Y(n4134) );
  OAI2BB2XL U3855 ( .B0(n6938), .B1(n22), .A0N(\ram[222][1] ), .A1N(n6388), 
        .Y(n4135) );
  OAI2BB2XL U3856 ( .B0(n6915), .B1(n22), .A0N(\ram[222][2] ), .A1N(n6388), 
        .Y(n4136) );
  OAI2BB2XL U3857 ( .B0(n6892), .B1(n22), .A0N(\ram[222][3] ), .A1N(n6388), 
        .Y(n4137) );
  OAI2BB2XL U3858 ( .B0(n6866), .B1(n22), .A0N(\ram[222][4] ), .A1N(n6388), 
        .Y(n4138) );
  OAI2BB2XL U3859 ( .B0(n6843), .B1(n22), .A0N(\ram[222][5] ), .A1N(n6388), 
        .Y(n4139) );
  OAI2BB2XL U3860 ( .B0(n6820), .B1(n22), .A0N(\ram[222][6] ), .A1N(n6388), 
        .Y(n4140) );
  OAI2BB2XL U3861 ( .B0(n6797), .B1(n22), .A0N(\ram[222][7] ), .A1N(n6388), 
        .Y(n4141) );
  OAI2BB2XL U3862 ( .B0(n6774), .B1(n22), .A0N(\ram[222][8] ), .A1N(n6388), 
        .Y(n4142) );
  OAI2BB2XL U3863 ( .B0(n6751), .B1(n22), .A0N(\ram[222][9] ), .A1N(n6388), 
        .Y(n4143) );
  OAI2BB2XL U3864 ( .B0(n6728), .B1(n22), .A0N(\ram[222][10] ), .A1N(n6388), 
        .Y(n4144) );
  OAI2BB2XL U3865 ( .B0(n6705), .B1(n22), .A0N(\ram[222][11] ), .A1N(n6388), 
        .Y(n4145) );
  OAI2BB2XL U3866 ( .B0(n6682), .B1(n22), .A0N(\ram[222][12] ), .A1N(n6388), 
        .Y(n4146) );
  OAI2BB2XL U3867 ( .B0(n6659), .B1(n22), .A0N(\ram[222][13] ), .A1N(n6388), 
        .Y(n4147) );
  OAI2BB2XL U3868 ( .B0(n6636), .B1(n22), .A0N(\ram[222][14] ), .A1N(n6388), 
        .Y(n4148) );
  OAI2BB2XL U3869 ( .B0(n6613), .B1(n22), .A0N(\ram[222][15] ), .A1N(n6388), 
        .Y(n4149) );
  OAI2BB2XL U3870 ( .B0(n6961), .B1(n23), .A0N(\ram[223][0] ), .A1N(n6387), 
        .Y(n4150) );
  OAI2BB2XL U3871 ( .B0(n6938), .B1(n23), .A0N(\ram[223][1] ), .A1N(n6387), 
        .Y(n4151) );
  OAI2BB2XL U3872 ( .B0(n6915), .B1(n23), .A0N(\ram[223][2] ), .A1N(n6387), 
        .Y(n4152) );
  OAI2BB2XL U3873 ( .B0(n6892), .B1(n23), .A0N(\ram[223][3] ), .A1N(n6387), 
        .Y(n4153) );
  OAI2BB2XL U3874 ( .B0(n6866), .B1(n23), .A0N(\ram[223][4] ), .A1N(n6387), 
        .Y(n4154) );
  OAI2BB2XL U3875 ( .B0(n6843), .B1(n23), .A0N(\ram[223][5] ), .A1N(n6387), 
        .Y(n4155) );
  OAI2BB2XL U3876 ( .B0(n6820), .B1(n23), .A0N(\ram[223][6] ), .A1N(n6387), 
        .Y(n4156) );
  OAI2BB2XL U3877 ( .B0(n6797), .B1(n23), .A0N(\ram[223][7] ), .A1N(n6387), 
        .Y(n4157) );
  OAI2BB2XL U3878 ( .B0(n6774), .B1(n23), .A0N(\ram[223][8] ), .A1N(n6387), 
        .Y(n4158) );
  OAI2BB2XL U3879 ( .B0(n6751), .B1(n23), .A0N(\ram[223][9] ), .A1N(n6387), 
        .Y(n4159) );
  OAI2BB2XL U3880 ( .B0(n6728), .B1(n23), .A0N(\ram[223][10] ), .A1N(n6387), 
        .Y(n4160) );
  OAI2BB2XL U3881 ( .B0(n6705), .B1(n23), .A0N(\ram[223][11] ), .A1N(n6387), 
        .Y(n4161) );
  OAI2BB2XL U3882 ( .B0(n6682), .B1(n23), .A0N(\ram[223][12] ), .A1N(n6387), 
        .Y(n4162) );
  OAI2BB2XL U3883 ( .B0(n6659), .B1(n23), .A0N(\ram[223][13] ), .A1N(n6387), 
        .Y(n4163) );
  OAI2BB2XL U3884 ( .B0(n6636), .B1(n23), .A0N(\ram[223][14] ), .A1N(n6387), 
        .Y(n4164) );
  OAI2BB2XL U3885 ( .B0(n6613), .B1(n23), .A0N(\ram[223][15] ), .A1N(n6387), 
        .Y(n4165) );
  OAI2BB2XL U3886 ( .B0(n6961), .B1(n24), .A0N(\ram[224][0] ), .A1N(n6386), 
        .Y(n4166) );
  OAI2BB2XL U3887 ( .B0(n6938), .B1(n24), .A0N(\ram[224][1] ), .A1N(n6386), 
        .Y(n4167) );
  OAI2BB2XL U3888 ( .B0(n6915), .B1(n24), .A0N(\ram[224][2] ), .A1N(n6386), 
        .Y(n4168) );
  OAI2BB2XL U3889 ( .B0(n6892), .B1(n24), .A0N(\ram[224][3] ), .A1N(n6386), 
        .Y(n4169) );
  OAI2BB2XL U3890 ( .B0(n6866), .B1(n24), .A0N(\ram[224][4] ), .A1N(n6386), 
        .Y(n4170) );
  OAI2BB2XL U3891 ( .B0(n6843), .B1(n24), .A0N(\ram[224][5] ), .A1N(n6386), 
        .Y(n4171) );
  OAI2BB2XL U3892 ( .B0(n6820), .B1(n24), .A0N(\ram[224][6] ), .A1N(n6386), 
        .Y(n4172) );
  OAI2BB2XL U3893 ( .B0(n6797), .B1(n24), .A0N(\ram[224][7] ), .A1N(n6386), 
        .Y(n4173) );
  OAI2BB2XL U3894 ( .B0(n6774), .B1(n24), .A0N(\ram[224][8] ), .A1N(n6386), 
        .Y(n4174) );
  OAI2BB2XL U3895 ( .B0(n6751), .B1(n24), .A0N(\ram[224][9] ), .A1N(n6386), 
        .Y(n4175) );
  OAI2BB2XL U3896 ( .B0(n6728), .B1(n24), .A0N(\ram[224][10] ), .A1N(n6386), 
        .Y(n4176) );
  OAI2BB2XL U3897 ( .B0(n6705), .B1(n24), .A0N(\ram[224][11] ), .A1N(n6386), 
        .Y(n4177) );
  OAI2BB2XL U3898 ( .B0(n6682), .B1(n24), .A0N(\ram[224][12] ), .A1N(n6386), 
        .Y(n4178) );
  OAI2BB2XL U3899 ( .B0(n6659), .B1(n24), .A0N(\ram[224][13] ), .A1N(n6386), 
        .Y(n4179) );
  OAI2BB2XL U3900 ( .B0(n6636), .B1(n24), .A0N(\ram[224][14] ), .A1N(n6386), 
        .Y(n4180) );
  OAI2BB2XL U3901 ( .B0(n6613), .B1(n24), .A0N(\ram[224][15] ), .A1N(n6386), 
        .Y(n4181) );
  OAI2BB2XL U3902 ( .B0(n6961), .B1(n25), .A0N(\ram[225][0] ), .A1N(n6385), 
        .Y(n4182) );
  OAI2BB2XL U3903 ( .B0(n6938), .B1(n25), .A0N(\ram[225][1] ), .A1N(n6385), 
        .Y(n4183) );
  OAI2BB2XL U3904 ( .B0(n6915), .B1(n25), .A0N(\ram[225][2] ), .A1N(n6385), 
        .Y(n4184) );
  OAI2BB2XL U3905 ( .B0(n6892), .B1(n25), .A0N(\ram[225][3] ), .A1N(n6385), 
        .Y(n4185) );
  OAI2BB2XL U3906 ( .B0(n6866), .B1(n25), .A0N(\ram[225][4] ), .A1N(n6385), 
        .Y(n4186) );
  OAI2BB2XL U3907 ( .B0(n6843), .B1(n25), .A0N(\ram[225][5] ), .A1N(n6385), 
        .Y(n4187) );
  OAI2BB2XL U3908 ( .B0(n6820), .B1(n25), .A0N(\ram[225][6] ), .A1N(n6385), 
        .Y(n4188) );
  OAI2BB2XL U3909 ( .B0(n6797), .B1(n25), .A0N(\ram[225][7] ), .A1N(n6385), 
        .Y(n4189) );
  OAI2BB2XL U3910 ( .B0(n6774), .B1(n25), .A0N(\ram[225][8] ), .A1N(n6385), 
        .Y(n4190) );
  OAI2BB2XL U3911 ( .B0(n6751), .B1(n25), .A0N(\ram[225][9] ), .A1N(n6385), 
        .Y(n4191) );
  OAI2BB2XL U3912 ( .B0(n6728), .B1(n25), .A0N(\ram[225][10] ), .A1N(n6385), 
        .Y(n4192) );
  OAI2BB2XL U3913 ( .B0(n6705), .B1(n25), .A0N(\ram[225][11] ), .A1N(n6385), 
        .Y(n4193) );
  OAI2BB2XL U3914 ( .B0(n6682), .B1(n25), .A0N(\ram[225][12] ), .A1N(n6385), 
        .Y(n4194) );
  OAI2BB2XL U3915 ( .B0(n6659), .B1(n25), .A0N(\ram[225][13] ), .A1N(n6385), 
        .Y(n4195) );
  OAI2BB2XL U3916 ( .B0(n6636), .B1(n25), .A0N(\ram[225][14] ), .A1N(n6385), 
        .Y(n4196) );
  OAI2BB2XL U3917 ( .B0(n6613), .B1(n25), .A0N(\ram[225][15] ), .A1N(n6385), 
        .Y(n4197) );
  OAI2BB2XL U3918 ( .B0(n6961), .B1(n26), .A0N(\ram[226][0] ), .A1N(n6384), 
        .Y(n4198) );
  OAI2BB2XL U3919 ( .B0(n6938), .B1(n26), .A0N(\ram[226][1] ), .A1N(n6384), 
        .Y(n4199) );
  OAI2BB2XL U3920 ( .B0(n6915), .B1(n26), .A0N(\ram[226][2] ), .A1N(n6384), 
        .Y(n4200) );
  OAI2BB2XL U3921 ( .B0(n6892), .B1(n26), .A0N(\ram[226][3] ), .A1N(n6384), 
        .Y(n4201) );
  OAI2BB2XL U3922 ( .B0(n6866), .B1(n26), .A0N(\ram[226][4] ), .A1N(n6384), 
        .Y(n4202) );
  OAI2BB2XL U3923 ( .B0(n6843), .B1(n26), .A0N(\ram[226][5] ), .A1N(n6384), 
        .Y(n4203) );
  OAI2BB2XL U3924 ( .B0(n6820), .B1(n26), .A0N(\ram[226][6] ), .A1N(n6384), 
        .Y(n4204) );
  OAI2BB2XL U3925 ( .B0(n6797), .B1(n26), .A0N(\ram[226][7] ), .A1N(n6384), 
        .Y(n4205) );
  OAI2BB2XL U3926 ( .B0(n6774), .B1(n26), .A0N(\ram[226][8] ), .A1N(n6384), 
        .Y(n4206) );
  OAI2BB2XL U3927 ( .B0(n6751), .B1(n26), .A0N(\ram[226][9] ), .A1N(n6384), 
        .Y(n4207) );
  OAI2BB2XL U3928 ( .B0(n6728), .B1(n26), .A0N(\ram[226][10] ), .A1N(n6384), 
        .Y(n4208) );
  OAI2BB2XL U3929 ( .B0(n6705), .B1(n26), .A0N(\ram[226][11] ), .A1N(n6384), 
        .Y(n4209) );
  OAI2BB2XL U3930 ( .B0(n6682), .B1(n26), .A0N(\ram[226][12] ), .A1N(n6384), 
        .Y(n4210) );
  OAI2BB2XL U3931 ( .B0(n6659), .B1(n26), .A0N(\ram[226][13] ), .A1N(n6384), 
        .Y(n4211) );
  OAI2BB2XL U3932 ( .B0(n6636), .B1(n26), .A0N(\ram[226][14] ), .A1N(n6384), 
        .Y(n4212) );
  OAI2BB2XL U3933 ( .B0(n6613), .B1(n26), .A0N(\ram[226][15] ), .A1N(n6384), 
        .Y(n4213) );
  OAI2BB2XL U3934 ( .B0(n6961), .B1(n28), .A0N(\ram[227][0] ), .A1N(n6383), 
        .Y(n4214) );
  OAI2BB2XL U3935 ( .B0(n6938), .B1(n28), .A0N(\ram[227][1] ), .A1N(n6383), 
        .Y(n4215) );
  OAI2BB2XL U3936 ( .B0(n6915), .B1(n28), .A0N(\ram[227][2] ), .A1N(n6383), 
        .Y(n4216) );
  OAI2BB2XL U3937 ( .B0(n6892), .B1(n28), .A0N(\ram[227][3] ), .A1N(n6383), 
        .Y(n4217) );
  OAI2BB2XL U3938 ( .B0(n6866), .B1(n28), .A0N(\ram[227][4] ), .A1N(n6383), 
        .Y(n4218) );
  OAI2BB2XL U3939 ( .B0(n6843), .B1(n28), .A0N(\ram[227][5] ), .A1N(n6383), 
        .Y(n4219) );
  OAI2BB2XL U3940 ( .B0(n6820), .B1(n28), .A0N(\ram[227][6] ), .A1N(n6383), 
        .Y(n4220) );
  OAI2BB2XL U3941 ( .B0(n6797), .B1(n28), .A0N(\ram[227][7] ), .A1N(n6383), 
        .Y(n4221) );
  OAI2BB2XL U3942 ( .B0(n6774), .B1(n28), .A0N(\ram[227][8] ), .A1N(n6383), 
        .Y(n4222) );
  OAI2BB2XL U3943 ( .B0(n6751), .B1(n28), .A0N(\ram[227][9] ), .A1N(n6383), 
        .Y(n4223) );
  OAI2BB2XL U3944 ( .B0(n6728), .B1(n28), .A0N(\ram[227][10] ), .A1N(n6383), 
        .Y(n4224) );
  OAI2BB2XL U3945 ( .B0(n6705), .B1(n28), .A0N(\ram[227][11] ), .A1N(n6383), 
        .Y(n4225) );
  OAI2BB2XL U3946 ( .B0(n6682), .B1(n28), .A0N(\ram[227][12] ), .A1N(n6383), 
        .Y(n4226) );
  OAI2BB2XL U3947 ( .B0(n6659), .B1(n28), .A0N(\ram[227][13] ), .A1N(n6383), 
        .Y(n4227) );
  OAI2BB2XL U3948 ( .B0(n6636), .B1(n28), .A0N(\ram[227][14] ), .A1N(n6383), 
        .Y(n4228) );
  OAI2BB2XL U3949 ( .B0(n6613), .B1(n28), .A0N(\ram[227][15] ), .A1N(n6383), 
        .Y(n4229) );
  OAI2BB2XL U3950 ( .B0(n6961), .B1(n29), .A0N(\ram[228][0] ), .A1N(n6382), 
        .Y(n4230) );
  OAI2BB2XL U3951 ( .B0(n6938), .B1(n29), .A0N(\ram[228][1] ), .A1N(n6382), 
        .Y(n4231) );
  OAI2BB2XL U3952 ( .B0(n6915), .B1(n29), .A0N(\ram[228][2] ), .A1N(n6382), 
        .Y(n4232) );
  OAI2BB2XL U3953 ( .B0(n6892), .B1(n29), .A0N(\ram[228][3] ), .A1N(n6382), 
        .Y(n4233) );
  OAI2BB2XL U3954 ( .B0(n6866), .B1(n29), .A0N(\ram[228][4] ), .A1N(n6382), 
        .Y(n4234) );
  OAI2BB2XL U3955 ( .B0(n6843), .B1(n29), .A0N(\ram[228][5] ), .A1N(n6382), 
        .Y(n4235) );
  OAI2BB2XL U3956 ( .B0(n6820), .B1(n29), .A0N(\ram[228][6] ), .A1N(n6382), 
        .Y(n4236) );
  OAI2BB2XL U3957 ( .B0(n6797), .B1(n29), .A0N(\ram[228][7] ), .A1N(n6382), 
        .Y(n4237) );
  OAI2BB2XL U3958 ( .B0(n6774), .B1(n29), .A0N(\ram[228][8] ), .A1N(n6382), 
        .Y(n4238) );
  OAI2BB2XL U3959 ( .B0(n6751), .B1(n29), .A0N(\ram[228][9] ), .A1N(n6382), 
        .Y(n4239) );
  OAI2BB2XL U3960 ( .B0(n6728), .B1(n29), .A0N(\ram[228][10] ), .A1N(n6382), 
        .Y(n4240) );
  OAI2BB2XL U3961 ( .B0(n6705), .B1(n29), .A0N(\ram[228][11] ), .A1N(n6382), 
        .Y(n4241) );
  OAI2BB2XL U3962 ( .B0(n6682), .B1(n29), .A0N(\ram[228][12] ), .A1N(n6382), 
        .Y(n4242) );
  OAI2BB2XL U3963 ( .B0(n6659), .B1(n29), .A0N(\ram[228][13] ), .A1N(n6382), 
        .Y(n4243) );
  OAI2BB2XL U3964 ( .B0(n6636), .B1(n29), .A0N(\ram[228][14] ), .A1N(n6382), 
        .Y(n4244) );
  OAI2BB2XL U3965 ( .B0(n6613), .B1(n29), .A0N(\ram[228][15] ), .A1N(n6382), 
        .Y(n4245) );
  OAI2BB2XL U3966 ( .B0(n6961), .B1(n31), .A0N(\ram[229][0] ), .A1N(n6381), 
        .Y(n4246) );
  OAI2BB2XL U3967 ( .B0(n6938), .B1(n31), .A0N(\ram[229][1] ), .A1N(n6381), 
        .Y(n4247) );
  OAI2BB2XL U3968 ( .B0(n6915), .B1(n31), .A0N(\ram[229][2] ), .A1N(n6381), 
        .Y(n4248) );
  OAI2BB2XL U3969 ( .B0(n6892), .B1(n31), .A0N(\ram[229][3] ), .A1N(n6381), 
        .Y(n4249) );
  OAI2BB2XL U3970 ( .B0(n6866), .B1(n31), .A0N(\ram[229][4] ), .A1N(n6381), 
        .Y(n4250) );
  OAI2BB2XL U3971 ( .B0(n6843), .B1(n31), .A0N(\ram[229][5] ), .A1N(n6381), 
        .Y(n4251) );
  OAI2BB2XL U3972 ( .B0(n6820), .B1(n31), .A0N(\ram[229][6] ), .A1N(n6381), 
        .Y(n4252) );
  OAI2BB2XL U3973 ( .B0(n6797), .B1(n31), .A0N(\ram[229][7] ), .A1N(n6381), 
        .Y(n4253) );
  OAI2BB2XL U3974 ( .B0(n6774), .B1(n31), .A0N(\ram[229][8] ), .A1N(n6381), 
        .Y(n4254) );
  OAI2BB2XL U3975 ( .B0(n6751), .B1(n31), .A0N(\ram[229][9] ), .A1N(n6381), 
        .Y(n4255) );
  OAI2BB2XL U3976 ( .B0(n6728), .B1(n31), .A0N(\ram[229][10] ), .A1N(n6381), 
        .Y(n4256) );
  OAI2BB2XL U3977 ( .B0(n6705), .B1(n31), .A0N(\ram[229][11] ), .A1N(n6381), 
        .Y(n4257) );
  OAI2BB2XL U3978 ( .B0(n6682), .B1(n31), .A0N(\ram[229][12] ), .A1N(n6381), 
        .Y(n4258) );
  OAI2BB2XL U3979 ( .B0(n6659), .B1(n31), .A0N(\ram[229][13] ), .A1N(n6381), 
        .Y(n4259) );
  OAI2BB2XL U3980 ( .B0(n6636), .B1(n31), .A0N(\ram[229][14] ), .A1N(n6381), 
        .Y(n4260) );
  OAI2BB2XL U3981 ( .B0(n6613), .B1(n31), .A0N(\ram[229][15] ), .A1N(n6381), 
        .Y(n4261) );
  OAI2BB2XL U3982 ( .B0(n6961), .B1(n32), .A0N(\ram[230][0] ), .A1N(n6380), 
        .Y(n4262) );
  OAI2BB2XL U3983 ( .B0(n6938), .B1(n32), .A0N(\ram[230][1] ), .A1N(n6380), 
        .Y(n4263) );
  OAI2BB2XL U3984 ( .B0(n6915), .B1(n32), .A0N(\ram[230][2] ), .A1N(n6380), 
        .Y(n4264) );
  OAI2BB2XL U3985 ( .B0(n6892), .B1(n32), .A0N(\ram[230][3] ), .A1N(n6380), 
        .Y(n4265) );
  OAI2BB2XL U3986 ( .B0(n6866), .B1(n32), .A0N(\ram[230][4] ), .A1N(n6380), 
        .Y(n4266) );
  OAI2BB2XL U3987 ( .B0(n6843), .B1(n32), .A0N(\ram[230][5] ), .A1N(n6380), 
        .Y(n4267) );
  OAI2BB2XL U3988 ( .B0(n6820), .B1(n32), .A0N(\ram[230][6] ), .A1N(n6380), 
        .Y(n4268) );
  OAI2BB2XL U3989 ( .B0(n6797), .B1(n32), .A0N(\ram[230][7] ), .A1N(n6380), 
        .Y(n4269) );
  OAI2BB2XL U3990 ( .B0(n6774), .B1(n32), .A0N(\ram[230][8] ), .A1N(n6380), 
        .Y(n4270) );
  OAI2BB2XL U3991 ( .B0(n6751), .B1(n32), .A0N(\ram[230][9] ), .A1N(n6380), 
        .Y(n4271) );
  OAI2BB2XL U3992 ( .B0(n6728), .B1(n32), .A0N(\ram[230][10] ), .A1N(n6380), 
        .Y(n4272) );
  OAI2BB2XL U3993 ( .B0(n6705), .B1(n32), .A0N(\ram[230][11] ), .A1N(n6380), 
        .Y(n4273) );
  OAI2BB2XL U3994 ( .B0(n6682), .B1(n32), .A0N(\ram[230][12] ), .A1N(n6380), 
        .Y(n4274) );
  OAI2BB2XL U3995 ( .B0(n6659), .B1(n32), .A0N(\ram[230][13] ), .A1N(n6380), 
        .Y(n4275) );
  OAI2BB2XL U3996 ( .B0(n6636), .B1(n32), .A0N(\ram[230][14] ), .A1N(n6380), 
        .Y(n4276) );
  OAI2BB2XL U3997 ( .B0(n6613), .B1(n32), .A0N(\ram[230][15] ), .A1N(n6380), 
        .Y(n4277) );
  OAI2BB2XL U3998 ( .B0(n6961), .B1(n34), .A0N(\ram[231][0] ), .A1N(n6379), 
        .Y(n4278) );
  OAI2BB2XL U3999 ( .B0(n6938), .B1(n34), .A0N(\ram[231][1] ), .A1N(n6379), 
        .Y(n4279) );
  OAI2BB2XL U4000 ( .B0(n6915), .B1(n34), .A0N(\ram[231][2] ), .A1N(n6379), 
        .Y(n4280) );
  OAI2BB2XL U4001 ( .B0(n6892), .B1(n34), .A0N(\ram[231][3] ), .A1N(n6379), 
        .Y(n4281) );
  OAI2BB2XL U4002 ( .B0(n6866), .B1(n34), .A0N(\ram[231][4] ), .A1N(n6379), 
        .Y(n4282) );
  OAI2BB2XL U4003 ( .B0(n6843), .B1(n34), .A0N(\ram[231][5] ), .A1N(n6379), 
        .Y(n4283) );
  OAI2BB2XL U4004 ( .B0(n6820), .B1(n34), .A0N(\ram[231][6] ), .A1N(n6379), 
        .Y(n4284) );
  OAI2BB2XL U4005 ( .B0(n6797), .B1(n34), .A0N(\ram[231][7] ), .A1N(n6379), 
        .Y(n4285) );
  OAI2BB2XL U4006 ( .B0(n6774), .B1(n34), .A0N(\ram[231][8] ), .A1N(n6379), 
        .Y(n4286) );
  OAI2BB2XL U4007 ( .B0(n6751), .B1(n34), .A0N(\ram[231][9] ), .A1N(n6379), 
        .Y(n4287) );
  OAI2BB2XL U4008 ( .B0(n6728), .B1(n34), .A0N(\ram[231][10] ), .A1N(n6379), 
        .Y(n4288) );
  OAI2BB2XL U4009 ( .B0(n6705), .B1(n34), .A0N(\ram[231][11] ), .A1N(n6379), 
        .Y(n4289) );
  OAI2BB2XL U4010 ( .B0(n6682), .B1(n34), .A0N(\ram[231][12] ), .A1N(n6379), 
        .Y(n4290) );
  OAI2BB2XL U4011 ( .B0(n6659), .B1(n34), .A0N(\ram[231][13] ), .A1N(n6379), 
        .Y(n4291) );
  OAI2BB2XL U4012 ( .B0(n6636), .B1(n34), .A0N(\ram[231][14] ), .A1N(n6379), 
        .Y(n4292) );
  OAI2BB2XL U4013 ( .B0(n6613), .B1(n34), .A0N(\ram[231][15] ), .A1N(n6379), 
        .Y(n4293) );
  OAI2BB2XL U4014 ( .B0(n6960), .B1(n35), .A0N(\ram[232][0] ), .A1N(n6378), 
        .Y(n4294) );
  OAI2BB2XL U4015 ( .B0(n6937), .B1(n35), .A0N(\ram[232][1] ), .A1N(n6378), 
        .Y(n4295) );
  OAI2BB2XL U4016 ( .B0(n6914), .B1(n35), .A0N(\ram[232][2] ), .A1N(n6378), 
        .Y(n4296) );
  OAI2BB2XL U4017 ( .B0(n6891), .B1(n35), .A0N(\ram[232][3] ), .A1N(n6378), 
        .Y(n4297) );
  OAI2BB2XL U4018 ( .B0(n6865), .B1(n35), .A0N(\ram[232][4] ), .A1N(n6378), 
        .Y(n4298) );
  OAI2BB2XL U4019 ( .B0(n6842), .B1(n35), .A0N(\ram[232][5] ), .A1N(n6378), 
        .Y(n4299) );
  OAI2BB2XL U4020 ( .B0(n6819), .B1(n35), .A0N(\ram[232][6] ), .A1N(n6378), 
        .Y(n4300) );
  OAI2BB2XL U4021 ( .B0(n6796), .B1(n35), .A0N(\ram[232][7] ), .A1N(n6378), 
        .Y(n4301) );
  OAI2BB2XL U4022 ( .B0(n6773), .B1(n35), .A0N(\ram[232][8] ), .A1N(n6378), 
        .Y(n4302) );
  OAI2BB2XL U4023 ( .B0(n6750), .B1(n35), .A0N(\ram[232][9] ), .A1N(n6378), 
        .Y(n4303) );
  OAI2BB2XL U4024 ( .B0(n6727), .B1(n35), .A0N(\ram[232][10] ), .A1N(n6378), 
        .Y(n4304) );
  OAI2BB2XL U4025 ( .B0(n6704), .B1(n35), .A0N(\ram[232][11] ), .A1N(n6378), 
        .Y(n4305) );
  OAI2BB2XL U4026 ( .B0(n6681), .B1(n35), .A0N(\ram[232][12] ), .A1N(n6378), 
        .Y(n4306) );
  OAI2BB2XL U4027 ( .B0(n6658), .B1(n35), .A0N(\ram[232][13] ), .A1N(n6378), 
        .Y(n4307) );
  OAI2BB2XL U4028 ( .B0(n6635), .B1(n35), .A0N(\ram[232][14] ), .A1N(n6378), 
        .Y(n4308) );
  OAI2BB2XL U4029 ( .B0(n6612), .B1(n35), .A0N(\ram[232][15] ), .A1N(n6378), 
        .Y(n4309) );
  OAI2BB2XL U4030 ( .B0(n6960), .B1(n37), .A0N(\ram[233][0] ), .A1N(n6377), 
        .Y(n4310) );
  OAI2BB2XL U4031 ( .B0(n6937), .B1(n37), .A0N(\ram[233][1] ), .A1N(n6377), 
        .Y(n4311) );
  OAI2BB2XL U4032 ( .B0(n6914), .B1(n37), .A0N(\ram[233][2] ), .A1N(n6377), 
        .Y(n4312) );
  OAI2BB2XL U4033 ( .B0(n6891), .B1(n37), .A0N(\ram[233][3] ), .A1N(n6377), 
        .Y(n4313) );
  OAI2BB2XL U4034 ( .B0(n6865), .B1(n37), .A0N(\ram[233][4] ), .A1N(n6377), 
        .Y(n4314) );
  OAI2BB2XL U4035 ( .B0(n6842), .B1(n37), .A0N(\ram[233][5] ), .A1N(n6377), 
        .Y(n4315) );
  OAI2BB2XL U4036 ( .B0(n6819), .B1(n37), .A0N(\ram[233][6] ), .A1N(n6377), 
        .Y(n4316) );
  OAI2BB2XL U4037 ( .B0(n6796), .B1(n37), .A0N(\ram[233][7] ), .A1N(n6377), 
        .Y(n4317) );
  OAI2BB2XL U4038 ( .B0(n6773), .B1(n37), .A0N(\ram[233][8] ), .A1N(n6377), 
        .Y(n4318) );
  OAI2BB2XL U4039 ( .B0(n6750), .B1(n37), .A0N(\ram[233][9] ), .A1N(n6377), 
        .Y(n4319) );
  OAI2BB2XL U4040 ( .B0(n6727), .B1(n37), .A0N(\ram[233][10] ), .A1N(n6377), 
        .Y(n4320) );
  OAI2BB2XL U4041 ( .B0(n6704), .B1(n37), .A0N(\ram[233][11] ), .A1N(n6377), 
        .Y(n4321) );
  OAI2BB2XL U4042 ( .B0(n6681), .B1(n37), .A0N(\ram[233][12] ), .A1N(n6377), 
        .Y(n4322) );
  OAI2BB2XL U4043 ( .B0(n6658), .B1(n37), .A0N(\ram[233][13] ), .A1N(n6377), 
        .Y(n4323) );
  OAI2BB2XL U4044 ( .B0(n6635), .B1(n37), .A0N(\ram[233][14] ), .A1N(n6377), 
        .Y(n4324) );
  OAI2BB2XL U4045 ( .B0(n6612), .B1(n37), .A0N(\ram[233][15] ), .A1N(n6377), 
        .Y(n4325) );
  OAI2BB2XL U4046 ( .B0(n6960), .B1(n38), .A0N(\ram[234][0] ), .A1N(n6376), 
        .Y(n4326) );
  OAI2BB2XL U4047 ( .B0(n6937), .B1(n38), .A0N(\ram[234][1] ), .A1N(n6376), 
        .Y(n4327) );
  OAI2BB2XL U4048 ( .B0(n6914), .B1(n38), .A0N(\ram[234][2] ), .A1N(n6376), 
        .Y(n4328) );
  OAI2BB2XL U4049 ( .B0(n6891), .B1(n38), .A0N(\ram[234][3] ), .A1N(n6376), 
        .Y(n4329) );
  OAI2BB2XL U4050 ( .B0(n6865), .B1(n38), .A0N(\ram[234][4] ), .A1N(n6376), 
        .Y(n4330) );
  OAI2BB2XL U4051 ( .B0(n6842), .B1(n38), .A0N(\ram[234][5] ), .A1N(n6376), 
        .Y(n4331) );
  OAI2BB2XL U4052 ( .B0(n6819), .B1(n38), .A0N(\ram[234][6] ), .A1N(n6376), 
        .Y(n4332) );
  OAI2BB2XL U4053 ( .B0(n6796), .B1(n38), .A0N(\ram[234][7] ), .A1N(n6376), 
        .Y(n4333) );
  OAI2BB2XL U4054 ( .B0(n6773), .B1(n38), .A0N(\ram[234][8] ), .A1N(n6376), 
        .Y(n4334) );
  OAI2BB2XL U4055 ( .B0(n6750), .B1(n38), .A0N(\ram[234][9] ), .A1N(n6376), 
        .Y(n4335) );
  OAI2BB2XL U4056 ( .B0(n6727), .B1(n38), .A0N(\ram[234][10] ), .A1N(n6376), 
        .Y(n4336) );
  OAI2BB2XL U4057 ( .B0(n6704), .B1(n38), .A0N(\ram[234][11] ), .A1N(n6376), 
        .Y(n4337) );
  OAI2BB2XL U4058 ( .B0(n6681), .B1(n38), .A0N(\ram[234][12] ), .A1N(n6376), 
        .Y(n4338) );
  OAI2BB2XL U4059 ( .B0(n6658), .B1(n38), .A0N(\ram[234][13] ), .A1N(n6376), 
        .Y(n4339) );
  OAI2BB2XL U4060 ( .B0(n6635), .B1(n38), .A0N(\ram[234][14] ), .A1N(n6376), 
        .Y(n4340) );
  OAI2BB2XL U4061 ( .B0(n6612), .B1(n38), .A0N(\ram[234][15] ), .A1N(n6376), 
        .Y(n4341) );
  OAI2BB2XL U4062 ( .B0(n6960), .B1(n419), .A0N(\ram[235][0] ), .A1N(n6375), 
        .Y(n4342) );
  OAI2BB2XL U4063 ( .B0(n6937), .B1(n419), .A0N(\ram[235][1] ), .A1N(n6375), 
        .Y(n4343) );
  OAI2BB2XL U4064 ( .B0(n6914), .B1(n419), .A0N(\ram[235][2] ), .A1N(n6375), 
        .Y(n4344) );
  OAI2BB2XL U4065 ( .B0(n6891), .B1(n419), .A0N(\ram[235][3] ), .A1N(n6375), 
        .Y(n4345) );
  OAI2BB2XL U4066 ( .B0(n6865), .B1(n419), .A0N(\ram[235][4] ), .A1N(n6375), 
        .Y(n4346) );
  OAI2BB2XL U4067 ( .B0(n6842), .B1(n419), .A0N(\ram[235][5] ), .A1N(n6375), 
        .Y(n4347) );
  OAI2BB2XL U4068 ( .B0(n6819), .B1(n419), .A0N(\ram[235][6] ), .A1N(n6375), 
        .Y(n4348) );
  OAI2BB2XL U4069 ( .B0(n6796), .B1(n419), .A0N(\ram[235][7] ), .A1N(n6375), 
        .Y(n4349) );
  OAI2BB2XL U4070 ( .B0(n6773), .B1(n419), .A0N(\ram[235][8] ), .A1N(n6375), 
        .Y(n4350) );
  OAI2BB2XL U4071 ( .B0(n6750), .B1(n419), .A0N(\ram[235][9] ), .A1N(n6375), 
        .Y(n4351) );
  OAI2BB2XL U4072 ( .B0(n6727), .B1(n419), .A0N(\ram[235][10] ), .A1N(n6375), 
        .Y(n4352) );
  OAI2BB2XL U4073 ( .B0(n6704), .B1(n419), .A0N(\ram[235][11] ), .A1N(n6375), 
        .Y(n4353) );
  OAI2BB2XL U4074 ( .B0(n6681), .B1(n419), .A0N(\ram[235][12] ), .A1N(n6375), 
        .Y(n4354) );
  OAI2BB2XL U4075 ( .B0(n6658), .B1(n419), .A0N(\ram[235][13] ), .A1N(n6375), 
        .Y(n4355) );
  OAI2BB2XL U4076 ( .B0(n6635), .B1(n419), .A0N(\ram[235][14] ), .A1N(n6375), 
        .Y(n4356) );
  OAI2BB2XL U4077 ( .B0(n6612), .B1(n419), .A0N(\ram[235][15] ), .A1N(n6375), 
        .Y(n4357) );
  OAI2BB2XL U4078 ( .B0(n6960), .B1(n421), .A0N(\ram[236][0] ), .A1N(n6374), 
        .Y(n4358) );
  OAI2BB2XL U4079 ( .B0(n6937), .B1(n421), .A0N(\ram[236][1] ), .A1N(n6374), 
        .Y(n4359) );
  OAI2BB2XL U4080 ( .B0(n6914), .B1(n421), .A0N(\ram[236][2] ), .A1N(n6374), 
        .Y(n4360) );
  OAI2BB2XL U4081 ( .B0(n6891), .B1(n421), .A0N(\ram[236][3] ), .A1N(n6374), 
        .Y(n4361) );
  OAI2BB2XL U4082 ( .B0(n6865), .B1(n421), .A0N(\ram[236][4] ), .A1N(n6374), 
        .Y(n4362) );
  OAI2BB2XL U4083 ( .B0(n6842), .B1(n421), .A0N(\ram[236][5] ), .A1N(n6374), 
        .Y(n4363) );
  OAI2BB2XL U4084 ( .B0(n6819), .B1(n421), .A0N(\ram[236][6] ), .A1N(n6374), 
        .Y(n4364) );
  OAI2BB2XL U4085 ( .B0(n6796), .B1(n421), .A0N(\ram[236][7] ), .A1N(n6374), 
        .Y(n4365) );
  OAI2BB2XL U4086 ( .B0(n6773), .B1(n421), .A0N(\ram[236][8] ), .A1N(n6374), 
        .Y(n4366) );
  OAI2BB2XL U4087 ( .B0(n6750), .B1(n421), .A0N(\ram[236][9] ), .A1N(n6374), 
        .Y(n4367) );
  OAI2BB2XL U4088 ( .B0(n6727), .B1(n421), .A0N(\ram[236][10] ), .A1N(n6374), 
        .Y(n4368) );
  OAI2BB2XL U4089 ( .B0(n6704), .B1(n421), .A0N(\ram[236][11] ), .A1N(n6374), 
        .Y(n4369) );
  OAI2BB2XL U4090 ( .B0(n6681), .B1(n421), .A0N(\ram[236][12] ), .A1N(n6374), 
        .Y(n4370) );
  OAI2BB2XL U4091 ( .B0(n6658), .B1(n421), .A0N(\ram[236][13] ), .A1N(n6374), 
        .Y(n4371) );
  OAI2BB2XL U4092 ( .B0(n6635), .B1(n421), .A0N(\ram[236][14] ), .A1N(n6374), 
        .Y(n4372) );
  OAI2BB2XL U4093 ( .B0(n6612), .B1(n421), .A0N(\ram[236][15] ), .A1N(n6374), 
        .Y(n4373) );
  OAI2BB2XL U4094 ( .B0(n6960), .B1(n423), .A0N(\ram[237][0] ), .A1N(n6373), 
        .Y(n4374) );
  OAI2BB2XL U4095 ( .B0(n6937), .B1(n423), .A0N(\ram[237][1] ), .A1N(n6373), 
        .Y(n4375) );
  OAI2BB2XL U4096 ( .B0(n6914), .B1(n423), .A0N(\ram[237][2] ), .A1N(n6373), 
        .Y(n4376) );
  OAI2BB2XL U4097 ( .B0(n6891), .B1(n423), .A0N(\ram[237][3] ), .A1N(n6373), 
        .Y(n4377) );
  OAI2BB2XL U4098 ( .B0(n6865), .B1(n423), .A0N(\ram[237][4] ), .A1N(n6373), 
        .Y(n4378) );
  OAI2BB2XL U4099 ( .B0(n6842), .B1(n423), .A0N(\ram[237][5] ), .A1N(n6373), 
        .Y(n4379) );
  OAI2BB2XL U4100 ( .B0(n6819), .B1(n423), .A0N(\ram[237][6] ), .A1N(n6373), 
        .Y(n4380) );
  OAI2BB2XL U4101 ( .B0(n6796), .B1(n423), .A0N(\ram[237][7] ), .A1N(n6373), 
        .Y(n4381) );
  OAI2BB2XL U4102 ( .B0(n6773), .B1(n423), .A0N(\ram[237][8] ), .A1N(n6373), 
        .Y(n4382) );
  OAI2BB2XL U4103 ( .B0(n6750), .B1(n423), .A0N(\ram[237][9] ), .A1N(n6373), 
        .Y(n4383) );
  OAI2BB2XL U4104 ( .B0(n6727), .B1(n423), .A0N(\ram[237][10] ), .A1N(n6373), 
        .Y(n4384) );
  OAI2BB2XL U4105 ( .B0(n6704), .B1(n423), .A0N(\ram[237][11] ), .A1N(n6373), 
        .Y(n4385) );
  OAI2BB2XL U4106 ( .B0(n6681), .B1(n423), .A0N(\ram[237][12] ), .A1N(n6373), 
        .Y(n4386) );
  OAI2BB2XL U4107 ( .B0(n6658), .B1(n423), .A0N(\ram[237][13] ), .A1N(n6373), 
        .Y(n4387) );
  OAI2BB2XL U4108 ( .B0(n6635), .B1(n423), .A0N(\ram[237][14] ), .A1N(n6373), 
        .Y(n4388) );
  OAI2BB2XL U4109 ( .B0(n6612), .B1(n423), .A0N(\ram[237][15] ), .A1N(n6373), 
        .Y(n4389) );
  OAI2BB2XL U4110 ( .B0(n6960), .B1(n425), .A0N(\ram[238][0] ), .A1N(n6372), 
        .Y(n4390) );
  OAI2BB2XL U4111 ( .B0(n6937), .B1(n425), .A0N(\ram[238][1] ), .A1N(n6372), 
        .Y(n4391) );
  OAI2BB2XL U4112 ( .B0(n6914), .B1(n425), .A0N(\ram[238][2] ), .A1N(n6372), 
        .Y(n4392) );
  OAI2BB2XL U4113 ( .B0(n6891), .B1(n425), .A0N(\ram[238][3] ), .A1N(n6372), 
        .Y(n4393) );
  OAI2BB2XL U4114 ( .B0(n6865), .B1(n425), .A0N(\ram[238][4] ), .A1N(n6372), 
        .Y(n4394) );
  OAI2BB2XL U4115 ( .B0(n6842), .B1(n425), .A0N(\ram[238][5] ), .A1N(n6372), 
        .Y(n4395) );
  OAI2BB2XL U4116 ( .B0(n6819), .B1(n425), .A0N(\ram[238][6] ), .A1N(n6372), 
        .Y(n4396) );
  OAI2BB2XL U4117 ( .B0(n6796), .B1(n425), .A0N(\ram[238][7] ), .A1N(n6372), 
        .Y(n4397) );
  OAI2BB2XL U4118 ( .B0(n6773), .B1(n425), .A0N(\ram[238][8] ), .A1N(n6372), 
        .Y(n4398) );
  OAI2BB2XL U4119 ( .B0(n6750), .B1(n425), .A0N(\ram[238][9] ), .A1N(n6372), 
        .Y(n4399) );
  OAI2BB2XL U4120 ( .B0(n6727), .B1(n425), .A0N(\ram[238][10] ), .A1N(n6372), 
        .Y(n4400) );
  OAI2BB2XL U4121 ( .B0(n6704), .B1(n425), .A0N(\ram[238][11] ), .A1N(n6372), 
        .Y(n4401) );
  OAI2BB2XL U4122 ( .B0(n6681), .B1(n425), .A0N(\ram[238][12] ), .A1N(n6372), 
        .Y(n4402) );
  OAI2BB2XL U4123 ( .B0(n6658), .B1(n425), .A0N(\ram[238][13] ), .A1N(n6372), 
        .Y(n4403) );
  OAI2BB2XL U4124 ( .B0(n6635), .B1(n425), .A0N(\ram[238][14] ), .A1N(n6372), 
        .Y(n4404) );
  OAI2BB2XL U4125 ( .B0(n6612), .B1(n425), .A0N(\ram[238][15] ), .A1N(n6372), 
        .Y(n4405) );
  OAI2BB2XL U4126 ( .B0(n6960), .B1(n427), .A0N(\ram[239][0] ), .A1N(n6371), 
        .Y(n4406) );
  OAI2BB2XL U4127 ( .B0(n6937), .B1(n427), .A0N(\ram[239][1] ), .A1N(n6371), 
        .Y(n4407) );
  OAI2BB2XL U4128 ( .B0(n6914), .B1(n427), .A0N(\ram[239][2] ), .A1N(n6371), 
        .Y(n4408) );
  OAI2BB2XL U4129 ( .B0(n6891), .B1(n427), .A0N(\ram[239][3] ), .A1N(n6371), 
        .Y(n4409) );
  OAI2BB2XL U4130 ( .B0(n6865), .B1(n427), .A0N(\ram[239][4] ), .A1N(n6371), 
        .Y(n4410) );
  OAI2BB2XL U4131 ( .B0(n6842), .B1(n427), .A0N(\ram[239][5] ), .A1N(n6371), 
        .Y(n4411) );
  OAI2BB2XL U4132 ( .B0(n6819), .B1(n427), .A0N(\ram[239][6] ), .A1N(n6371), 
        .Y(n4412) );
  OAI2BB2XL U4133 ( .B0(n6796), .B1(n427), .A0N(\ram[239][7] ), .A1N(n6371), 
        .Y(n4413) );
  OAI2BB2XL U4134 ( .B0(n6773), .B1(n427), .A0N(\ram[239][8] ), .A1N(n6371), 
        .Y(n4414) );
  OAI2BB2XL U4135 ( .B0(n6750), .B1(n427), .A0N(\ram[239][9] ), .A1N(n6371), 
        .Y(n4415) );
  OAI2BB2XL U4136 ( .B0(n6727), .B1(n427), .A0N(\ram[239][10] ), .A1N(n6371), 
        .Y(n4416) );
  OAI2BB2XL U4137 ( .B0(n6704), .B1(n427), .A0N(\ram[239][11] ), .A1N(n6371), 
        .Y(n4417) );
  OAI2BB2XL U4138 ( .B0(n6681), .B1(n427), .A0N(\ram[239][12] ), .A1N(n6371), 
        .Y(n4418) );
  OAI2BB2XL U4139 ( .B0(n6658), .B1(n427), .A0N(\ram[239][13] ), .A1N(n6371), 
        .Y(n4419) );
  OAI2BB2XL U4140 ( .B0(n6635), .B1(n427), .A0N(\ram[239][14] ), .A1N(n6371), 
        .Y(n4420) );
  OAI2BB2XL U4141 ( .B0(n6612), .B1(n427), .A0N(\ram[239][15] ), .A1N(n6371), 
        .Y(n4421) );
  OAI2BB2XL U4142 ( .B0(n6960), .B1(n429), .A0N(\ram[240][0] ), .A1N(n6370), 
        .Y(n4422) );
  OAI2BB2XL U4143 ( .B0(n6937), .B1(n429), .A0N(\ram[240][1] ), .A1N(n6370), 
        .Y(n4423) );
  OAI2BB2XL U4144 ( .B0(n6914), .B1(n429), .A0N(\ram[240][2] ), .A1N(n6370), 
        .Y(n4424) );
  OAI2BB2XL U4145 ( .B0(n6891), .B1(n429), .A0N(\ram[240][3] ), .A1N(n6370), 
        .Y(n4425) );
  OAI2BB2XL U4146 ( .B0(n6865), .B1(n429), .A0N(\ram[240][4] ), .A1N(n6370), 
        .Y(n4426) );
  OAI2BB2XL U4147 ( .B0(n6842), .B1(n429), .A0N(\ram[240][5] ), .A1N(n6370), 
        .Y(n4427) );
  OAI2BB2XL U4148 ( .B0(n6819), .B1(n429), .A0N(\ram[240][6] ), .A1N(n6370), 
        .Y(n4428) );
  OAI2BB2XL U4149 ( .B0(n6796), .B1(n429), .A0N(\ram[240][7] ), .A1N(n6370), 
        .Y(n4429) );
  OAI2BB2XL U4150 ( .B0(n6773), .B1(n429), .A0N(\ram[240][8] ), .A1N(n6370), 
        .Y(n4430) );
  OAI2BB2XL U4151 ( .B0(n6750), .B1(n429), .A0N(\ram[240][9] ), .A1N(n6370), 
        .Y(n4431) );
  OAI2BB2XL U4152 ( .B0(n6727), .B1(n429), .A0N(\ram[240][10] ), .A1N(n6370), 
        .Y(n4432) );
  OAI2BB2XL U4153 ( .B0(n6704), .B1(n429), .A0N(\ram[240][11] ), .A1N(n6370), 
        .Y(n4433) );
  OAI2BB2XL U4154 ( .B0(n6681), .B1(n429), .A0N(\ram[240][12] ), .A1N(n6370), 
        .Y(n4434) );
  OAI2BB2XL U4155 ( .B0(n6658), .B1(n429), .A0N(\ram[240][13] ), .A1N(n6370), 
        .Y(n4435) );
  OAI2BB2XL U4156 ( .B0(n6635), .B1(n429), .A0N(\ram[240][14] ), .A1N(n6370), 
        .Y(n4436) );
  OAI2BB2XL U4157 ( .B0(n6612), .B1(n429), .A0N(\ram[240][15] ), .A1N(n6370), 
        .Y(n4437) );
  OAI2BB2XL U4158 ( .B0(n6960), .B1(n431), .A0N(\ram[241][0] ), .A1N(n6369), 
        .Y(n4438) );
  OAI2BB2XL U4159 ( .B0(n6937), .B1(n431), .A0N(\ram[241][1] ), .A1N(n6369), 
        .Y(n4439) );
  OAI2BB2XL U4160 ( .B0(n6914), .B1(n431), .A0N(\ram[241][2] ), .A1N(n6369), 
        .Y(n4440) );
  OAI2BB2XL U4161 ( .B0(n6891), .B1(n431), .A0N(\ram[241][3] ), .A1N(n6369), 
        .Y(n4441) );
  OAI2BB2XL U4162 ( .B0(n6865), .B1(n431), .A0N(\ram[241][4] ), .A1N(n6369), 
        .Y(n4442) );
  OAI2BB2XL U4163 ( .B0(n6842), .B1(n431), .A0N(\ram[241][5] ), .A1N(n6369), 
        .Y(n4443) );
  OAI2BB2XL U4164 ( .B0(n6819), .B1(n431), .A0N(\ram[241][6] ), .A1N(n6369), 
        .Y(n4444) );
  OAI2BB2XL U4165 ( .B0(n6796), .B1(n431), .A0N(\ram[241][7] ), .A1N(n6369), 
        .Y(n4445) );
  OAI2BB2XL U4166 ( .B0(n6773), .B1(n431), .A0N(\ram[241][8] ), .A1N(n6369), 
        .Y(n4446) );
  OAI2BB2XL U4167 ( .B0(n6750), .B1(n431), .A0N(\ram[241][9] ), .A1N(n6369), 
        .Y(n4447) );
  OAI2BB2XL U4168 ( .B0(n6727), .B1(n431), .A0N(\ram[241][10] ), .A1N(n6369), 
        .Y(n4448) );
  OAI2BB2XL U4169 ( .B0(n6704), .B1(n431), .A0N(\ram[241][11] ), .A1N(n6369), 
        .Y(n4449) );
  OAI2BB2XL U4170 ( .B0(n6681), .B1(n431), .A0N(\ram[241][12] ), .A1N(n6369), 
        .Y(n4450) );
  OAI2BB2XL U4171 ( .B0(n6658), .B1(n431), .A0N(\ram[241][13] ), .A1N(n6369), 
        .Y(n4451) );
  OAI2BB2XL U4172 ( .B0(n6635), .B1(n431), .A0N(\ram[241][14] ), .A1N(n6369), 
        .Y(n4452) );
  OAI2BB2XL U4173 ( .B0(n6612), .B1(n431), .A0N(\ram[241][15] ), .A1N(n6369), 
        .Y(n4453) );
  OAI2BB2XL U4174 ( .B0(n6960), .B1(n433), .A0N(\ram[242][0] ), .A1N(n6368), 
        .Y(n4454) );
  OAI2BB2XL U4175 ( .B0(n6937), .B1(n433), .A0N(\ram[242][1] ), .A1N(n6368), 
        .Y(n4455) );
  OAI2BB2XL U4176 ( .B0(n6914), .B1(n433), .A0N(\ram[242][2] ), .A1N(n6368), 
        .Y(n4456) );
  OAI2BB2XL U4177 ( .B0(n6891), .B1(n433), .A0N(\ram[242][3] ), .A1N(n6368), 
        .Y(n4457) );
  OAI2BB2XL U4178 ( .B0(n6865), .B1(n433), .A0N(\ram[242][4] ), .A1N(n6368), 
        .Y(n4458) );
  OAI2BB2XL U4179 ( .B0(n6842), .B1(n433), .A0N(\ram[242][5] ), .A1N(n6368), 
        .Y(n4459) );
  OAI2BB2XL U4180 ( .B0(n6819), .B1(n433), .A0N(\ram[242][6] ), .A1N(n6368), 
        .Y(n4460) );
  OAI2BB2XL U4181 ( .B0(n6796), .B1(n433), .A0N(\ram[242][7] ), .A1N(n6368), 
        .Y(n4461) );
  OAI2BB2XL U4182 ( .B0(n6773), .B1(n433), .A0N(\ram[242][8] ), .A1N(n6368), 
        .Y(n4462) );
  OAI2BB2XL U4183 ( .B0(n6750), .B1(n433), .A0N(\ram[242][9] ), .A1N(n6368), 
        .Y(n4463) );
  OAI2BB2XL U4184 ( .B0(n6727), .B1(n433), .A0N(\ram[242][10] ), .A1N(n6368), 
        .Y(n4464) );
  OAI2BB2XL U4185 ( .B0(n6704), .B1(n433), .A0N(\ram[242][11] ), .A1N(n6368), 
        .Y(n4465) );
  OAI2BB2XL U4186 ( .B0(n6681), .B1(n433), .A0N(\ram[242][12] ), .A1N(n6368), 
        .Y(n4466) );
  OAI2BB2XL U4187 ( .B0(n6658), .B1(n433), .A0N(\ram[242][13] ), .A1N(n6368), 
        .Y(n4467) );
  OAI2BB2XL U4188 ( .B0(n6635), .B1(n433), .A0N(\ram[242][14] ), .A1N(n6368), 
        .Y(n4468) );
  OAI2BB2XL U4189 ( .B0(n6612), .B1(n433), .A0N(\ram[242][15] ), .A1N(n6368), 
        .Y(n4469) );
  OAI2BB2XL U4190 ( .B0(n6960), .B1(n435), .A0N(\ram[243][0] ), .A1N(n6367), 
        .Y(n4470) );
  OAI2BB2XL U4191 ( .B0(n6937), .B1(n435), .A0N(\ram[243][1] ), .A1N(n6367), 
        .Y(n4471) );
  OAI2BB2XL U4192 ( .B0(n6914), .B1(n435), .A0N(\ram[243][2] ), .A1N(n6367), 
        .Y(n4472) );
  OAI2BB2XL U4193 ( .B0(n6891), .B1(n435), .A0N(\ram[243][3] ), .A1N(n6367), 
        .Y(n4473) );
  OAI2BB2XL U4194 ( .B0(n6865), .B1(n435), .A0N(\ram[243][4] ), .A1N(n6367), 
        .Y(n4474) );
  OAI2BB2XL U4195 ( .B0(n6842), .B1(n435), .A0N(\ram[243][5] ), .A1N(n6367), 
        .Y(n4475) );
  OAI2BB2XL U4196 ( .B0(n6819), .B1(n435), .A0N(\ram[243][6] ), .A1N(n6367), 
        .Y(n4476) );
  OAI2BB2XL U4197 ( .B0(n6796), .B1(n435), .A0N(\ram[243][7] ), .A1N(n6367), 
        .Y(n4477) );
  OAI2BB2XL U4198 ( .B0(n6773), .B1(n435), .A0N(\ram[243][8] ), .A1N(n6367), 
        .Y(n4478) );
  OAI2BB2XL U4199 ( .B0(n6750), .B1(n435), .A0N(\ram[243][9] ), .A1N(n6367), 
        .Y(n4479) );
  OAI2BB2XL U4200 ( .B0(n6727), .B1(n435), .A0N(\ram[243][10] ), .A1N(n6367), 
        .Y(n4480) );
  OAI2BB2XL U4201 ( .B0(n6704), .B1(n435), .A0N(\ram[243][11] ), .A1N(n6367), 
        .Y(n4481) );
  OAI2BB2XL U4202 ( .B0(n6681), .B1(n435), .A0N(\ram[243][12] ), .A1N(n6367), 
        .Y(n4482) );
  OAI2BB2XL U4203 ( .B0(n6658), .B1(n435), .A0N(\ram[243][13] ), .A1N(n6367), 
        .Y(n4483) );
  OAI2BB2XL U4204 ( .B0(n6635), .B1(n435), .A0N(\ram[243][14] ), .A1N(n6367), 
        .Y(n4484) );
  OAI2BB2XL U4205 ( .B0(n6612), .B1(n435), .A0N(\ram[243][15] ), .A1N(n6367), 
        .Y(n4485) );
  OAI2BB2XL U4206 ( .B0(n6959), .B1(n437), .A0N(\ram[244][0] ), .A1N(n6366), 
        .Y(n4486) );
  OAI2BB2XL U4207 ( .B0(n6936), .B1(n437), .A0N(\ram[244][1] ), .A1N(n6366), 
        .Y(n4487) );
  OAI2BB2XL U4208 ( .B0(n6913), .B1(n437), .A0N(\ram[244][2] ), .A1N(n6366), 
        .Y(n4488) );
  OAI2BB2XL U4209 ( .B0(n6890), .B1(n437), .A0N(\ram[244][3] ), .A1N(n6366), 
        .Y(n4489) );
  OAI2BB2XL U4210 ( .B0(n6865), .B1(n437), .A0N(\ram[244][4] ), .A1N(n6366), 
        .Y(n4490) );
  OAI2BB2XL U4211 ( .B0(n6842), .B1(n437), .A0N(\ram[244][5] ), .A1N(n6366), 
        .Y(n4491) );
  OAI2BB2XL U4212 ( .B0(n6819), .B1(n437), .A0N(\ram[244][6] ), .A1N(n6366), 
        .Y(n4492) );
  OAI2BB2XL U4213 ( .B0(n6796), .B1(n437), .A0N(\ram[244][7] ), .A1N(n6366), 
        .Y(n4493) );
  OAI2BB2XL U4214 ( .B0(n6773), .B1(n437), .A0N(\ram[244][8] ), .A1N(n6366), 
        .Y(n4494) );
  OAI2BB2XL U4215 ( .B0(n6750), .B1(n437), .A0N(\ram[244][9] ), .A1N(n6366), 
        .Y(n4495) );
  OAI2BB2XL U4216 ( .B0(n6727), .B1(n437), .A0N(\ram[244][10] ), .A1N(n6366), 
        .Y(n4496) );
  OAI2BB2XL U4217 ( .B0(n6704), .B1(n437), .A0N(\ram[244][11] ), .A1N(n6366), 
        .Y(n4497) );
  OAI2BB2XL U4218 ( .B0(n6681), .B1(n437), .A0N(\ram[244][12] ), .A1N(n6366), 
        .Y(n4498) );
  OAI2BB2XL U4219 ( .B0(n6658), .B1(n437), .A0N(\ram[244][13] ), .A1N(n6366), 
        .Y(n4499) );
  OAI2BB2XL U4220 ( .B0(n6635), .B1(n437), .A0N(\ram[244][14] ), .A1N(n6366), 
        .Y(n4500) );
  OAI2BB2XL U4221 ( .B0(n6612), .B1(n437), .A0N(\ram[244][15] ), .A1N(n6366), 
        .Y(n4501) );
  OAI2BB2XL U4222 ( .B0(n6959), .B1(n439), .A0N(\ram[245][0] ), .A1N(n6365), 
        .Y(n4502) );
  OAI2BB2XL U4223 ( .B0(n6936), .B1(n439), .A0N(\ram[245][1] ), .A1N(n6365), 
        .Y(n4503) );
  OAI2BB2XL U4224 ( .B0(n6913), .B1(n439), .A0N(\ram[245][2] ), .A1N(n6365), 
        .Y(n4504) );
  OAI2BB2XL U4225 ( .B0(n6890), .B1(n439), .A0N(\ram[245][3] ), .A1N(n6365), 
        .Y(n4505) );
  OAI2BB2XL U4226 ( .B0(n6866), .B1(n439), .A0N(\ram[245][4] ), .A1N(n6365), 
        .Y(n4506) );
  OAI2BB2XL U4227 ( .B0(n6843), .B1(n439), .A0N(\ram[245][5] ), .A1N(n6365), 
        .Y(n4507) );
  OAI2BB2XL U4228 ( .B0(n6820), .B1(n439), .A0N(\ram[245][6] ), .A1N(n6365), 
        .Y(n4508) );
  OAI2BB2XL U4229 ( .B0(n6797), .B1(n439), .A0N(\ram[245][7] ), .A1N(n6365), 
        .Y(n4509) );
  OAI2BB2XL U4230 ( .B0(n6774), .B1(n439), .A0N(\ram[245][8] ), .A1N(n6365), 
        .Y(n4510) );
  OAI2BB2XL U4231 ( .B0(n6751), .B1(n439), .A0N(\ram[245][9] ), .A1N(n6365), 
        .Y(n4511) );
  OAI2BB2XL U4232 ( .B0(n6728), .B1(n439), .A0N(\ram[245][10] ), .A1N(n6365), 
        .Y(n4512) );
  OAI2BB2XL U4233 ( .B0(n6705), .B1(n439), .A0N(\ram[245][11] ), .A1N(n6365), 
        .Y(n4513) );
  OAI2BB2XL U4234 ( .B0(n6682), .B1(n439), .A0N(\ram[245][12] ), .A1N(n6365), 
        .Y(n4514) );
  OAI2BB2XL U4235 ( .B0(n6659), .B1(n439), .A0N(\ram[245][13] ), .A1N(n6365), 
        .Y(n4515) );
  OAI2BB2XL U4236 ( .B0(n6636), .B1(n439), .A0N(\ram[245][14] ), .A1N(n6365), 
        .Y(n4516) );
  OAI2BB2XL U4237 ( .B0(n6613), .B1(n439), .A0N(\ram[245][15] ), .A1N(n6365), 
        .Y(n4517) );
  OAI2BB2XL U4238 ( .B0(n6959), .B1(n441), .A0N(\ram[246][0] ), .A1N(n6364), 
        .Y(n4518) );
  OAI2BB2XL U4239 ( .B0(n6936), .B1(n441), .A0N(\ram[246][1] ), .A1N(n6364), 
        .Y(n4519) );
  OAI2BB2XL U4240 ( .B0(n6913), .B1(n441), .A0N(\ram[246][2] ), .A1N(n6364), 
        .Y(n4520) );
  OAI2BB2XL U4241 ( .B0(n6890), .B1(n441), .A0N(\ram[246][3] ), .A1N(n6364), 
        .Y(n4521) );
  OAI2BB2XL U4242 ( .B0(n6871), .B1(n441), .A0N(\ram[246][4] ), .A1N(n6364), 
        .Y(n4522) );
  OAI2BB2XL U4243 ( .B0(n6848), .B1(n441), .A0N(\ram[246][5] ), .A1N(n6364), 
        .Y(n4523) );
  OAI2BB2XL U4244 ( .B0(n6825), .B1(n441), .A0N(\ram[246][6] ), .A1N(n6364), 
        .Y(n4524) );
  OAI2BB2XL U4245 ( .B0(n6802), .B1(n441), .A0N(\ram[246][7] ), .A1N(n6364), 
        .Y(n4525) );
  OAI2BB2XL U4246 ( .B0(n6779), .B1(n441), .A0N(\ram[246][8] ), .A1N(n6364), 
        .Y(n4526) );
  OAI2BB2XL U4247 ( .B0(n6756), .B1(n441), .A0N(\ram[246][9] ), .A1N(n6364), 
        .Y(n4527) );
  OAI2BB2XL U4248 ( .B0(n6733), .B1(n441), .A0N(\ram[246][10] ), .A1N(n6364), 
        .Y(n4528) );
  OAI2BB2XL U4249 ( .B0(n6710), .B1(n441), .A0N(\ram[246][11] ), .A1N(n6364), 
        .Y(n4529) );
  OAI2BB2XL U4250 ( .B0(n6687), .B1(n441), .A0N(\ram[246][12] ), .A1N(n6364), 
        .Y(n4530) );
  OAI2BB2XL U4251 ( .B0(n6664), .B1(n441), .A0N(\ram[246][13] ), .A1N(n6364), 
        .Y(n4531) );
  OAI2BB2XL U4252 ( .B0(n6641), .B1(n441), .A0N(\ram[246][14] ), .A1N(n6364), 
        .Y(n4532) );
  OAI2BB2XL U4253 ( .B0(n6618), .B1(n441), .A0N(\ram[246][15] ), .A1N(n6364), 
        .Y(n4533) );
  OAI2BB2XL U4254 ( .B0(n6959), .B1(n443), .A0N(\ram[247][0] ), .A1N(n6363), 
        .Y(n4534) );
  OAI2BB2XL U4255 ( .B0(n6936), .B1(n443), .A0N(\ram[247][1] ), .A1N(n6363), 
        .Y(n4535) );
  OAI2BB2XL U4256 ( .B0(n6913), .B1(n443), .A0N(\ram[247][2] ), .A1N(n6363), 
        .Y(n4536) );
  OAI2BB2XL U4257 ( .B0(n6890), .B1(n443), .A0N(\ram[247][3] ), .A1N(n6363), 
        .Y(n4537) );
  OAI2BB2XL U4258 ( .B0(n6870), .B1(n443), .A0N(\ram[247][4] ), .A1N(n6363), 
        .Y(n4538) );
  OAI2BB2XL U4259 ( .B0(n6847), .B1(n443), .A0N(\ram[247][5] ), .A1N(n6363), 
        .Y(n4539) );
  OAI2BB2XL U4260 ( .B0(n6824), .B1(n443), .A0N(\ram[247][6] ), .A1N(n6363), 
        .Y(n4540) );
  OAI2BB2XL U4261 ( .B0(n6801), .B1(n443), .A0N(\ram[247][7] ), .A1N(n6363), 
        .Y(n4541) );
  OAI2BB2XL U4262 ( .B0(n6778), .B1(n443), .A0N(\ram[247][8] ), .A1N(n6363), 
        .Y(n4542) );
  OAI2BB2XL U4263 ( .B0(n6755), .B1(n443), .A0N(\ram[247][9] ), .A1N(n6363), 
        .Y(n4543) );
  OAI2BB2XL U4264 ( .B0(n6732), .B1(n443), .A0N(\ram[247][10] ), .A1N(n6363), 
        .Y(n4544) );
  OAI2BB2XL U4265 ( .B0(n6709), .B1(n443), .A0N(\ram[247][11] ), .A1N(n6363), 
        .Y(n4545) );
  OAI2BB2XL U4266 ( .B0(n6686), .B1(n443), .A0N(\ram[247][12] ), .A1N(n6363), 
        .Y(n4546) );
  OAI2BB2XL U4267 ( .B0(n6663), .B1(n443), .A0N(\ram[247][13] ), .A1N(n6363), 
        .Y(n4547) );
  OAI2BB2XL U4268 ( .B0(n6640), .B1(n443), .A0N(\ram[247][14] ), .A1N(n6363), 
        .Y(n4548) );
  OAI2BB2XL U4269 ( .B0(n6617), .B1(n443), .A0N(\ram[247][15] ), .A1N(n6363), 
        .Y(n4549) );
  OAI2BB2XL U4270 ( .B0(n6959), .B1(n444), .A0N(\ram[248][0] ), .A1N(n6362), 
        .Y(n4550) );
  OAI2BB2XL U4271 ( .B0(n6936), .B1(n444), .A0N(\ram[248][1] ), .A1N(n6362), 
        .Y(n4551) );
  OAI2BB2XL U4272 ( .B0(n6913), .B1(n444), .A0N(\ram[248][2] ), .A1N(n6362), 
        .Y(n4552) );
  OAI2BB2XL U4273 ( .B0(n6890), .B1(n444), .A0N(\ram[248][3] ), .A1N(n6362), 
        .Y(n4553) );
  OAI2BB2XL U4274 ( .B0(n6865), .B1(n444), .A0N(\ram[248][4] ), .A1N(n6362), 
        .Y(n4554) );
  OAI2BB2XL U4275 ( .B0(n6842), .B1(n444), .A0N(\ram[248][5] ), .A1N(n6362), 
        .Y(n4555) );
  OAI2BB2XL U4276 ( .B0(n6819), .B1(n444), .A0N(\ram[248][6] ), .A1N(n6362), 
        .Y(n4556) );
  OAI2BB2XL U4277 ( .B0(n6796), .B1(n444), .A0N(\ram[248][7] ), .A1N(n6362), 
        .Y(n4557) );
  OAI2BB2XL U4278 ( .B0(n6773), .B1(n444), .A0N(\ram[248][8] ), .A1N(n6362), 
        .Y(n4558) );
  OAI2BB2XL U4279 ( .B0(n6750), .B1(n444), .A0N(\ram[248][9] ), .A1N(n6362), 
        .Y(n4559) );
  OAI2BB2XL U4280 ( .B0(n6727), .B1(n444), .A0N(\ram[248][10] ), .A1N(n6362), 
        .Y(n4560) );
  OAI2BB2XL U4281 ( .B0(n6704), .B1(n444), .A0N(\ram[248][11] ), .A1N(n6362), 
        .Y(n4561) );
  OAI2BB2XL U4282 ( .B0(n6681), .B1(n444), .A0N(\ram[248][12] ), .A1N(n6362), 
        .Y(n4562) );
  OAI2BB2XL U4283 ( .B0(n6658), .B1(n444), .A0N(\ram[248][13] ), .A1N(n6362), 
        .Y(n4563) );
  OAI2BB2XL U4284 ( .B0(n6635), .B1(n444), .A0N(\ram[248][14] ), .A1N(n6362), 
        .Y(n4564) );
  OAI2BB2XL U4285 ( .B0(n6612), .B1(n444), .A0N(\ram[248][15] ), .A1N(n6362), 
        .Y(n4565) );
  OAI2BB2XL U4286 ( .B0(n6959), .B1(n446), .A0N(\ram[249][0] ), .A1N(n6361), 
        .Y(n4566) );
  OAI2BB2XL U4287 ( .B0(n6936), .B1(n446), .A0N(\ram[249][1] ), .A1N(n6361), 
        .Y(n4567) );
  OAI2BB2XL U4288 ( .B0(n6913), .B1(n446), .A0N(\ram[249][2] ), .A1N(n6361), 
        .Y(n4568) );
  OAI2BB2XL U4289 ( .B0(n6890), .B1(n446), .A0N(\ram[249][3] ), .A1N(n6361), 
        .Y(n4569) );
  OAI2BB2XL U4290 ( .B0(n6866), .B1(n446), .A0N(\ram[249][4] ), .A1N(n6361), 
        .Y(n4570) );
  OAI2BB2XL U4291 ( .B0(n6843), .B1(n446), .A0N(\ram[249][5] ), .A1N(n6361), 
        .Y(n4571) );
  OAI2BB2XL U4292 ( .B0(n6820), .B1(n446), .A0N(\ram[249][6] ), .A1N(n6361), 
        .Y(n4572) );
  OAI2BB2XL U4293 ( .B0(n6797), .B1(n446), .A0N(\ram[249][7] ), .A1N(n6361), 
        .Y(n4573) );
  OAI2BB2XL U4294 ( .B0(n6774), .B1(n446), .A0N(\ram[249][8] ), .A1N(n6361), 
        .Y(n4574) );
  OAI2BB2XL U4295 ( .B0(n6751), .B1(n446), .A0N(\ram[249][9] ), .A1N(n6361), 
        .Y(n4575) );
  OAI2BB2XL U4296 ( .B0(n6728), .B1(n446), .A0N(\ram[249][10] ), .A1N(n6361), 
        .Y(n4576) );
  OAI2BB2XL U4297 ( .B0(n6705), .B1(n446), .A0N(\ram[249][11] ), .A1N(n6361), 
        .Y(n4577) );
  OAI2BB2XL U4298 ( .B0(n6682), .B1(n446), .A0N(\ram[249][12] ), .A1N(n6361), 
        .Y(n4578) );
  OAI2BB2XL U4299 ( .B0(n6659), .B1(n446), .A0N(\ram[249][13] ), .A1N(n6361), 
        .Y(n4579) );
  OAI2BB2XL U4300 ( .B0(n6636), .B1(n446), .A0N(\ram[249][14] ), .A1N(n6361), 
        .Y(n4580) );
  OAI2BB2XL U4301 ( .B0(n6613), .B1(n446), .A0N(\ram[249][15] ), .A1N(n6361), 
        .Y(n4581) );
  OAI2BB2XL U4302 ( .B0(n6959), .B1(n448), .A0N(\ram[250][0] ), .A1N(n6360), 
        .Y(n4582) );
  OAI2BB2XL U4303 ( .B0(n6936), .B1(n448), .A0N(\ram[250][1] ), .A1N(n6360), 
        .Y(n4583) );
  OAI2BB2XL U4304 ( .B0(n6913), .B1(n448), .A0N(\ram[250][2] ), .A1N(n6360), 
        .Y(n4584) );
  OAI2BB2XL U4305 ( .B0(n6890), .B1(n448), .A0N(\ram[250][3] ), .A1N(n6360), 
        .Y(n4585) );
  OAI2BB2XL U4306 ( .B0(n6871), .B1(n448), .A0N(\ram[250][4] ), .A1N(n6360), 
        .Y(n4586) );
  OAI2BB2XL U4307 ( .B0(n6848), .B1(n448), .A0N(\ram[250][5] ), .A1N(n6360), 
        .Y(n4587) );
  OAI2BB2XL U4308 ( .B0(n6825), .B1(n448), .A0N(\ram[250][6] ), .A1N(n6360), 
        .Y(n4588) );
  OAI2BB2XL U4309 ( .B0(n6802), .B1(n448), .A0N(\ram[250][7] ), .A1N(n6360), 
        .Y(n4589) );
  OAI2BB2XL U4310 ( .B0(n6779), .B1(n448), .A0N(\ram[250][8] ), .A1N(n6360), 
        .Y(n4590) );
  OAI2BB2XL U4311 ( .B0(n6756), .B1(n448), .A0N(\ram[250][9] ), .A1N(n6360), 
        .Y(n4591) );
  OAI2BB2XL U4312 ( .B0(n6733), .B1(n448), .A0N(\ram[250][10] ), .A1N(n6360), 
        .Y(n4592) );
  OAI2BB2XL U4313 ( .B0(n6710), .B1(n448), .A0N(\ram[250][11] ), .A1N(n6360), 
        .Y(n4593) );
  OAI2BB2XL U4314 ( .B0(n6687), .B1(n448), .A0N(\ram[250][12] ), .A1N(n6360), 
        .Y(n4594) );
  OAI2BB2XL U4315 ( .B0(n6664), .B1(n448), .A0N(\ram[250][13] ), .A1N(n6360), 
        .Y(n4595) );
  OAI2BB2XL U4316 ( .B0(n6641), .B1(n448), .A0N(\ram[250][14] ), .A1N(n6360), 
        .Y(n4596) );
  OAI2BB2XL U4317 ( .B0(n6618), .B1(n448), .A0N(\ram[250][15] ), .A1N(n6360), 
        .Y(n4597) );
  OAI2BB2XL U4318 ( .B0(n6959), .B1(n450), .A0N(\ram[251][0] ), .A1N(n6359), 
        .Y(n4598) );
  OAI2BB2XL U4319 ( .B0(n6936), .B1(n450), .A0N(\ram[251][1] ), .A1N(n6359), 
        .Y(n4599) );
  OAI2BB2XL U4320 ( .B0(n6913), .B1(n450), .A0N(\ram[251][2] ), .A1N(n6359), 
        .Y(n4600) );
  OAI2BB2XL U4321 ( .B0(n6890), .B1(n450), .A0N(\ram[251][3] ), .A1N(n6359), 
        .Y(n4601) );
  OAI2BB2XL U4322 ( .B0(n6870), .B1(n450), .A0N(\ram[251][4] ), .A1N(n6359), 
        .Y(n4602) );
  OAI2BB2XL U4323 ( .B0(n6847), .B1(n450), .A0N(\ram[251][5] ), .A1N(n6359), 
        .Y(n4603) );
  OAI2BB2XL U4324 ( .B0(n6824), .B1(n450), .A0N(\ram[251][6] ), .A1N(n6359), 
        .Y(n4604) );
  OAI2BB2XL U4325 ( .B0(n6801), .B1(n450), .A0N(\ram[251][7] ), .A1N(n6359), 
        .Y(n4605) );
  OAI2BB2XL U4326 ( .B0(n6778), .B1(n450), .A0N(\ram[251][8] ), .A1N(n6359), 
        .Y(n4606) );
  OAI2BB2XL U4327 ( .B0(n6755), .B1(n450), .A0N(\ram[251][9] ), .A1N(n6359), 
        .Y(n4607) );
  OAI2BB2XL U4328 ( .B0(n6732), .B1(n450), .A0N(\ram[251][10] ), .A1N(n6359), 
        .Y(n4608) );
  OAI2BB2XL U4329 ( .B0(n6709), .B1(n450), .A0N(\ram[251][11] ), .A1N(n6359), 
        .Y(n4609) );
  OAI2BB2XL U4330 ( .B0(n6686), .B1(n450), .A0N(\ram[251][12] ), .A1N(n6359), 
        .Y(n4610) );
  OAI2BB2XL U4331 ( .B0(n6663), .B1(n450), .A0N(\ram[251][13] ), .A1N(n6359), 
        .Y(n4611) );
  OAI2BB2XL U4332 ( .B0(n6640), .B1(n450), .A0N(\ram[251][14] ), .A1N(n6359), 
        .Y(n4612) );
  OAI2BB2XL U4333 ( .B0(n6617), .B1(n450), .A0N(\ram[251][15] ), .A1N(n6359), 
        .Y(n4613) );
  OAI2BB2XL U4334 ( .B0(n6959), .B1(n452), .A0N(\ram[252][0] ), .A1N(n6358), 
        .Y(n4614) );
  OAI2BB2XL U4335 ( .B0(n6936), .B1(n452), .A0N(\ram[252][1] ), .A1N(n6358), 
        .Y(n4615) );
  OAI2BB2XL U4336 ( .B0(n6913), .B1(n452), .A0N(\ram[252][2] ), .A1N(n6358), 
        .Y(n4616) );
  OAI2BB2XL U4337 ( .B0(n6890), .B1(n452), .A0N(\ram[252][3] ), .A1N(n6358), 
        .Y(n4617) );
  OAI2BB2XL U4338 ( .B0(n6865), .B1(n452), .A0N(\ram[252][4] ), .A1N(n6358), 
        .Y(n4618) );
  OAI2BB2XL U4339 ( .B0(n6842), .B1(n452), .A0N(\ram[252][5] ), .A1N(n6358), 
        .Y(n4619) );
  OAI2BB2XL U4340 ( .B0(n6819), .B1(n452), .A0N(\ram[252][6] ), .A1N(n6358), 
        .Y(n4620) );
  OAI2BB2XL U4341 ( .B0(n6796), .B1(n452), .A0N(\ram[252][7] ), .A1N(n6358), 
        .Y(n4621) );
  OAI2BB2XL U4342 ( .B0(n6773), .B1(n452), .A0N(\ram[252][8] ), .A1N(n6358), 
        .Y(n4622) );
  OAI2BB2XL U4343 ( .B0(n6750), .B1(n452), .A0N(\ram[252][9] ), .A1N(n6358), 
        .Y(n4623) );
  OAI2BB2XL U4344 ( .B0(n6727), .B1(n452), .A0N(\ram[252][10] ), .A1N(n6358), 
        .Y(n4624) );
  OAI2BB2XL U4345 ( .B0(n6704), .B1(n452), .A0N(\ram[252][11] ), .A1N(n6358), 
        .Y(n4625) );
  OAI2BB2XL U4346 ( .B0(n6681), .B1(n452), .A0N(\ram[252][12] ), .A1N(n6358), 
        .Y(n4626) );
  OAI2BB2XL U4347 ( .B0(n6658), .B1(n452), .A0N(\ram[252][13] ), .A1N(n6358), 
        .Y(n4627) );
  OAI2BB2XL U4348 ( .B0(n6635), .B1(n452), .A0N(\ram[252][14] ), .A1N(n6358), 
        .Y(n4628) );
  OAI2BB2XL U4349 ( .B0(n6612), .B1(n452), .A0N(\ram[252][15] ), .A1N(n6358), 
        .Y(n4629) );
  OAI2BB2XL U4350 ( .B0(n6959), .B1(n454), .A0N(\ram[253][0] ), .A1N(n6357), 
        .Y(n4630) );
  OAI2BB2XL U4351 ( .B0(n6936), .B1(n454), .A0N(\ram[253][1] ), .A1N(n6357), 
        .Y(n4631) );
  OAI2BB2XL U4352 ( .B0(n6913), .B1(n454), .A0N(\ram[253][2] ), .A1N(n6357), 
        .Y(n4632) );
  OAI2BB2XL U4353 ( .B0(n6890), .B1(n454), .A0N(\ram[253][3] ), .A1N(n6357), 
        .Y(n4633) );
  OAI2BB2XL U4354 ( .B0(n6866), .B1(n454), .A0N(\ram[253][4] ), .A1N(n6357), 
        .Y(n4634) );
  OAI2BB2XL U4355 ( .B0(n6843), .B1(n454), .A0N(\ram[253][5] ), .A1N(n6357), 
        .Y(n4635) );
  OAI2BB2XL U4356 ( .B0(n6820), .B1(n454), .A0N(\ram[253][6] ), .A1N(n6357), 
        .Y(n4636) );
  OAI2BB2XL U4357 ( .B0(n6797), .B1(n454), .A0N(\ram[253][7] ), .A1N(n6357), 
        .Y(n4637) );
  OAI2BB2XL U4358 ( .B0(n6774), .B1(n454), .A0N(\ram[253][8] ), .A1N(n6357), 
        .Y(n4638) );
  OAI2BB2XL U4359 ( .B0(n6751), .B1(n454), .A0N(\ram[253][9] ), .A1N(n6357), 
        .Y(n4639) );
  OAI2BB2XL U4360 ( .B0(n6728), .B1(n454), .A0N(\ram[253][10] ), .A1N(n6357), 
        .Y(n4640) );
  OAI2BB2XL U4361 ( .B0(n6705), .B1(n454), .A0N(\ram[253][11] ), .A1N(n6357), 
        .Y(n4641) );
  OAI2BB2XL U4362 ( .B0(n6682), .B1(n454), .A0N(\ram[253][12] ), .A1N(n6357), 
        .Y(n4642) );
  OAI2BB2XL U4363 ( .B0(n6659), .B1(n454), .A0N(\ram[253][13] ), .A1N(n6357), 
        .Y(n4643) );
  OAI2BB2XL U4364 ( .B0(n6636), .B1(n454), .A0N(\ram[253][14] ), .A1N(n6357), 
        .Y(n4644) );
  OAI2BB2XL U4365 ( .B0(n6613), .B1(n454), .A0N(\ram[253][15] ), .A1N(n6357), 
        .Y(n4645) );
  OAI2BB2XL U4366 ( .B0(n6959), .B1(n456), .A0N(\ram[254][0] ), .A1N(n6356), 
        .Y(n4646) );
  OAI2BB2XL U4367 ( .B0(n6936), .B1(n456), .A0N(\ram[254][1] ), .A1N(n6356), 
        .Y(n4647) );
  OAI2BB2XL U4368 ( .B0(n6913), .B1(n456), .A0N(\ram[254][2] ), .A1N(n6356), 
        .Y(n4648) );
  OAI2BB2XL U4369 ( .B0(n6890), .B1(n456), .A0N(\ram[254][3] ), .A1N(n6356), 
        .Y(n4649) );
  OAI2BB2XL U4370 ( .B0(n6871), .B1(n456), .A0N(\ram[254][4] ), .A1N(n6356), 
        .Y(n4650) );
  OAI2BB2XL U4371 ( .B0(n6848), .B1(n456), .A0N(\ram[254][5] ), .A1N(n6356), 
        .Y(n4651) );
  OAI2BB2XL U4372 ( .B0(n6825), .B1(n456), .A0N(\ram[254][6] ), .A1N(n6356), 
        .Y(n4652) );
  OAI2BB2XL U4373 ( .B0(n6802), .B1(n456), .A0N(\ram[254][7] ), .A1N(n6356), 
        .Y(n4653) );
  OAI2BB2XL U4374 ( .B0(n6779), .B1(n456), .A0N(\ram[254][8] ), .A1N(n6356), 
        .Y(n4654) );
  OAI2BB2XL U4375 ( .B0(n6756), .B1(n456), .A0N(\ram[254][9] ), .A1N(n6356), 
        .Y(n4655) );
  OAI2BB2XL U4376 ( .B0(n6733), .B1(n456), .A0N(\ram[254][10] ), .A1N(n6356), 
        .Y(n4656) );
  OAI2BB2XL U4377 ( .B0(n6710), .B1(n456), .A0N(\ram[254][11] ), .A1N(n6356), 
        .Y(n4657) );
  OAI2BB2XL U4378 ( .B0(n6687), .B1(n456), .A0N(\ram[254][12] ), .A1N(n6356), 
        .Y(n4658) );
  OAI2BB2XL U4379 ( .B0(n6664), .B1(n456), .A0N(\ram[254][13] ), .A1N(n6356), 
        .Y(n4659) );
  OAI2BB2XL U4380 ( .B0(n6641), .B1(n456), .A0N(\ram[254][14] ), .A1N(n6356), 
        .Y(n4660) );
  OAI2BB2XL U4381 ( .B0(n6618), .B1(n456), .A0N(\ram[254][15] ), .A1N(n6356), 
        .Y(n4661) );
  OAI2BB2XL U4382 ( .B0(n6959), .B1(n458), .A0N(\ram[255][0] ), .A1N(n6355), 
        .Y(n4662) );
  OAI2BB2XL U4383 ( .B0(n6936), .B1(n458), .A0N(\ram[255][1] ), .A1N(n6355), 
        .Y(n4663) );
  OAI2BB2XL U4384 ( .B0(n6913), .B1(n458), .A0N(\ram[255][2] ), .A1N(n6355), 
        .Y(n4664) );
  OAI2BB2XL U4385 ( .B0(n6890), .B1(n458), .A0N(\ram[255][3] ), .A1N(n6355), 
        .Y(n4665) );
  OAI2BB2XL U4386 ( .B0(n6870), .B1(n458), .A0N(\ram[255][4] ), .A1N(n6355), 
        .Y(n4666) );
  OAI2BB2XL U4387 ( .B0(n6847), .B1(n458), .A0N(\ram[255][5] ), .A1N(n6355), 
        .Y(n4667) );
  OAI2BB2XL U4388 ( .B0(n6824), .B1(n458), .A0N(\ram[255][6] ), .A1N(n6355), 
        .Y(n4668) );
  OAI2BB2XL U4389 ( .B0(n6801), .B1(n458), .A0N(\ram[255][7] ), .A1N(n6355), 
        .Y(n4669) );
  OAI2BB2XL U4390 ( .B0(n6778), .B1(n458), .A0N(\ram[255][8] ), .A1N(n6355), 
        .Y(n4670) );
  OAI2BB2XL U4391 ( .B0(n6755), .B1(n458), .A0N(\ram[255][9] ), .A1N(n6355), 
        .Y(n4671) );
  OAI2BB2XL U4392 ( .B0(n6732), .B1(n458), .A0N(\ram[255][10] ), .A1N(n6355), 
        .Y(n4672) );
  OAI2BB2XL U4393 ( .B0(n6709), .B1(n458), .A0N(\ram[255][11] ), .A1N(n6355), 
        .Y(n4673) );
  OAI2BB2XL U4394 ( .B0(n6686), .B1(n458), .A0N(\ram[255][12] ), .A1N(n6355), 
        .Y(n4674) );
  OAI2BB2XL U4395 ( .B0(n6663), .B1(n458), .A0N(\ram[255][13] ), .A1N(n6355), 
        .Y(n4675) );
  OAI2BB2XL U4396 ( .B0(n6640), .B1(n458), .A0N(\ram[255][14] ), .A1N(n6355), 
        .Y(n4676) );
  OAI2BB2XL U4397 ( .B0(n6617), .B1(n458), .A0N(\ram[255][15] ), .A1N(n6355), 
        .Y(n4677) );
  CLKINVX3 U4398 ( .A(n6266), .Y(n6269) );
  CLKINVX3 U4399 ( .A(n6266), .Y(n6270) );
  CLKINVX3 U4400 ( .A(n6265), .Y(n6271) );
  CLKINVX3 U4401 ( .A(n6265), .Y(n6272) );
  CLKINVX3 U4402 ( .A(n6264), .Y(n6273) );
  CLKINVX3 U4403 ( .A(n6263), .Y(n6276) );
  CLKINVX3 U4404 ( .A(n6264), .Y(n6274) );
  CLKINVX3 U4405 ( .A(n6263), .Y(n6275) );
  CLKINVX3 U4406 ( .A(n6262), .Y(n6277) );
  CLKINVX3 U4407 ( .A(n6262), .Y(n6278) );
  CLKINVX3 U4408 ( .A(n6260), .Y(n6281) );
  CLKINVX3 U4409 ( .A(n6261), .Y(n6279) );
  CLKINVX3 U4410 ( .A(n6261), .Y(n6280) );
  CLKINVX3 U4411 ( .A(n6260), .Y(n6282) );
  CLKINVX3 U4412 ( .A(n6259), .Y(n6283) );
  CLKINVX3 U4413 ( .A(n6259), .Y(n6284) );
  CLKINVX3 U4414 ( .A(n6257), .Y(n6287) );
  CLKINVX3 U4415 ( .A(n6257), .Y(n6288) );
  CLKINVX3 U4416 ( .A(n6258), .Y(n6285) );
  CLKINVX3 U4417 ( .A(n6258), .Y(n6286) );
  CLKINVX3 U4418 ( .A(n6256), .Y(n6289) );
  CLKINVX3 U4419 ( .A(n6255), .Y(n6292) );
  CLKINVX3 U4420 ( .A(n6256), .Y(n6290) );
  CLKINVX3 U4421 ( .A(n6255), .Y(n6291) );
  CLKINVX3 U4422 ( .A(n6254), .Y(n6293) );
  CLKINVX3 U4423 ( .A(n6254), .Y(n6294) );
  CLKINVX3 U4424 ( .A(n6252), .Y(n6297) );
  CLKINVX3 U4425 ( .A(n6253), .Y(n6295) );
  CLKINVX3 U4426 ( .A(n6253), .Y(n6296) );
  CLKINVX3 U4427 ( .A(n6252), .Y(n6298) );
  CLKINVX3 U4428 ( .A(n6251), .Y(n6299) );
  CLKINVX3 U4429 ( .A(n6251), .Y(n6300) );
  CLKINVX3 U4430 ( .A(n6250), .Y(n6301) );
  CLKINVX3 U4431 ( .A(n6250), .Y(n6302) );
  CLKINVX3 U4432 ( .A(n6249), .Y(n6303) );
  CLKINVX3 U4433 ( .A(n6249), .Y(n6304) );
  CLKINVX3 U4434 ( .A(n6248), .Y(n6305) );
  CLKINVX3 U4435 ( .A(n6247), .Y(n6308) );
  CLKINVX3 U4436 ( .A(n6248), .Y(n6306) );
  CLKINVX3 U4437 ( .A(n6247), .Y(n6307) );
  CLKINVX3 U4438 ( .A(n6246), .Y(n6309) );
  CLKINVX3 U4439 ( .A(n6246), .Y(n6310) );
  CLKINVX3 U4440 ( .A(n6244), .Y(n6313) );
  CLKINVX3 U4441 ( .A(n6245), .Y(n6311) );
  CLKINVX3 U4442 ( .A(n6245), .Y(n6312) );
  CLKINVX3 U4443 ( .A(n6245), .Y(n6314) );
  CLKINVX3 U4444 ( .A(n6244), .Y(n6315) );
  CLKINVX3 U4445 ( .A(n6244), .Y(n6316) );
  CLKINVX3 U4446 ( .A(n6243), .Y(n6317) );
  CLKINVX3 U4447 ( .A(n6243), .Y(n6318) );
  CLKINVX3 U4448 ( .A(n6242), .Y(n6319) );
  CLKINVX3 U4449 ( .A(n6242), .Y(n6320) );
  CLKINVX3 U4450 ( .A(n6243), .Y(n6321) );
  CLKINVX3 U4451 ( .A(n6242), .Y(n6322) );
  CLKINVX3 U4452 ( .A(n6231), .Y(n6268) );
  CLKINVX3 U4453 ( .A(n6241), .Y(n6323) );
  CLKINVX3 U4454 ( .A(n6241), .Y(n6324) );
  CLKINVX3 U4455 ( .A(n6240), .Y(n6325) );
  CLKINVX3 U4456 ( .A(n6240), .Y(n6326) );
  CLKINVX3 U4457 ( .A(n6239), .Y(n6329) );
  CLKINVX3 U4458 ( .A(n6240), .Y(n6327) );
  CLKINVX3 U4459 ( .A(n6241), .Y(n6328) );
  CLKINVX3 U4460 ( .A(n6239), .Y(n6330) );
  CLKINVX3 U4461 ( .A(n6238), .Y(n6331) );
  CLKINVX3 U4462 ( .A(n6238), .Y(n6332) );
  CLKINVX3 U4463 ( .A(n6237), .Y(n6333) );
  CLKINVX3 U4464 ( .A(n6237), .Y(n6334) );
  CLKINVX3 U4465 ( .A(n6236), .Y(n6335) );
  CLKINVX3 U4466 ( .A(n6236), .Y(n6336) );
  CLKINVX3 U4467 ( .A(n6235), .Y(n6337) );
  CLKINVX3 U4468 ( .A(n6234), .Y(n6340) );
  CLKINVX3 U4469 ( .A(n6235), .Y(n6338) );
  CLKINVX3 U4470 ( .A(n6234), .Y(n6339) );
  CLKINVX3 U4471 ( .A(n6233), .Y(n6341) );
  CLKINVX3 U4472 ( .A(n6233), .Y(n6342) );
  CLKINVX3 U4473 ( .A(n6231), .Y(n6345) );
  CLKINVX3 U4474 ( .A(n6232), .Y(n6343) );
  CLKINVX3 U4475 ( .A(n6232), .Y(n6344) );
  CLKINVX3 U4476 ( .A(n6231), .Y(n6346) );
  INVX1 U4477 ( .A(n6217), .Y(n6266) );
  INVX1 U4478 ( .A(n6217), .Y(n6265) );
  INVX1 U4479 ( .A(n6217), .Y(n6264) );
  INVX1 U4480 ( .A(n6218), .Y(n6263) );
  INVX1 U4481 ( .A(n6218), .Y(n6262) );
  INVX1 U4482 ( .A(n6218), .Y(n6261) );
  INVX1 U4483 ( .A(n6219), .Y(n6260) );
  INVX1 U4484 ( .A(n6219), .Y(n6259) );
  INVX1 U4485 ( .A(n6220), .Y(n6257) );
  INVX1 U4486 ( .A(n6219), .Y(n6258) );
  INVX1 U4487 ( .A(n6220), .Y(n6256) );
  INVX1 U4488 ( .A(n6220), .Y(n6255) );
  INVX1 U4489 ( .A(n6221), .Y(n6254) );
  INVX1 U4490 ( .A(n6221), .Y(n6253) );
  INVX1 U4491 ( .A(n6221), .Y(n6252) );
  INVX1 U4492 ( .A(n6222), .Y(n6251) );
  INVX1 U4493 ( .A(n6222), .Y(n6250) );
  INVX1 U4494 ( .A(n6222), .Y(n6249) );
  INVX1 U4495 ( .A(n6223), .Y(n6248) );
  INVX1 U4496 ( .A(n6223), .Y(n6247) );
  INVX1 U4497 ( .A(n6223), .Y(n6246) );
  INVX1 U4498 ( .A(n6223), .Y(n6245) );
  INVX1 U4499 ( .A(n6222), .Y(n6244) );
  INVX1 U4500 ( .A(n6224), .Y(n6243) );
  INVX1 U4501 ( .A(n6224), .Y(n6242) );
  INVX1 U4502 ( .A(n6229), .Y(n6267) );
  CLKINVX3 U4503 ( .A(n6230), .Y(n6347) );
  CLKINVX3 U4504 ( .A(n6230), .Y(n6348) );
  CLKINVX3 U4505 ( .A(n6229), .Y(n6349) );
  CLKINVX3 U4506 ( .A(n6229), .Y(n6350) );
  CLKINVX3 U4507 ( .A(n6228), .Y(n6351) );
  CLKINVX3 U4508 ( .A(n6228), .Y(n6352) );
  INVX1 U4509 ( .A(n6215), .Y(n6217) );
  INVX1 U4510 ( .A(n6215), .Y(n6218) );
  INVX1 U4511 ( .A(n6215), .Y(n6219) );
  INVX1 U4512 ( .A(n6216), .Y(n6220) );
  INVX1 U4513 ( .A(n6216), .Y(n6221) );
  INVX1 U4514 ( .A(n6216), .Y(n6222) );
  INVX1 U4515 ( .A(n6216), .Y(n6223) );
  INVX1 U4516 ( .A(n6216), .Y(n6224) );
  INVX1 U4517 ( .A(n6219), .Y(n6241) );
  INVX1 U4518 ( .A(n6218), .Y(n6240) );
  INVX1 U4519 ( .A(n6225), .Y(n6239) );
  INVX1 U4520 ( .A(n6225), .Y(n6238) );
  INVX1 U4521 ( .A(n6225), .Y(n6237) );
  INVX1 U4522 ( .A(n6226), .Y(n6236) );
  INVX1 U4523 ( .A(n6226), .Y(n6235) );
  INVX1 U4524 ( .A(n6226), .Y(n6234) );
  INVX1 U4525 ( .A(n6227), .Y(n6233) );
  INVX1 U4526 ( .A(n6227), .Y(n6232) );
  INVX1 U4527 ( .A(n6227), .Y(n6231) );
  CLKINVX3 U4528 ( .A(n6132), .Y(n6135) );
  CLKINVX3 U4529 ( .A(n6132), .Y(n6136) );
  CLKINVX3 U4530 ( .A(n6131), .Y(n6137) );
  CLKINVX3 U4531 ( .A(n6131), .Y(n6138) );
  CLKINVX3 U4532 ( .A(n6094), .Y(n6139) );
  CLKINVX3 U4533 ( .A(n6130), .Y(n6142) );
  CLKINVX3 U4534 ( .A(n6094), .Y(n6140) );
  CLKINVX3 U4535 ( .A(n6130), .Y(n6141) );
  CLKINVX3 U4536 ( .A(n6129), .Y(n6143) );
  CLKINVX3 U4537 ( .A(n6129), .Y(n6144) );
  CLKINVX3 U4538 ( .A(n6127), .Y(n6147) );
  CLKINVX3 U4539 ( .A(n6128), .Y(n6145) );
  CLKINVX3 U4540 ( .A(n6128), .Y(n6146) );
  CLKINVX3 U4541 ( .A(n6127), .Y(n6148) );
  CLKINVX3 U4542 ( .A(n6126), .Y(n6149) );
  CLKINVX3 U4543 ( .A(n6126), .Y(n6150) );
  CLKINVX3 U4544 ( .A(n6124), .Y(n6153) );
  CLKINVX3 U4545 ( .A(n6124), .Y(n6154) );
  CLKINVX3 U4546 ( .A(n6125), .Y(n6151) );
  CLKINVX3 U4547 ( .A(n6125), .Y(n6152) );
  CLKINVX3 U4548 ( .A(n6123), .Y(n6155) );
  CLKINVX3 U4549 ( .A(n6122), .Y(n6158) );
  CLKINVX3 U4550 ( .A(n6123), .Y(n6156) );
  CLKINVX3 U4551 ( .A(n6122), .Y(n6157) );
  CLKINVX3 U4552 ( .A(n6121), .Y(n6159) );
  CLKINVX3 U4553 ( .A(n6121), .Y(n6160) );
  CLKINVX3 U4554 ( .A(n6119), .Y(n6163) );
  CLKINVX3 U4555 ( .A(n6120), .Y(n6161) );
  CLKINVX3 U4556 ( .A(n6120), .Y(n6162) );
  CLKINVX3 U4557 ( .A(n6119), .Y(n6164) );
  CLKINVX3 U4558 ( .A(n6118), .Y(n6165) );
  CLKINVX3 U4559 ( .A(n6118), .Y(n6166) );
  CLKINVX3 U4560 ( .A(n6117), .Y(n6167) );
  CLKINVX3 U4561 ( .A(n6117), .Y(n6168) );
  CLKINVX3 U4562 ( .A(n6116), .Y(n6169) );
  CLKINVX3 U4563 ( .A(n6116), .Y(n6170) );
  CLKINVX3 U4564 ( .A(n6115), .Y(n6171) );
  CLKINVX3 U4565 ( .A(n6114), .Y(n6174) );
  CLKINVX3 U4566 ( .A(n6115), .Y(n6172) );
  CLKINVX3 U4567 ( .A(n6114), .Y(n6173) );
  CLKINVX3 U4568 ( .A(n6113), .Y(n6175) );
  CLKINVX3 U4569 ( .A(n6113), .Y(n6176) );
  CLKINVX3 U4570 ( .A(n6111), .Y(n6179) );
  CLKINVX3 U4571 ( .A(n6112), .Y(n6177) );
  CLKINVX3 U4572 ( .A(n6112), .Y(n6178) );
  CLKINVX3 U4573 ( .A(n6111), .Y(n6180) );
  CLKINVX3 U4574 ( .A(n6110), .Y(n6181) );
  CLKINVX3 U4575 ( .A(n6110), .Y(n6182) );
  CLKINVX3 U4576 ( .A(n6109), .Y(n6183) );
  CLKINVX3 U4577 ( .A(n6109), .Y(n6184) );
  CLKINVX3 U4578 ( .A(n6108), .Y(n6185) );
  CLKINVX3 U4579 ( .A(n6108), .Y(n6186) );
  CLKINVX3 U4580 ( .A(n6107), .Y(n6187) );
  CLKINVX3 U4581 ( .A(n6107), .Y(n6188) );
  CLKINVX3 U4582 ( .A(n6054), .Y(n6056) );
  CLKINVX3 U4583 ( .A(n6053), .Y(n6057) );
  CLKINVX3 U4584 ( .A(n6055), .Y(n6058) );
  CLKINVX3 U4585 ( .A(n6055), .Y(n6059) );
  CLKINVX3 U4586 ( .A(n6050), .Y(n6060) );
  CLKINVX3 U4587 ( .A(n7011), .Y(n6061) );
  CLKINVX3 U4588 ( .A(n6055), .Y(n6062) );
  CLKINVX3 U4589 ( .A(n7009), .Y(n6063) );
  CLKINVX3 U4590 ( .A(n6054), .Y(n6064) );
  CLKINVX3 U4591 ( .A(n6054), .Y(n6065) );
  CLKINVX3 U4592 ( .A(n6053), .Y(n6066) );
  CLKINVX3 U4593 ( .A(n6053), .Y(n6067) );
  CLKINVX3 U4594 ( .A(n6052), .Y(n6068) );
  CLKINVX3 U4595 ( .A(n6054), .Y(n6069) );
  CLKINVX3 U4596 ( .A(n6052), .Y(n6070) );
  CLKINVX3 U4597 ( .A(n6052), .Y(n6071) );
  CLKINVX3 U4598 ( .A(n6052), .Y(n6072) );
  CLKINVX3 U4599 ( .A(n7009), .Y(n6073) );
  INVX1 U4600 ( .A(n6215), .Y(n6225) );
  INVX1 U4601 ( .A(n6215), .Y(n6226) );
  INVX1 U4602 ( .A(n6215), .Y(n6227) );
  INVX1 U4603 ( .A(n6354), .Y(n6216) );
  INVX1 U4604 ( .A(n6226), .Y(n6230) );
  INVX1 U4605 ( .A(n6227), .Y(n6229) );
  INVX1 U4606 ( .A(n6226), .Y(n6228) );
  CLKINVX3 U4607 ( .A(n6132), .Y(n6134) );
  CLKINVX3 U4608 ( .A(n6106), .Y(n6189) );
  CLKINVX3 U4609 ( .A(n6106), .Y(n6190) );
  CLKINVX3 U4610 ( .A(n6105), .Y(n6191) );
  CLKINVX3 U4611 ( .A(n6105), .Y(n6192) );
  CLKINVX3 U4612 ( .A(n6103), .Y(n6195) );
  CLKINVX3 U4613 ( .A(n6104), .Y(n6193) );
  CLKINVX3 U4614 ( .A(n6104), .Y(n6194) );
  CLKINVX3 U4615 ( .A(n6103), .Y(n6196) );
  CLKINVX3 U4616 ( .A(n6102), .Y(n6197) );
  CLKINVX3 U4617 ( .A(n6102), .Y(n6198) );
  CLKINVX3 U4618 ( .A(n6101), .Y(n6199) );
  CLKINVX3 U4619 ( .A(n6101), .Y(n6200) );
  CLKINVX3 U4620 ( .A(n6100), .Y(n6201) );
  CLKINVX3 U4621 ( .A(n6100), .Y(n6202) );
  CLKINVX3 U4622 ( .A(n6099), .Y(n6203) );
  CLKINVX3 U4623 ( .A(n6098), .Y(n6206) );
  CLKINVX3 U4624 ( .A(n6099), .Y(n6204) );
  CLKINVX3 U4625 ( .A(n6098), .Y(n6205) );
  CLKINVX3 U4626 ( .A(n6097), .Y(n6207) );
  CLKINVX3 U4627 ( .A(n6097), .Y(n6208) );
  CLKINVX3 U4628 ( .A(n6095), .Y(n6211) );
  CLKINVX3 U4629 ( .A(n6096), .Y(n6209) );
  CLKINVX3 U4630 ( .A(n6096), .Y(n6210) );
  CLKINVX3 U4631 ( .A(n6095), .Y(n6212) );
  INVX1 U4632 ( .A(n6131), .Y(n6133) );
  INVX1 U4633 ( .A(n6082), .Y(n6132) );
  INVX1 U4634 ( .A(n6083), .Y(n6131) );
  INVX1 U4635 ( .A(n6082), .Y(n6130) );
  INVX1 U4636 ( .A(n6082), .Y(n6129) );
  INVX1 U4637 ( .A(n6082), .Y(n6128) );
  INVX1 U4638 ( .A(n6083), .Y(n6127) );
  INVX1 U4639 ( .A(n6083), .Y(n6126) );
  INVX1 U4640 ( .A(n6084), .Y(n6124) );
  INVX1 U4641 ( .A(n6083), .Y(n6125) );
  INVX1 U4642 ( .A(n6084), .Y(n6123) );
  INVX1 U4643 ( .A(n6084), .Y(n6122) );
  INVX1 U4644 ( .A(n6085), .Y(n6121) );
  INVX1 U4645 ( .A(n6085), .Y(n6120) );
  INVX1 U4646 ( .A(n6085), .Y(n6119) );
  INVX1 U4647 ( .A(n6086), .Y(n6118) );
  INVX1 U4648 ( .A(n6086), .Y(n6117) );
  INVX1 U4649 ( .A(n6086), .Y(n6116) );
  INVX1 U4650 ( .A(n6087), .Y(n6115) );
  INVX1 U4651 ( .A(n6087), .Y(n6114) );
  INVX1 U4652 ( .A(n6087), .Y(n6113) );
  INVX1 U4653 ( .A(n6088), .Y(n6112) );
  INVX1 U4654 ( .A(n6088), .Y(n6111) );
  INVX1 U4655 ( .A(n6088), .Y(n6110) );
  INVX1 U4656 ( .A(n6089), .Y(n6109) );
  INVX1 U4657 ( .A(n6089), .Y(n6108) );
  INVX1 U4658 ( .A(n6089), .Y(n6107) );
  INVX1 U4659 ( .A(n6051), .Y(n6055) );
  INVX1 U4660 ( .A(n6051), .Y(n6054) );
  INVX1 U4661 ( .A(n6051), .Y(n6053) );
  INVX1 U4662 ( .A(n6051), .Y(n6052) );
  INVX1 U4663 ( .A(n6354), .Y(n6215) );
  CLKINVX3 U4664 ( .A(n6024), .Y(n6033) );
  CLKINVX3 U4665 ( .A(n6024), .Y(n6034) );
  CLKINVX3 U4666 ( .A(n6024), .Y(n6035) );
  CLKINVX3 U4667 ( .A(n6032), .Y(n6036) );
  CLKINVX3 U4668 ( .A(n6032), .Y(n6037) );
  CLKINVX3 U4669 ( .A(n6031), .Y(n6038) );
  CLKINVX3 U4670 ( .A(n6031), .Y(n6039) );
  CLKINVX3 U4671 ( .A(n6030), .Y(n6040) );
  CLKINVX3 U4672 ( .A(n6030), .Y(n6041) );
  CLKINVX3 U4673 ( .A(n6029), .Y(n6042) );
  CLKINVX3 U4674 ( .A(n6029), .Y(n6043) );
  CLKINVX3 U4675 ( .A(n6028), .Y(n6044) );
  CLKINVX3 U4676 ( .A(n6028), .Y(n6045) );
  CLKINVX3 U4677 ( .A(n6027), .Y(n6046) );
  CLKINVX3 U4678 ( .A(n6027), .Y(n6047) );
  CLKINVX3 U4679 ( .A(n6094), .Y(n6213) );
  CLKINVX3 U4680 ( .A(n6094), .Y(n6214) );
  INVX1 U4681 ( .A(n6081), .Y(n6082) );
  INVX1 U4682 ( .A(n6081), .Y(n6083) );
  INVX1 U4683 ( .A(n6080), .Y(n6084) );
  INVX1 U4684 ( .A(n6080), .Y(n6085) );
  INVX1 U4685 ( .A(n6079), .Y(n6086) );
  INVX1 U4686 ( .A(n6079), .Y(n6087) );
  INVX1 U4687 ( .A(n6079), .Y(n6088) );
  INVX1 U4688 ( .A(n6080), .Y(n6089) );
  INVX1 U4689 ( .A(n6050), .Y(n6051) );
  INVX1 U4690 ( .A(n6090), .Y(n6106) );
  INVX1 U4691 ( .A(n6090), .Y(n6105) );
  INVX1 U4692 ( .A(n6090), .Y(n6104) );
  INVX1 U4693 ( .A(n6091), .Y(n6103) );
  INVX1 U4694 ( .A(n6091), .Y(n6102) );
  INVX1 U4695 ( .A(n6091), .Y(n6101) );
  INVX1 U4696 ( .A(n6092), .Y(n6100) );
  INVX1 U4697 ( .A(n6092), .Y(n6099) );
  INVX1 U4698 ( .A(n6092), .Y(n6098) );
  INVX1 U4699 ( .A(n6093), .Y(n6097) );
  INVX1 U4700 ( .A(n6093), .Y(n6096) );
  INVX1 U4701 ( .A(n6093), .Y(n6095) );
  CLKINVX3 U4702 ( .A(n7014), .Y(n6021) );
  CLKINVX3 U4703 ( .A(n7014), .Y(n6022) );
  CLKINVX3 U4704 ( .A(n7014), .Y(n6023) );
  INVX1 U4705 ( .A(n6078), .Y(n6090) );
  INVX1 U4706 ( .A(n6078), .Y(n6091) );
  INVX1 U4707 ( .A(n6077), .Y(n6092) );
  INVX1 U4708 ( .A(n6077), .Y(n6093) );
  INVX1 U4709 ( .A(n6075), .Y(n6081) );
  INVX1 U4710 ( .A(n7010), .Y(n6050) );
  INVX1 U4711 ( .A(n6075), .Y(n6080) );
  INVX1 U4712 ( .A(n6075), .Y(n6079) );
  INVX1 U4713 ( .A(n6076), .Y(n6094) );
  INVX1 U4714 ( .A(n6025), .Y(n6032) );
  INVX1 U4715 ( .A(n6025), .Y(n6031) );
  INVX1 U4716 ( .A(n6025), .Y(n6030) );
  INVX1 U4717 ( .A(n6026), .Y(n6029) );
  INVX1 U4718 ( .A(n6026), .Y(n6028) );
  INVX1 U4719 ( .A(n6026), .Y(n6027) );
  CLKINVX3 U4720 ( .A(n6994), .Y(n6989) );
  CLKINVX3 U4721 ( .A(n6994), .Y(n6988) );
  CLKINVX3 U4722 ( .A(n6995), .Y(n6987) );
  CLKINVX3 U4723 ( .A(n6995), .Y(n6986) );
  CLKINVX3 U4724 ( .A(n6996), .Y(n6984) );
  CLKINVX3 U4725 ( .A(n6996), .Y(n6983) );
  CLKINVX3 U4726 ( .A(n6997), .Y(n6982) );
  CLKINVX3 U4727 ( .A(n6997), .Y(n6981) );
  CLKINVX3 U4728 ( .A(n6995), .Y(n6985) );
  CLKINVX3 U4729 ( .A(n6994), .Y(n6990) );
  CLKINVX3 U4730 ( .A(n6993), .Y(n6991) );
  CLKINVX3 U4731 ( .A(n6993), .Y(n6992) );
  INVX1 U4732 ( .A(n6353), .Y(n6354) );
  INVX1 U4733 ( .A(n7004), .Y(n6353) );
  INVX1 U4734 ( .A(n6074), .Y(n6075) );
  INVX1 U4735 ( .A(n6024), .Y(n6025) );
  INVX1 U4736 ( .A(n6024), .Y(n6026) );
  INVX1 U4737 ( .A(n6076), .Y(n6078) );
  INVX1 U4738 ( .A(n6076), .Y(n6077) );
  CLKINVX3 U4739 ( .A(n7016), .Y(n6017) );
  CLKINVX3 U4740 ( .A(n7016), .Y(n6018) );
  CLKINVX3 U4741 ( .A(n7016), .Y(n6019) );
  CLKINVX3 U4742 ( .A(n7016), .Y(n6020) );
  CLKINVX3 U4743 ( .A(n6883), .Y(n6882) );
  CLKINVX3 U4744 ( .A(n6860), .Y(n6859) );
  CLKINVX3 U4745 ( .A(n6837), .Y(n6836) );
  CLKINVX3 U4746 ( .A(n6814), .Y(n6813) );
  CLKINVX3 U4747 ( .A(n6791), .Y(n6790) );
  CLKINVX3 U4748 ( .A(n6768), .Y(n6767) );
  CLKINVX3 U4749 ( .A(n6745), .Y(n6744) );
  CLKINVX3 U4750 ( .A(n6722), .Y(n6721) );
  CLKINVX3 U4751 ( .A(n6699), .Y(n6698) );
  CLKINVX3 U4752 ( .A(n6676), .Y(n6675) );
  CLKINVX3 U4753 ( .A(n6653), .Y(n6652) );
  CLKINVX3 U4754 ( .A(n6630), .Y(n6629) );
  CLKINVX3 U4755 ( .A(n6883), .Y(n6881) );
  CLKINVX3 U4756 ( .A(n6860), .Y(n6858) );
  CLKINVX3 U4757 ( .A(n6837), .Y(n6835) );
  CLKINVX3 U4758 ( .A(n6814), .Y(n6812) );
  CLKINVX3 U4759 ( .A(n6791), .Y(n6789) );
  CLKINVX3 U4760 ( .A(n6768), .Y(n6766) );
  CLKINVX3 U4761 ( .A(n6745), .Y(n6743) );
  CLKINVX3 U4762 ( .A(n6722), .Y(n6720) );
  CLKINVX3 U4763 ( .A(n6699), .Y(n6697) );
  CLKINVX3 U4764 ( .A(n6676), .Y(n6674) );
  CLKINVX3 U4765 ( .A(n6653), .Y(n6651) );
  CLKINVX3 U4766 ( .A(n6630), .Y(n6628) );
  CLKINVX3 U4767 ( .A(n6883), .Y(n6880) );
  CLKINVX3 U4768 ( .A(n6860), .Y(n6857) );
  CLKINVX3 U4769 ( .A(n6837), .Y(n6834) );
  CLKINVX3 U4770 ( .A(n6814), .Y(n6811) );
  CLKINVX3 U4771 ( .A(n6791), .Y(n6788) );
  CLKINVX3 U4772 ( .A(n6768), .Y(n6765) );
  CLKINVX3 U4773 ( .A(n6745), .Y(n6742) );
  CLKINVX3 U4774 ( .A(n6722), .Y(n6719) );
  CLKINVX3 U4775 ( .A(n6699), .Y(n6696) );
  CLKINVX3 U4776 ( .A(n6676), .Y(n6673) );
  CLKINVX3 U4777 ( .A(n6653), .Y(n6650) );
  CLKINVX3 U4778 ( .A(n6630), .Y(n6627) );
  CLKINVX3 U4779 ( .A(n6883), .Y(n6879) );
  CLKINVX3 U4780 ( .A(n6860), .Y(n6856) );
  CLKINVX3 U4781 ( .A(n6837), .Y(n6833) );
  CLKINVX3 U4782 ( .A(n6814), .Y(n6810) );
  CLKINVX3 U4783 ( .A(n6791), .Y(n6787) );
  CLKINVX3 U4784 ( .A(n6768), .Y(n6764) );
  CLKINVX3 U4785 ( .A(n6745), .Y(n6741) );
  CLKINVX3 U4786 ( .A(n6722), .Y(n6718) );
  CLKINVX3 U4787 ( .A(n6699), .Y(n6695) );
  CLKINVX3 U4788 ( .A(n6676), .Y(n6672) );
  CLKINVX3 U4789 ( .A(n6653), .Y(n6649) );
  CLKINVX3 U4790 ( .A(n6630), .Y(n6626) );
  CLKINVX3 U4791 ( .A(n6884), .Y(n6878) );
  CLKINVX3 U4792 ( .A(n6861), .Y(n6855) );
  CLKINVX3 U4793 ( .A(n6838), .Y(n6832) );
  CLKINVX3 U4794 ( .A(n6815), .Y(n6809) );
  CLKINVX3 U4795 ( .A(n6792), .Y(n6786) );
  CLKINVX3 U4796 ( .A(n6769), .Y(n6763) );
  CLKINVX3 U4797 ( .A(n6746), .Y(n6740) );
  CLKINVX3 U4798 ( .A(n6723), .Y(n6717) );
  CLKINVX3 U4799 ( .A(n6700), .Y(n6694) );
  CLKINVX3 U4800 ( .A(n6677), .Y(n6671) );
  CLKINVX3 U4801 ( .A(n6654), .Y(n6648) );
  CLKINVX3 U4802 ( .A(n6631), .Y(n6625) );
  CLKINVX3 U4803 ( .A(n6975), .Y(n6974) );
  CLKINVX3 U4804 ( .A(n6952), .Y(n6951) );
  CLKINVX3 U4805 ( .A(n6929), .Y(n6928) );
  CLKINVX3 U4806 ( .A(n6906), .Y(n6905) );
  CLKINVX3 U4807 ( .A(n6884), .Y(n6877) );
  CLKINVX3 U4808 ( .A(n6861), .Y(n6854) );
  CLKINVX3 U4809 ( .A(n6838), .Y(n6831) );
  CLKINVX3 U4810 ( .A(n6815), .Y(n6808) );
  CLKINVX3 U4811 ( .A(n6792), .Y(n6785) );
  CLKINVX3 U4812 ( .A(n6769), .Y(n6762) );
  CLKINVX3 U4813 ( .A(n6746), .Y(n6739) );
  CLKINVX3 U4814 ( .A(n6723), .Y(n6716) );
  CLKINVX3 U4815 ( .A(n6700), .Y(n6693) );
  CLKINVX3 U4816 ( .A(n6677), .Y(n6670) );
  CLKINVX3 U4817 ( .A(n6654), .Y(n6647) );
  CLKINVX3 U4818 ( .A(n6631), .Y(n6624) );
  CLKINVX3 U4819 ( .A(n6975), .Y(n6973) );
  CLKINVX3 U4820 ( .A(n6952), .Y(n6950) );
  CLKINVX3 U4821 ( .A(n6929), .Y(n6927) );
  CLKINVX3 U4822 ( .A(n6906), .Y(n6904) );
  CLKINVX3 U4823 ( .A(n6884), .Y(n6876) );
  CLKINVX3 U4824 ( .A(n6861), .Y(n6853) );
  CLKINVX3 U4825 ( .A(n6838), .Y(n6830) );
  CLKINVX3 U4826 ( .A(n6815), .Y(n6807) );
  CLKINVX3 U4827 ( .A(n6792), .Y(n6784) );
  CLKINVX3 U4828 ( .A(n6769), .Y(n6761) );
  CLKINVX3 U4829 ( .A(n6746), .Y(n6738) );
  CLKINVX3 U4830 ( .A(n6723), .Y(n6715) );
  CLKINVX3 U4831 ( .A(n6700), .Y(n6692) );
  CLKINVX3 U4832 ( .A(n6677), .Y(n6669) );
  CLKINVX3 U4833 ( .A(n6654), .Y(n6646) );
  CLKINVX3 U4834 ( .A(n6631), .Y(n6623) );
  CLKINVX3 U4835 ( .A(n6976), .Y(n6972) );
  CLKINVX3 U4836 ( .A(n6953), .Y(n6949) );
  CLKINVX3 U4837 ( .A(n6930), .Y(n6926) );
  CLKINVX3 U4838 ( .A(n6907), .Y(n6903) );
  CLKINVX3 U4839 ( .A(n6884), .Y(n6875) );
  CLKINVX3 U4840 ( .A(n6861), .Y(n6852) );
  CLKINVX3 U4841 ( .A(n6838), .Y(n6829) );
  CLKINVX3 U4842 ( .A(n6815), .Y(n6806) );
  CLKINVX3 U4843 ( .A(n6792), .Y(n6783) );
  CLKINVX3 U4844 ( .A(n6769), .Y(n6760) );
  CLKINVX3 U4845 ( .A(n6746), .Y(n6737) );
  CLKINVX3 U4846 ( .A(n6723), .Y(n6714) );
  CLKINVX3 U4847 ( .A(n6700), .Y(n6691) );
  CLKINVX3 U4848 ( .A(n6677), .Y(n6668) );
  CLKINVX3 U4849 ( .A(n6654), .Y(n6645) );
  CLKINVX3 U4850 ( .A(n6631), .Y(n6622) );
  CLKINVX3 U4851 ( .A(n6976), .Y(n6971) );
  CLKINVX3 U4852 ( .A(n6953), .Y(n6948) );
  CLKINVX3 U4853 ( .A(n6930), .Y(n6925) );
  CLKINVX3 U4854 ( .A(n6907), .Y(n6902) );
  CLKINVX3 U4855 ( .A(n6883), .Y(n6874) );
  CLKINVX3 U4856 ( .A(n6860), .Y(n6851) );
  CLKINVX3 U4857 ( .A(n6837), .Y(n6828) );
  CLKINVX3 U4858 ( .A(n6814), .Y(n6805) );
  CLKINVX3 U4859 ( .A(n6791), .Y(n6782) );
  CLKINVX3 U4860 ( .A(n6768), .Y(n6759) );
  CLKINVX3 U4861 ( .A(n6745), .Y(n6736) );
  CLKINVX3 U4862 ( .A(n6722), .Y(n6713) );
  CLKINVX3 U4863 ( .A(n6699), .Y(n6690) );
  CLKINVX3 U4864 ( .A(n6676), .Y(n6667) );
  CLKINVX3 U4865 ( .A(n6653), .Y(n6644) );
  CLKINVX3 U4866 ( .A(n6630), .Y(n6621) );
  CLKINVX3 U4867 ( .A(n6975), .Y(n6970) );
  CLKINVX3 U4868 ( .A(n6952), .Y(n6947) );
  CLKINVX3 U4869 ( .A(n6929), .Y(n6924) );
  CLKINVX3 U4870 ( .A(n6906), .Y(n6901) );
  CLKINVX3 U4871 ( .A(n6884), .Y(n6873) );
  CLKINVX3 U4872 ( .A(n6861), .Y(n6850) );
  CLKINVX3 U4873 ( .A(n6838), .Y(n6827) );
  CLKINVX3 U4874 ( .A(n6815), .Y(n6804) );
  CLKINVX3 U4875 ( .A(n6792), .Y(n6781) );
  CLKINVX3 U4876 ( .A(n6769), .Y(n6758) );
  CLKINVX3 U4877 ( .A(n6746), .Y(n6735) );
  CLKINVX3 U4878 ( .A(n6723), .Y(n6712) );
  CLKINVX3 U4879 ( .A(n6700), .Y(n6689) );
  CLKINVX3 U4880 ( .A(n6677), .Y(n6666) );
  CLKINVX3 U4881 ( .A(n6654), .Y(n6643) );
  CLKINVX3 U4882 ( .A(n6631), .Y(n6620) );
  CLKINVX3 U4883 ( .A(n6976), .Y(n6969) );
  CLKINVX3 U4884 ( .A(n6953), .Y(n6946) );
  CLKINVX3 U4885 ( .A(n6930), .Y(n6923) );
  CLKINVX3 U4886 ( .A(n6907), .Y(n6900) );
  CLKINVX3 U4887 ( .A(n6886), .Y(n6872) );
  CLKINVX3 U4888 ( .A(n6863), .Y(n6849) );
  CLKINVX3 U4889 ( .A(n6840), .Y(n6826) );
  CLKINVX3 U4890 ( .A(n6817), .Y(n6803) );
  CLKINVX3 U4891 ( .A(n6794), .Y(n6780) );
  CLKINVX3 U4892 ( .A(n6771), .Y(n6757) );
  CLKINVX3 U4893 ( .A(n6748), .Y(n6734) );
  CLKINVX3 U4894 ( .A(n6725), .Y(n6711) );
  CLKINVX3 U4895 ( .A(n6702), .Y(n6688) );
  CLKINVX3 U4896 ( .A(n6679), .Y(n6665) );
  CLKINVX3 U4897 ( .A(n6656), .Y(n6642) );
  CLKINVX3 U4898 ( .A(n6633), .Y(n6619) );
  CLKINVX3 U4899 ( .A(n6977), .Y(n6968) );
  CLKINVX3 U4900 ( .A(n6954), .Y(n6945) );
  CLKINVX3 U4901 ( .A(n6931), .Y(n6922) );
  CLKINVX3 U4902 ( .A(n6908), .Y(n6899) );
  CLKINVX3 U4903 ( .A(n6885), .Y(n6871) );
  CLKINVX3 U4904 ( .A(n6862), .Y(n6848) );
  CLKINVX3 U4905 ( .A(n6839), .Y(n6825) );
  CLKINVX3 U4906 ( .A(n6816), .Y(n6802) );
  CLKINVX3 U4907 ( .A(n6793), .Y(n6779) );
  CLKINVX3 U4908 ( .A(n6770), .Y(n6756) );
  CLKINVX3 U4909 ( .A(n6747), .Y(n6733) );
  CLKINVX3 U4910 ( .A(n6724), .Y(n6710) );
  CLKINVX3 U4911 ( .A(n6701), .Y(n6687) );
  CLKINVX3 U4912 ( .A(n6678), .Y(n6664) );
  CLKINVX3 U4913 ( .A(n6655), .Y(n6641) );
  CLKINVX3 U4914 ( .A(n6632), .Y(n6618) );
  CLKINVX3 U4915 ( .A(n6977), .Y(n6967) );
  CLKINVX3 U4916 ( .A(n6954), .Y(n6944) );
  CLKINVX3 U4917 ( .A(n6931), .Y(n6921) );
  CLKINVX3 U4918 ( .A(n6908), .Y(n6898) );
  CLKINVX3 U4919 ( .A(n6885), .Y(n6870) );
  CLKINVX3 U4920 ( .A(n6862), .Y(n6847) );
  CLKINVX3 U4921 ( .A(n6839), .Y(n6824) );
  CLKINVX3 U4922 ( .A(n6816), .Y(n6801) );
  CLKINVX3 U4923 ( .A(n6793), .Y(n6778) );
  CLKINVX3 U4924 ( .A(n6770), .Y(n6755) );
  CLKINVX3 U4925 ( .A(n6747), .Y(n6732) );
  CLKINVX3 U4926 ( .A(n6724), .Y(n6709) );
  CLKINVX3 U4927 ( .A(n6701), .Y(n6686) );
  CLKINVX3 U4928 ( .A(n6678), .Y(n6663) );
  CLKINVX3 U4929 ( .A(n6655), .Y(n6640) );
  CLKINVX3 U4930 ( .A(n6632), .Y(n6617) );
  CLKINVX3 U4931 ( .A(n6978), .Y(n6966) );
  CLKINVX3 U4932 ( .A(n6955), .Y(n6943) );
  CLKINVX3 U4933 ( .A(n6932), .Y(n6920) );
  CLKINVX3 U4934 ( .A(n6909), .Y(n6897) );
  CLKINVX3 U4935 ( .A(n6886), .Y(n6869) );
  CLKINVX3 U4936 ( .A(n6863), .Y(n6846) );
  CLKINVX3 U4937 ( .A(n6840), .Y(n6823) );
  CLKINVX3 U4938 ( .A(n6817), .Y(n6800) );
  CLKINVX3 U4939 ( .A(n6794), .Y(n6777) );
  CLKINVX3 U4940 ( .A(n6771), .Y(n6754) );
  CLKINVX3 U4941 ( .A(n6748), .Y(n6731) );
  CLKINVX3 U4942 ( .A(n6725), .Y(n6708) );
  CLKINVX3 U4943 ( .A(n6702), .Y(n6685) );
  CLKINVX3 U4944 ( .A(n6679), .Y(n6662) );
  CLKINVX3 U4945 ( .A(n6656), .Y(n6639) );
  CLKINVX3 U4946 ( .A(n6633), .Y(n6616) );
  CLKINVX3 U4947 ( .A(n6978), .Y(n6965) );
  CLKINVX3 U4948 ( .A(n6955), .Y(n6942) );
  CLKINVX3 U4949 ( .A(n6932), .Y(n6919) );
  CLKINVX3 U4950 ( .A(n6909), .Y(n6896) );
  CLKINVX3 U4951 ( .A(n6977), .Y(n6964) );
  CLKINVX3 U4952 ( .A(n6954), .Y(n6941) );
  CLKINVX3 U4953 ( .A(n6931), .Y(n6918) );
  CLKINVX3 U4954 ( .A(n6908), .Y(n6895) );
  CLKINVX3 U4955 ( .A(n6886), .Y(n6868) );
  CLKINVX3 U4956 ( .A(n6863), .Y(n6845) );
  CLKINVX3 U4957 ( .A(n6840), .Y(n6822) );
  CLKINVX3 U4958 ( .A(n6817), .Y(n6799) );
  CLKINVX3 U4959 ( .A(n6794), .Y(n6776) );
  CLKINVX3 U4960 ( .A(n6771), .Y(n6753) );
  CLKINVX3 U4961 ( .A(n6748), .Y(n6730) );
  CLKINVX3 U4962 ( .A(n6725), .Y(n6707) );
  CLKINVX3 U4963 ( .A(n6702), .Y(n6684) );
  CLKINVX3 U4964 ( .A(n6679), .Y(n6661) );
  CLKINVX3 U4965 ( .A(n6656), .Y(n6638) );
  CLKINVX3 U4966 ( .A(n6633), .Y(n6615) );
  CLKINVX3 U4967 ( .A(n6978), .Y(n6963) );
  CLKINVX3 U4968 ( .A(n6955), .Y(n6940) );
  CLKINVX3 U4969 ( .A(n6932), .Y(n6917) );
  CLKINVX3 U4970 ( .A(n6909), .Y(n6894) );
  CLKINVX3 U4971 ( .A(n6886), .Y(n6867) );
  CLKINVX3 U4972 ( .A(n6863), .Y(n6844) );
  CLKINVX3 U4973 ( .A(n6840), .Y(n6821) );
  CLKINVX3 U4974 ( .A(n6817), .Y(n6798) );
  CLKINVX3 U4975 ( .A(n6794), .Y(n6775) );
  CLKINVX3 U4976 ( .A(n6771), .Y(n6752) );
  CLKINVX3 U4977 ( .A(n6748), .Y(n6729) );
  CLKINVX3 U4978 ( .A(n6725), .Y(n6706) );
  CLKINVX3 U4979 ( .A(n6702), .Y(n6683) );
  CLKINVX3 U4980 ( .A(n6679), .Y(n6660) );
  CLKINVX3 U4981 ( .A(n6656), .Y(n6637) );
  CLKINVX3 U4982 ( .A(n6633), .Y(n6614) );
  CLKINVX3 U4983 ( .A(n6977), .Y(n6962) );
  CLKINVX3 U4984 ( .A(n6954), .Y(n6939) );
  CLKINVX3 U4985 ( .A(n6931), .Y(n6916) );
  CLKINVX3 U4986 ( .A(n6908), .Y(n6893) );
  CLKINVX3 U4987 ( .A(n6978), .Y(n6961) );
  CLKINVX3 U4988 ( .A(n6955), .Y(n6938) );
  CLKINVX3 U4989 ( .A(n6932), .Y(n6915) );
  CLKINVX3 U4990 ( .A(n6909), .Y(n6892) );
  CLKINVX3 U4991 ( .A(n6885), .Y(n6866) );
  CLKINVX3 U4992 ( .A(n6862), .Y(n6843) );
  CLKINVX3 U4993 ( .A(n6839), .Y(n6820) );
  CLKINVX3 U4994 ( .A(n6816), .Y(n6797) );
  CLKINVX3 U4995 ( .A(n6793), .Y(n6774) );
  CLKINVX3 U4996 ( .A(n6770), .Y(n6751) );
  CLKINVX3 U4997 ( .A(n6747), .Y(n6728) );
  CLKINVX3 U4998 ( .A(n6724), .Y(n6705) );
  CLKINVX3 U4999 ( .A(n6701), .Y(n6682) );
  CLKINVX3 U5000 ( .A(n6678), .Y(n6659) );
  CLKINVX3 U5001 ( .A(n6655), .Y(n6636) );
  CLKINVX3 U5002 ( .A(n6632), .Y(n6613) );
  CLKINVX3 U5003 ( .A(n6975), .Y(n6960) );
  CLKINVX3 U5004 ( .A(n6952), .Y(n6937) );
  CLKINVX3 U5005 ( .A(n6929), .Y(n6914) );
  CLKINVX3 U5006 ( .A(n6906), .Y(n6891) );
  CLKINVX3 U5007 ( .A(n6885), .Y(n6865) );
  CLKINVX3 U5008 ( .A(n6862), .Y(n6842) );
  CLKINVX3 U5009 ( .A(n6839), .Y(n6819) );
  CLKINVX3 U5010 ( .A(n6816), .Y(n6796) );
  CLKINVX3 U5011 ( .A(n6793), .Y(n6773) );
  CLKINVX3 U5012 ( .A(n6770), .Y(n6750) );
  CLKINVX3 U5013 ( .A(n6747), .Y(n6727) );
  CLKINVX3 U5014 ( .A(n6724), .Y(n6704) );
  CLKINVX3 U5015 ( .A(n6701), .Y(n6681) );
  CLKINVX3 U5016 ( .A(n6678), .Y(n6658) );
  CLKINVX3 U5017 ( .A(n6655), .Y(n6635) );
  CLKINVX3 U5018 ( .A(n6632), .Y(n6612) );
  CLKINVX3 U5019 ( .A(n6976), .Y(n6959) );
  CLKINVX3 U5020 ( .A(n6953), .Y(n6936) );
  CLKINVX3 U5021 ( .A(n6930), .Y(n6913) );
  CLKINVX3 U5022 ( .A(n6907), .Y(n6890) );
  INVX1 U5023 ( .A(n7000), .Y(n6993) );
  INVX1 U5024 ( .A(n6998), .Y(n6996) );
  INVX1 U5025 ( .A(n6998), .Y(n6997) );
  INVX1 U5026 ( .A(n6999), .Y(n6995) );
  INVX1 U5027 ( .A(n6999), .Y(n6994) );
  INVX1 U5028 ( .A(n7005), .Y(n7004) );
  BUFX3 U5029 ( .A(n8), .Y(n6610) );
  NAND2BX1 U5030 ( .AN(n21), .B(n6990), .Y(n8) );
  BUFX3 U5031 ( .A(n27), .Y(n6609) );
  NAND2BXL U5032 ( .AN(n18), .B(n6990), .Y(n27) );
  BUFX3 U5033 ( .A(n30), .Y(n6608) );
  NAND2BXL U5034 ( .AN(n19), .B(n6990), .Y(n30) );
  BUFX3 U5035 ( .A(n33), .Y(n6607) );
  NAND2BXL U5036 ( .AN(n20), .B(n6990), .Y(n33) );
  BUFX3 U5037 ( .A(n36), .Y(n6606) );
  NAND2BXL U5038 ( .AN(n40), .B(n6990), .Y(n36) );
  BUFX3 U5039 ( .A(n39), .Y(n6605) );
  NAND2BXL U5040 ( .AN(n41), .B(n6990), .Y(n39) );
  BUFX3 U5041 ( .A(n42), .Y(n6604) );
  NAND2BXL U5042 ( .AN(n43), .B(n6990), .Y(n42) );
  BUFX3 U5043 ( .A(n45), .Y(n6603) );
  NAND2BXL U5044 ( .AN(n44), .B(n6989), .Y(n45) );
  BUFX3 U5045 ( .A(n48), .Y(n6602) );
  NAND2BXL U5046 ( .AN(n46), .B(n6989), .Y(n48) );
  BUFX3 U5047 ( .A(n51), .Y(n6601) );
  NAND2BXL U5048 ( .AN(n47), .B(n6989), .Y(n51) );
  BUFX3 U5049 ( .A(n54), .Y(n6600) );
  NAND2BXL U5050 ( .AN(n49), .B(n6989), .Y(n54) );
  BUFX3 U5051 ( .A(n57), .Y(n6599) );
  NAND2BXL U5052 ( .AN(n50), .B(n6989), .Y(n57) );
  BUFX3 U5053 ( .A(n60), .Y(n6598) );
  NAND2BXL U5054 ( .AN(n52), .B(n6989), .Y(n60) );
  BUFX3 U5055 ( .A(n63), .Y(n6597) );
  NAND2BXL U5056 ( .AN(n53), .B(n6989), .Y(n63) );
  BUFX3 U5057 ( .A(n66), .Y(n6596) );
  NAND2BXL U5058 ( .AN(n494), .B(n6989), .Y(n66) );
  BUFX3 U5059 ( .A(n69), .Y(n6595) );
  NAND2BXL U5060 ( .AN(n55), .B(n6989), .Y(n69) );
  BUFX3 U5061 ( .A(n74), .Y(n6594) );
  NAND2BXL U5062 ( .AN(n56), .B(n6989), .Y(n74) );
  BUFX3 U5063 ( .A(n77), .Y(n6593) );
  NAND2BXL U5064 ( .AN(n58), .B(n6989), .Y(n77) );
  BUFX3 U5065 ( .A(n79), .Y(n6592) );
  NAND2BXL U5066 ( .AN(n59), .B(n6989), .Y(n79) );
  BUFX3 U5067 ( .A(n81), .Y(n6591) );
  NAND2BXL U5068 ( .AN(n61), .B(n6989), .Y(n81) );
  BUFX3 U5069 ( .A(n83), .Y(n6590) );
  NAND2BXL U5070 ( .AN(n62), .B(n6988), .Y(n83) );
  BUFX3 U5071 ( .A(n85), .Y(n6589) );
  NAND2BXL U5072 ( .AN(n64), .B(n6988), .Y(n85) );
  BUFX3 U5073 ( .A(n87), .Y(n6588) );
  NAND2BXL U5074 ( .AN(n65), .B(n6988), .Y(n87) );
  BUFX3 U5075 ( .A(n89), .Y(n6587) );
  NAND2BXL U5076 ( .AN(n67), .B(n6988), .Y(n89) );
  BUFX3 U5077 ( .A(n91), .Y(n6586) );
  NAND2BXL U5078 ( .AN(n68), .B(n6988), .Y(n91) );
  BUFX3 U5079 ( .A(n93), .Y(n6585) );
  NAND2BXL U5080 ( .AN(n70), .B(n6988), .Y(n93) );
  BUFX3 U5081 ( .A(n95), .Y(n6584) );
  NAND2BXL U5082 ( .AN(n73), .B(n6988), .Y(n95) );
  BUFX3 U5083 ( .A(n97), .Y(n6583) );
  NAND2BXL U5084 ( .AN(n75), .B(n6988), .Y(n97) );
  BUFX3 U5085 ( .A(n99), .Y(n6582) );
  NAND2BXL U5086 ( .AN(n76), .B(n6988), .Y(n99) );
  BUFX3 U5087 ( .A(n101), .Y(n6581) );
  NAND2BXL U5088 ( .AN(n541), .B(n6988), .Y(n101) );
  BUFX3 U5089 ( .A(n103), .Y(n6580) );
  NAND2BXL U5090 ( .AN(n543), .B(n6988), .Y(n103) );
  BUFX3 U5091 ( .A(n105), .Y(n6579) );
  NAND2BXL U5092 ( .AN(n546), .B(n6988), .Y(n105) );
  BUFX3 U5093 ( .A(n108), .Y(n6578) );
  NAND2BXL U5094 ( .AN(n78), .B(n6988), .Y(n108) );
  BUFX3 U5095 ( .A(n111), .Y(n6577) );
  NAND2BXL U5096 ( .AN(n80), .B(n6987), .Y(n111) );
  BUFX3 U5097 ( .A(n113), .Y(n6576) );
  NAND2BXL U5098 ( .AN(n82), .B(n6987), .Y(n113) );
  BUFX3 U5099 ( .A(n115), .Y(n6575) );
  NAND2BXL U5100 ( .AN(n84), .B(n6987), .Y(n115) );
  BUFX3 U5101 ( .A(n117), .Y(n6574) );
  NAND2BXL U5102 ( .AN(n86), .B(n6987), .Y(n117) );
  BUFX3 U5103 ( .A(n119), .Y(n6573) );
  NAND2BXL U5104 ( .AN(n88), .B(n6987), .Y(n119) );
  BUFX3 U5105 ( .A(n121), .Y(n6572) );
  NAND2BXL U5106 ( .AN(n90), .B(n6987), .Y(n121) );
  BUFX3 U5107 ( .A(n123), .Y(n6571) );
  NAND2BXL U5108 ( .AN(n92), .B(n6987), .Y(n123) );
  BUFX3 U5109 ( .A(n125), .Y(n6570) );
  NAND2BXL U5110 ( .AN(n94), .B(n6987), .Y(n125) );
  BUFX3 U5111 ( .A(n127), .Y(n6569) );
  NAND2BXL U5112 ( .AN(n96), .B(n6987), .Y(n127) );
  BUFX3 U5113 ( .A(n131), .Y(n6567) );
  NAND2BXL U5114 ( .AN(n98), .B(n6987), .Y(n131) );
  BUFX3 U5115 ( .A(n133), .Y(n6566) );
  NAND2BXL U5116 ( .AN(n100), .B(n6987), .Y(n133) );
  BUFX3 U5117 ( .A(n135), .Y(n6565) );
  NAND2BXL U5118 ( .AN(n102), .B(n6987), .Y(n135) );
  BUFX3 U5119 ( .A(n137), .Y(n6564) );
  NAND2BXL U5120 ( .AN(n496), .B(n6986), .Y(n137) );
  BUFX3 U5121 ( .A(n139), .Y(n6563) );
  NAND2BXL U5122 ( .AN(n104), .B(n6986), .Y(n139) );
  BUFX3 U5123 ( .A(n142), .Y(n6562) );
  NAND2BXL U5124 ( .AN(n107), .B(n6986), .Y(n142) );
  BUFX3 U5125 ( .A(n145), .Y(n6561) );
  NAND2BXL U5126 ( .AN(n109), .B(n6986), .Y(n145) );
  BUFX3 U5127 ( .A(n147), .Y(n6560) );
  NAND2BXL U5128 ( .AN(n110), .B(n6986), .Y(n147) );
  BUFX3 U5129 ( .A(n149), .Y(n6559) );
  NAND2BXL U5130 ( .AN(n112), .B(n6986), .Y(n149) );
  BUFX3 U5131 ( .A(n151), .Y(n6558) );
  NAND2BXL U5132 ( .AN(n114), .B(n6986), .Y(n151) );
  BUFX3 U5133 ( .A(n153), .Y(n6557) );
  NAND2BXL U5134 ( .AN(n116), .B(n6986), .Y(n153) );
  BUFX3 U5135 ( .A(n155), .Y(n6556) );
  NAND2BXL U5136 ( .AN(n118), .B(n6986), .Y(n155) );
  BUFX3 U5137 ( .A(n157), .Y(n6555) );
  NAND2BXL U5138 ( .AN(n120), .B(n6986), .Y(n157) );
  BUFX3 U5139 ( .A(n159), .Y(n6554) );
  NAND2BXL U5140 ( .AN(n122), .B(n6986), .Y(n159) );
  BUFX3 U5141 ( .A(n161), .Y(n6553) );
  NAND2BXL U5142 ( .AN(n124), .B(n6986), .Y(n161) );
  BUFX3 U5143 ( .A(n163), .Y(n6552) );
  NAND2BXL U5144 ( .AN(n126), .B(n6986), .Y(n163) );
  BUFX3 U5145 ( .A(n165), .Y(n6551) );
  NAND2BXL U5146 ( .AN(n128), .B(n6985), .Y(n165) );
  BUFX3 U5147 ( .A(n167), .Y(n6550) );
  NAND2BXL U5148 ( .AN(n130), .B(n6985), .Y(n167) );
  BUFX3 U5149 ( .A(n169), .Y(n6549) );
  NAND2BXL U5150 ( .AN(n132), .B(n6985), .Y(n169) );
  BUFX3 U5151 ( .A(n171), .Y(n6548) );
  NAND2BXL U5152 ( .AN(n498), .B(n6985), .Y(n171) );
  BUFX3 U5153 ( .A(n173), .Y(n6547) );
  NAND2BXL U5154 ( .AN(n134), .B(n6985), .Y(n173) );
  BUFX3 U5155 ( .A(n176), .Y(n6546) );
  NAND2BXL U5156 ( .AN(n136), .B(n6985), .Y(n176) );
  BUFX3 U5157 ( .A(n179), .Y(n6545) );
  NAND2BXL U5158 ( .AN(n138), .B(n6985), .Y(n179) );
  BUFX3 U5159 ( .A(n181), .Y(n6544) );
  NAND2BXL U5160 ( .AN(n141), .B(n6985), .Y(n181) );
  BUFX3 U5161 ( .A(n183), .Y(n6543) );
  NAND2BXL U5162 ( .AN(n143), .B(n6985), .Y(n183) );
  BUFX3 U5163 ( .A(n185), .Y(n6542) );
  NAND2BXL U5164 ( .AN(n144), .B(n6985), .Y(n185) );
  BUFX3 U5165 ( .A(n187), .Y(n6541) );
  NAND2BXL U5166 ( .AN(n146), .B(n6985), .Y(n187) );
  BUFX3 U5167 ( .A(n189), .Y(n6540) );
  NAND2BXL U5168 ( .AN(n148), .B(n6985), .Y(n189) );
  BUFX3 U5169 ( .A(n191), .Y(n6539) );
  NAND2BXL U5170 ( .AN(n150), .B(n6984), .Y(n191) );
  BUFX3 U5171 ( .A(n193), .Y(n6538) );
  NAND2BXL U5172 ( .AN(n152), .B(n6984), .Y(n193) );
  BUFX3 U5173 ( .A(n195), .Y(n6537) );
  NAND2BXL U5174 ( .AN(n154), .B(n6984), .Y(n195) );
  BUFX3 U5175 ( .A(n197), .Y(n6536) );
  NAND2BXL U5176 ( .AN(n156), .B(n6984), .Y(n197) );
  BUFX3 U5177 ( .A(n199), .Y(n6535) );
  NAND2BXL U5178 ( .AN(n158), .B(n6984), .Y(n199) );
  BUFX3 U5179 ( .A(n201), .Y(n6534) );
  NAND2BXL U5180 ( .AN(n160), .B(n6984), .Y(n201) );
  BUFX3 U5181 ( .A(n203), .Y(n6533) );
  NAND2BXL U5182 ( .AN(n162), .B(n6984), .Y(n203) );
  BUFX3 U5183 ( .A(n205), .Y(n6532) );
  NAND2BXL U5184 ( .AN(n164), .B(n6984), .Y(n205) );
  BUFX3 U5185 ( .A(n207), .Y(n6531) );
  NAND2BXL U5186 ( .AN(n166), .B(n6984), .Y(n207) );
  BUFX3 U5187 ( .A(n210), .Y(n6530) );
  NAND2BXL U5188 ( .AN(n168), .B(n6984), .Y(n210) );
  BUFX3 U5189 ( .A(n213), .Y(n6529) );
  NAND2BXL U5190 ( .AN(n170), .B(n6984), .Y(n213) );
  BUFX3 U5191 ( .A(n215), .Y(n6528) );
  NAND2BXL U5192 ( .AN(n172), .B(n6984), .Y(n215) );
  BUFX3 U5193 ( .A(n217), .Y(n6527) );
  NAND2BXL U5194 ( .AN(n175), .B(n6984), .Y(n217) );
  BUFX3 U5195 ( .A(n219), .Y(n6526) );
  NAND2BXL U5196 ( .AN(n177), .B(n6983), .Y(n219) );
  BUFX3 U5197 ( .A(n221), .Y(n6525) );
  NAND2BXL U5198 ( .AN(n178), .B(n6983), .Y(n221) );
  BUFX3 U5199 ( .A(n223), .Y(n6524) );
  NAND2BXL U5200 ( .AN(n180), .B(n6983), .Y(n223) );
  BUFX3 U5201 ( .A(n225), .Y(n6523) );
  NAND2BXL U5202 ( .AN(n182), .B(n6983), .Y(n225) );
  BUFX3 U5203 ( .A(n227), .Y(n6522) );
  NAND2BXL U5204 ( .AN(n184), .B(n6983), .Y(n227) );
  BUFX3 U5205 ( .A(n229), .Y(n6521) );
  NAND2BXL U5206 ( .AN(n186), .B(n6983), .Y(n229) );
  BUFX3 U5207 ( .A(n231), .Y(n6520) );
  NAND2BXL U5208 ( .AN(n188), .B(n6983), .Y(n231) );
  BUFX3 U5209 ( .A(n233), .Y(n6519) );
  NAND2BXL U5210 ( .AN(n190), .B(n6983), .Y(n233) );
  BUFX3 U5211 ( .A(n235), .Y(n6518) );
  NAND2BXL U5212 ( .AN(n192), .B(n6983), .Y(n235) );
  BUFX3 U5213 ( .A(n237), .Y(n6517) );
  NAND2BXL U5214 ( .AN(n194), .B(n6983), .Y(n237) );
  BUFX3 U5215 ( .A(n239), .Y(n6516) );
  NAND2BXL U5216 ( .AN(n196), .B(n6983), .Y(n239) );
  BUFX3 U5217 ( .A(n241), .Y(n6515) );
  NAND2BXL U5218 ( .AN(n198), .B(n6983), .Y(n241) );
  BUFX3 U5219 ( .A(n243), .Y(n6514) );
  NAND2BXL U5220 ( .AN(n200), .B(n6983), .Y(n243) );
  BUFX3 U5221 ( .A(n246), .Y(n6513) );
  NAND2BXL U5222 ( .AN(n202), .B(n6982), .Y(n246) );
  BUFX3 U5223 ( .A(n248), .Y(n6512) );
  NAND2BXL U5224 ( .AN(n204), .B(n6982), .Y(n248) );
  BUFX3 U5225 ( .A(n250), .Y(n6511) );
  NAND2BXL U5226 ( .AN(n206), .B(n6982), .Y(n250) );
  BUFX3 U5227 ( .A(n252), .Y(n6510) );
  NAND2BXL U5228 ( .AN(n209), .B(n6982), .Y(n252) );
  BUFX3 U5229 ( .A(n254), .Y(n6509) );
  NAND2BXL U5230 ( .AN(n211), .B(n6982), .Y(n254) );
  BUFX3 U5231 ( .A(n256), .Y(n6508) );
  NAND2BXL U5232 ( .AN(n212), .B(n6982), .Y(n256) );
  BUFX3 U5233 ( .A(n258), .Y(n6507) );
  NAND2BXL U5234 ( .AN(n214), .B(n6982), .Y(n258) );
  BUFX3 U5235 ( .A(n260), .Y(n6506) );
  NAND2BXL U5236 ( .AN(n216), .B(n6982), .Y(n260) );
  BUFX3 U5237 ( .A(n262), .Y(n6505) );
  NAND2BXL U5238 ( .AN(n218), .B(n6982), .Y(n262) );
  BUFX3 U5239 ( .A(n266), .Y(n6503) );
  NAND2BXL U5240 ( .AN(n220), .B(n6982), .Y(n266) );
  BUFX3 U5241 ( .A(n268), .Y(n6502) );
  NAND2BXL U5242 ( .AN(n222), .B(n6982), .Y(n268) );
  BUFX3 U5243 ( .A(n270), .Y(n6501) );
  NAND2BXL U5244 ( .AN(n224), .B(n6982), .Y(n270) );
  BUFX3 U5245 ( .A(n272), .Y(n6500) );
  NAND2BXL U5246 ( .AN(n226), .B(n6981), .Y(n272) );
  BUFX3 U5247 ( .A(n274), .Y(n6499) );
  NAND2BXL U5248 ( .AN(n228), .B(n6981), .Y(n274) );
  BUFX3 U5249 ( .A(n276), .Y(n6498) );
  NAND2BXL U5250 ( .AN(n230), .B(n6981), .Y(n276) );
  BUFX3 U5251 ( .A(n279), .Y(n6497) );
  NAND2BXL U5252 ( .AN(n232), .B(n6981), .Y(n279) );
  BUFX3 U5253 ( .A(n281), .Y(n6496) );
  NAND2BXL U5254 ( .AN(n234), .B(n6981), .Y(n281) );
  BUFX3 U5255 ( .A(n283), .Y(n6495) );
  NAND2BXL U5256 ( .AN(n236), .B(n6981), .Y(n283) );
  BUFX3 U5257 ( .A(n285), .Y(n6494) );
  NAND2BXL U5258 ( .AN(n238), .B(n6981), .Y(n285) );
  BUFX3 U5259 ( .A(n287), .Y(n6493) );
  NAND2BXL U5260 ( .AN(n240), .B(n6981), .Y(n287) );
  BUFX3 U5261 ( .A(n289), .Y(n6492) );
  NAND2BXL U5262 ( .AN(n242), .B(n6981), .Y(n289) );
  BUFX3 U5263 ( .A(n291), .Y(n6491) );
  NAND2BXL U5264 ( .AN(n244), .B(n6981), .Y(n291) );
  BUFX3 U5265 ( .A(n293), .Y(n6490) );
  NAND2BXL U5266 ( .AN(n245), .B(n6981), .Y(n293) );
  BUFX3 U5267 ( .A(n295), .Y(n6489) );
  NAND2BXL U5268 ( .AN(n247), .B(n6981), .Y(n295) );
  BUFX3 U5269 ( .A(n297), .Y(n6488) );
  NAND2BXL U5270 ( .AN(n249), .B(n6981), .Y(n297) );
  BUFX3 U5271 ( .A(n299), .Y(n6487) );
  NAND2BXL U5272 ( .AN(n251), .B(n6990), .Y(n299) );
  BUFX3 U5273 ( .A(n301), .Y(n6486) );
  NAND2BXL U5274 ( .AN(n253), .B(n6985), .Y(n301) );
  BUFX3 U5275 ( .A(n303), .Y(n6485) );
  NAND2BXL U5276 ( .AN(n255), .B(n6983), .Y(n303) );
  BUFX3 U5277 ( .A(n305), .Y(n6484) );
  NAND2BXL U5278 ( .AN(n257), .B(n6987), .Y(n305) );
  BUFX3 U5279 ( .A(n307), .Y(n6483) );
  NAND2BXL U5280 ( .AN(n259), .B(n6991), .Y(n307) );
  BUFX3 U5281 ( .A(n309), .Y(n6482) );
  NAND2BXL U5282 ( .AN(n261), .B(n6988), .Y(n309) );
  BUFX3 U5283 ( .A(n312), .Y(n6481) );
  NAND2BXL U5284 ( .AN(n263), .B(n6986), .Y(n312) );
  BUFX3 U5285 ( .A(n314), .Y(n6480) );
  NAND2BXL U5286 ( .AN(n265), .B(n7000), .Y(n314) );
  BUFX3 U5287 ( .A(n316), .Y(n6479) );
  NAND2BXL U5288 ( .AN(n267), .B(n6986), .Y(n316) );
  BUFX3 U5289 ( .A(n318), .Y(n6478) );
  NAND2BXL U5290 ( .AN(n269), .B(n6982), .Y(n318) );
  BUFX3 U5291 ( .A(n320), .Y(n6477) );
  NAND2BXL U5292 ( .AN(n500), .B(n6988), .Y(n320) );
  BUFX3 U5293 ( .A(n322), .Y(n6476) );
  NAND2BXL U5294 ( .AN(n502), .B(n6986), .Y(n322) );
  BUFX3 U5295 ( .A(n324), .Y(n6475) );
  NAND2BXL U5296 ( .AN(n504), .B(n6985), .Y(n324) );
  BUFX3 U5297 ( .A(n326), .Y(n6474) );
  NAND2BXL U5298 ( .AN(n271), .B(mem_write_en), .Y(n326) );
  BUFX3 U5299 ( .A(n328), .Y(n6473) );
  NAND2BXL U5300 ( .AN(n273), .B(n6991), .Y(n328) );
  BUFX3 U5301 ( .A(n330), .Y(n6472) );
  NAND2BXL U5302 ( .AN(n275), .B(n6991), .Y(n330) );
  BUFX3 U5303 ( .A(n332), .Y(n6471) );
  NAND2BXL U5304 ( .AN(n277), .B(n6991), .Y(n332) );
  BUFX3 U5305 ( .A(n334), .Y(n6470) );
  NAND2BXL U5306 ( .AN(n278), .B(n6991), .Y(n334) );
  BUFX3 U5307 ( .A(n336), .Y(n6469) );
  NAND2BXL U5308 ( .AN(n280), .B(n6991), .Y(n336) );
  BUFX3 U5309 ( .A(n338), .Y(n6468) );
  NAND2BXL U5310 ( .AN(n282), .B(n6991), .Y(n338) );
  BUFX3 U5311 ( .A(n340), .Y(n6467) );
  NAND2BXL U5312 ( .AN(n284), .B(n6991), .Y(n340) );
  BUFX3 U5313 ( .A(n343), .Y(n6466) );
  NAND2BXL U5314 ( .AN(n286), .B(n6991), .Y(n343) );
  BUFX3 U5315 ( .A(n346), .Y(n6465) );
  NAND2BXL U5316 ( .AN(n288), .B(n6991), .Y(n346) );
  BUFX3 U5317 ( .A(n348), .Y(n6464) );
  NAND2BXL U5318 ( .AN(n290), .B(mem_write_en), .Y(n348) );
  BUFX3 U5319 ( .A(n350), .Y(n6463) );
  NAND2BXL U5320 ( .AN(n292), .B(mem_write_en), .Y(n350) );
  BUFX3 U5321 ( .A(n352), .Y(n6462) );
  NAND2BXL U5322 ( .AN(n294), .B(n6979), .Y(n352) );
  BUFX3 U5323 ( .A(n354), .Y(n6461) );
  NAND2BXL U5324 ( .AN(n506), .B(n6979), .Y(n354) );
  BUFX3 U5325 ( .A(n356), .Y(n6460) );
  NAND2BXL U5326 ( .AN(n508), .B(n6979), .Y(n356) );
  BUFX3 U5327 ( .A(n358), .Y(n6459) );
  NAND2BXL U5328 ( .AN(n510), .B(n6979), .Y(n358) );
  BUFX3 U5329 ( .A(n360), .Y(n6458) );
  NAND2BXL U5330 ( .AN(n296), .B(n6979), .Y(n360) );
  BUFX3 U5331 ( .A(n362), .Y(n6457) );
  NAND2BXL U5332 ( .AN(n298), .B(n6979), .Y(n362) );
  BUFX3 U5333 ( .A(n364), .Y(n6456) );
  NAND2BXL U5334 ( .AN(n300), .B(n7000), .Y(n364) );
  BUFX3 U5335 ( .A(n366), .Y(n6455) );
  NAND2BXL U5336 ( .AN(n302), .B(n7000), .Y(n366) );
  BUFX3 U5337 ( .A(n368), .Y(n6454) );
  NAND2BXL U5338 ( .AN(n304), .B(n7000), .Y(n368) );
  BUFX3 U5339 ( .A(n370), .Y(n6453) );
  NAND2BXL U5340 ( .AN(n306), .B(n7000), .Y(n370) );
  BUFX3 U5341 ( .A(n372), .Y(n6452) );
  NAND2BXL U5342 ( .AN(n308), .B(n6990), .Y(n372) );
  BUFX3 U5343 ( .A(n374), .Y(n6451) );
  NAND2BXL U5344 ( .AN(n310), .B(n6987), .Y(n374) );
  BUFX3 U5345 ( .A(n376), .Y(n6450) );
  NAND2BXL U5346 ( .AN(n311), .B(n6985), .Y(n376) );
  BUFX3 U5347 ( .A(n379), .Y(n6449) );
  NAND2BXL U5348 ( .AN(n313), .B(n6988), .Y(n379) );
  BUFX3 U5349 ( .A(n381), .Y(n6448) );
  NAND2BXL U5350 ( .AN(n315), .B(n6986), .Y(n381) );
  BUFX3 U5351 ( .A(n383), .Y(n6447) );
  NAND2BXL U5352 ( .AN(n317), .B(n6989), .Y(n383) );
  BUFX3 U5353 ( .A(n385), .Y(n6446) );
  NAND2BXL U5354 ( .AN(n319), .B(n6990), .Y(n385) );
  BUFX3 U5355 ( .A(n387), .Y(n6445) );
  NAND2BXL U5356 ( .AN(n549), .B(n6987), .Y(n387) );
  BUFX3 U5357 ( .A(n389), .Y(n6444) );
  NAND2BXL U5358 ( .AN(n552), .B(n6985), .Y(n389) );
  BUFX3 U5359 ( .A(n391), .Y(n6443) );
  NAND2BXL U5360 ( .AN(n555), .B(n6988), .Y(n391) );
  BUFX3 U5361 ( .A(n393), .Y(n6442) );
  NAND2BXL U5362 ( .AN(n321), .B(n6986), .Y(n393) );
  BUFX3 U5363 ( .A(n395), .Y(n6441) );
  NAND2BXL U5364 ( .AN(n323), .B(n6989), .Y(n395) );
  BUFX3 U5365 ( .A(n399), .Y(n6439) );
  NAND2BXL U5366 ( .AN(n325), .B(n6987), .Y(n399) );
  BUFX3 U5367 ( .A(n401), .Y(n6438) );
  NAND2BXL U5368 ( .AN(n327), .B(n6986), .Y(n401) );
  BUFX3 U5369 ( .A(n403), .Y(n6437) );
  NAND2BXL U5370 ( .AN(n329), .B(n6989), .Y(n403) );
  BUFX3 U5371 ( .A(n405), .Y(n6436) );
  NAND2BXL U5372 ( .AN(n331), .B(n6990), .Y(n405) );
  BUFX3 U5373 ( .A(n407), .Y(n6435) );
  NAND2BXL U5374 ( .AN(n333), .B(n6985), .Y(n407) );
  BUFX3 U5375 ( .A(n409), .Y(n6434) );
  NAND2BXL U5376 ( .AN(n335), .B(n6988), .Y(n409) );
  BUFX3 U5377 ( .A(n412), .Y(n6433) );
  NAND2BXL U5378 ( .AN(n337), .B(n6987), .Y(n412) );
  BUFX3 U5379 ( .A(n414), .Y(n6432) );
  NAND2BXL U5380 ( .AN(n339), .B(n6986), .Y(n414) );
  BUFX3 U5381 ( .A(n416), .Y(n6431) );
  NAND2BXL U5382 ( .AN(n342), .B(n6989), .Y(n416) );
  BUFX3 U5383 ( .A(n418), .Y(n6430) );
  NAND2BXL U5384 ( .AN(n344), .B(n6990), .Y(n418) );
  BUFX3 U5385 ( .A(n420), .Y(n6429) );
  NAND2BXL U5386 ( .AN(n511), .B(n6985), .Y(n420) );
  BUFX3 U5387 ( .A(n422), .Y(n6428) );
  NAND2BXL U5388 ( .AN(n513), .B(n6988), .Y(n422) );
  BUFX3 U5389 ( .A(n424), .Y(n6427) );
  NAND2BXL U5390 ( .AN(n515), .B(n6987), .Y(n424) );
  BUFX3 U5391 ( .A(n426), .Y(n6426) );
  NAND2BXL U5392 ( .AN(n345), .B(n6981), .Y(n426) );
  BUFX3 U5393 ( .A(n428), .Y(n6425) );
  NAND2BXL U5394 ( .AN(n347), .B(n6984), .Y(n428) );
  BUFX3 U5395 ( .A(n430), .Y(n6424) );
  NAND2BXL U5396 ( .AN(n349), .B(n6983), .Y(n430) );
  BUFX3 U5397 ( .A(n432), .Y(n6423) );
  NAND2BXL U5398 ( .AN(n351), .B(n6982), .Y(n432) );
  BUFX3 U5399 ( .A(n434), .Y(n6422) );
  NAND2BXL U5400 ( .AN(n353), .B(n6981), .Y(n434) );
  BUFX3 U5401 ( .A(n436), .Y(n6421) );
  NAND2BXL U5402 ( .AN(n355), .B(n6984), .Y(n436) );
  BUFX3 U5403 ( .A(n438), .Y(n6420) );
  NAND2BXL U5404 ( .AN(n357), .B(n6983), .Y(n438) );
  BUFX3 U5405 ( .A(n440), .Y(n6419) );
  NAND2BXL U5406 ( .AN(n359), .B(n6982), .Y(n440) );
  BUFX3 U5407 ( .A(n442), .Y(n6418) );
  NAND2BXL U5408 ( .AN(n361), .B(n6981), .Y(n442) );
  BUFX3 U5409 ( .A(n445), .Y(n6417) );
  NAND2BXL U5410 ( .AN(n363), .B(n6984), .Y(n445) );
  BUFX3 U5411 ( .A(n447), .Y(n6416) );
  NAND2BXL U5412 ( .AN(n365), .B(n6983), .Y(n447) );
  BUFX3 U5413 ( .A(n449), .Y(n6415) );
  NAND2BXL U5414 ( .AN(n367), .B(n6982), .Y(n449) );
  BUFX3 U5415 ( .A(n451), .Y(n6414) );
  NAND2BXL U5416 ( .AN(n369), .B(n6999), .Y(n451) );
  BUFX3 U5417 ( .A(n453), .Y(n6413) );
  NAND2BXL U5418 ( .AN(n371), .B(n6992), .Y(n453) );
  BUFX3 U5419 ( .A(n455), .Y(n6412) );
  NAND2BXL U5420 ( .AN(n373), .B(n6992), .Y(n455) );
  BUFX3 U5421 ( .A(n457), .Y(n6411) );
  NAND2BXL U5422 ( .AN(n375), .B(n6999), .Y(n457) );
  BUFX3 U5423 ( .A(n459), .Y(n6410) );
  NAND2BXL U5424 ( .AN(n377), .B(n6992), .Y(n459) );
  BUFX3 U5425 ( .A(n461), .Y(n6409) );
  NAND2BXL U5426 ( .AN(n378), .B(n6992), .Y(n461) );
  BUFX3 U5427 ( .A(n463), .Y(n6408) );
  NAND2BXL U5428 ( .AN(n380), .B(n6999), .Y(n463) );
  BUFX3 U5429 ( .A(n465), .Y(n6407) );
  NAND2BXL U5430 ( .AN(n382), .B(n6992), .Y(n465) );
  BUFX3 U5431 ( .A(n467), .Y(n6406) );
  NAND2BXL U5432 ( .AN(n384), .B(n6999), .Y(n467) );
  BUFX3 U5433 ( .A(n469), .Y(n6405) );
  NAND2BXL U5434 ( .AN(n386), .B(n6992), .Y(n469) );
  BUFX3 U5435 ( .A(n471), .Y(n6404) );
  NAND2BXL U5436 ( .AN(n388), .B(n6992), .Y(n471) );
  BUFX3 U5437 ( .A(n473), .Y(n6403) );
  NAND2BXL U5438 ( .AN(n390), .B(n6999), .Y(n473) );
  BUFX3 U5439 ( .A(n476), .Y(n6402) );
  NAND2BXL U5440 ( .AN(n392), .B(n6985), .Y(n476) );
  BUFX3 U5441 ( .A(n479), .Y(n6401) );
  NAND2BXL U5442 ( .AN(n394), .B(n6981), .Y(n479) );
  BUFX3 U5443 ( .A(n481), .Y(n6400) );
  NAND2BXL U5444 ( .AN(n396), .B(n6984), .Y(n481) );
  BUFX3 U5445 ( .A(n483), .Y(n6399) );
  NAND2BXL U5446 ( .AN(n398), .B(n6998), .Y(n483) );
  BUFX3 U5447 ( .A(n485), .Y(n6398) );
  NAND2BXL U5448 ( .AN(n400), .B(n6984), .Y(n485) );
  BUFX3 U5449 ( .A(n487), .Y(n6397) );
  NAND2BXL U5450 ( .AN(n402), .B(n6983), .Y(n487) );
  BUFX3 U5451 ( .A(n489), .Y(n6396) );
  NAND2BXL U5452 ( .AN(n404), .B(n6998), .Y(n489) );
  BUFX3 U5453 ( .A(n491), .Y(n6395) );
  NAND2BXL U5454 ( .AN(n406), .B(n6983), .Y(n491) );
  BUFX3 U5455 ( .A(n493), .Y(n6394) );
  NAND2BXL U5456 ( .AN(n408), .B(n6982), .Y(n493) );
  BUFX3 U5457 ( .A(n495), .Y(n6393) );
  NAND2BXL U5458 ( .AN(n410), .B(n6998), .Y(n495) );
  BUFX3 U5459 ( .A(n497), .Y(n6392) );
  NAND2BXL U5460 ( .AN(n411), .B(n6982), .Y(n497) );
  BUFX3 U5461 ( .A(n499), .Y(n6391) );
  NAND2BXL U5462 ( .AN(n413), .B(n6981), .Y(n499) );
  BUFX3 U5463 ( .A(n501), .Y(n6390) );
  NAND2BXL U5464 ( .AN(n415), .B(n6985), .Y(n501) );
  BUFX3 U5465 ( .A(n503), .Y(n6389) );
  NAND2BXL U5466 ( .AN(n417), .B(n6981), .Y(n503) );
  BUFX3 U5467 ( .A(n505), .Y(n6388) );
  NAND2BXL U5468 ( .AN(n22), .B(mem_write_en), .Y(n505) );
  BUFX3 U5469 ( .A(n507), .Y(n6387) );
  NAND2BXL U5470 ( .AN(n23), .B(n6987), .Y(n507) );
  BUFX3 U5471 ( .A(n509), .Y(n6386) );
  NAND2BXL U5472 ( .AN(n24), .B(n6992), .Y(n509) );
  BUFX3 U5473 ( .A(n512), .Y(n6385) );
  NAND2BXL U5474 ( .AN(n25), .B(n6998), .Y(n512) );
  BUFX3 U5475 ( .A(n514), .Y(n6384) );
  NAND2BXL U5476 ( .AN(n26), .B(mem_write_en), .Y(n514) );
  BUFX3 U5477 ( .A(n516), .Y(n6383) );
  NAND2BXL U5478 ( .AN(n28), .B(n6988), .Y(n516) );
  BUFX3 U5479 ( .A(n518), .Y(n6382) );
  NAND2BXL U5480 ( .AN(n29), .B(n6984), .Y(n518) );
  BUFX3 U5481 ( .A(n520), .Y(n6381) );
  NAND2BXL U5482 ( .AN(n31), .B(mem_write_en), .Y(n520) );
  BUFX3 U5483 ( .A(n522), .Y(n6380) );
  NAND2BXL U5484 ( .AN(n32), .B(n6989), .Y(n522) );
  BUFX3 U5485 ( .A(n524), .Y(n6379) );
  NAND2BXL U5486 ( .AN(n34), .B(n6992), .Y(n524) );
  BUFX3 U5487 ( .A(n526), .Y(n6378) );
  NAND2BXL U5488 ( .AN(n35), .B(n6987), .Y(n526) );
  BUFX3 U5489 ( .A(n528), .Y(n6377) );
  NAND2BXL U5490 ( .AN(n37), .B(n6998), .Y(n528) );
  BUFX3 U5491 ( .A(n532), .Y(n6375) );
  NAND2BXL U5492 ( .AN(n419), .B(n6985), .Y(n532) );
  BUFX3 U5493 ( .A(n534), .Y(n6374) );
  NAND2BXL U5494 ( .AN(n421), .B(n6986), .Y(n534) );
  BUFX3 U5495 ( .A(n536), .Y(n6373) );
  NAND2BXL U5496 ( .AN(n423), .B(n6981), .Y(n536) );
  BUFX3 U5497 ( .A(n538), .Y(n6372) );
  NAND2BXL U5498 ( .AN(n425), .B(n6989), .Y(n538) );
  BUFX3 U5499 ( .A(n540), .Y(n6371) );
  NAND2BXL U5500 ( .AN(n427), .B(n6988), .Y(n540) );
  BUFX3 U5501 ( .A(n542), .Y(n6370) );
  NAND2BXL U5502 ( .AN(n429), .B(n6989), .Y(n542) );
  BUFX3 U5503 ( .A(n547), .Y(n6369) );
  NAND2BXL U5504 ( .AN(n431), .B(n6990), .Y(n547) );
  BUFX3 U5505 ( .A(n550), .Y(n6368) );
  NAND2BXL U5506 ( .AN(n433), .B(n6984), .Y(n550) );
  BUFX3 U5507 ( .A(n553), .Y(n6367) );
  NAND2BXL U5508 ( .AN(n435), .B(n6983), .Y(n553) );
  BUFX3 U5509 ( .A(n556), .Y(n6366) );
  NAND2BXL U5510 ( .AN(n437), .B(n6982), .Y(n556) );
  BUFX3 U5511 ( .A(n559), .Y(n6365) );
  NAND2BXL U5512 ( .AN(n439), .B(n6981), .Y(n559) );
  BUFX3 U5513 ( .A(n561), .Y(n6364) );
  NAND2BXL U5514 ( .AN(n441), .B(n6984), .Y(n561) );
  BUFX3 U5515 ( .A(n563), .Y(n6363) );
  NAND2BXL U5516 ( .AN(n443), .B(n6983), .Y(n563) );
  BUFX3 U5517 ( .A(n565), .Y(n6362) );
  NAND2BXL U5518 ( .AN(n444), .B(n6982), .Y(n565) );
  BUFX3 U5519 ( .A(n568), .Y(n6361) );
  NAND2BXL U5520 ( .AN(n446), .B(n6990), .Y(n568) );
  BUFX3 U5521 ( .A(n570), .Y(n6360) );
  NAND2BXL U5522 ( .AN(n448), .B(n6990), .Y(n570) );
  BUFX3 U5523 ( .A(n572), .Y(n6359) );
  NAND2BXL U5524 ( .AN(n450), .B(n6990), .Y(n572) );
  BUFX3 U5525 ( .A(n574), .Y(n6358) );
  NAND2BXL U5526 ( .AN(n452), .B(n6990), .Y(n574) );
  BUFX3 U5527 ( .A(n577), .Y(n6357) );
  NAND2BXL U5528 ( .AN(n454), .B(n6990), .Y(n577) );
  BUFX3 U5529 ( .A(n579), .Y(n6356) );
  NAND2BXL U5530 ( .AN(n456), .B(n6990), .Y(n579) );
  BUFX3 U5531 ( .A(n581), .Y(n6355) );
  NAND2BXL U5532 ( .AN(n458), .B(n6990), .Y(n581) );
  INVX1 U5533 ( .A(n7011), .Y(n7010) );
  INVX1 U5534 ( .A(n7014), .Y(n7015) );
  INVX1 U5535 ( .A(n6049), .Y(n6024) );
  INVX1 U5536 ( .A(n6074), .Y(n6076) );
  INVX1 U5537 ( .A(n7006), .Y(n6074) );
  BUFX3 U5538 ( .A(n129), .Y(n6568) );
  NAND2BXL U5539 ( .AN(n460), .B(n6987), .Y(n129) );
  BUFX3 U5540 ( .A(n264), .Y(n6504) );
  NAND2BXL U5541 ( .AN(n462), .B(n6982), .Y(n264) );
  BUFX3 U5542 ( .A(n397), .Y(n6440) );
  NAND2BXL U5543 ( .AN(n464), .B(n6990), .Y(n397) );
  BUFX3 U5544 ( .A(n530), .Y(n6376) );
  NAND2BXL U5545 ( .AN(n38), .B(n6989), .Y(n530) );
  INVX1 U5546 ( .A(n7001), .Y(n6998) );
  INVX1 U5547 ( .A(n6993), .Y(n6999) );
  INVX1 U5548 ( .A(n6864), .Y(n6883) );
  INVX1 U5549 ( .A(n6841), .Y(n6860) );
  INVX1 U5550 ( .A(n6818), .Y(n6837) );
  INVX1 U5551 ( .A(n6795), .Y(n6814) );
  INVX1 U5552 ( .A(n6772), .Y(n6791) );
  INVX1 U5553 ( .A(n6749), .Y(n6768) );
  INVX1 U5554 ( .A(n6726), .Y(n6745) );
  INVX1 U5555 ( .A(n6703), .Y(n6722) );
  INVX1 U5556 ( .A(n6680), .Y(n6699) );
  INVX1 U5557 ( .A(n6657), .Y(n6676) );
  INVX1 U5558 ( .A(n6634), .Y(n6653) );
  INVX1 U5559 ( .A(n6611), .Y(n6630) );
  INVX1 U5560 ( .A(n6956), .Y(n6975) );
  INVX1 U5561 ( .A(n6933), .Y(n6952) );
  INVX1 U5562 ( .A(n6910), .Y(n6929) );
  INVX1 U5563 ( .A(n6887), .Y(n6906) );
  INVX1 U5564 ( .A(n6864), .Y(n6884) );
  INVX1 U5565 ( .A(n6841), .Y(n6861) );
  INVX1 U5566 ( .A(n6818), .Y(n6838) );
  INVX1 U5567 ( .A(n6795), .Y(n6815) );
  INVX1 U5568 ( .A(n6772), .Y(n6792) );
  INVX1 U5569 ( .A(n6749), .Y(n6769) );
  INVX1 U5570 ( .A(n6726), .Y(n6746) );
  INVX1 U5571 ( .A(n6703), .Y(n6723) );
  INVX1 U5572 ( .A(n6680), .Y(n6700) );
  INVX1 U5573 ( .A(n6657), .Y(n6677) );
  INVX1 U5574 ( .A(n6634), .Y(n6654) );
  INVX1 U5575 ( .A(n6611), .Y(n6631) );
  INVX1 U5576 ( .A(n6956), .Y(n6976) );
  INVX1 U5577 ( .A(n6933), .Y(n6953) );
  INVX1 U5578 ( .A(n6910), .Y(n6930) );
  INVX1 U5579 ( .A(n6887), .Y(n6907) );
  INVX1 U5580 ( .A(n6957), .Y(n6977) );
  INVX1 U5581 ( .A(n6934), .Y(n6954) );
  INVX1 U5582 ( .A(n6911), .Y(n6931) );
  INVX1 U5583 ( .A(n6888), .Y(n6908) );
  INVX1 U5584 ( .A(n6864), .Y(n6885) );
  INVX1 U5585 ( .A(n6841), .Y(n6862) );
  INVX1 U5586 ( .A(n6818), .Y(n6839) );
  INVX1 U5587 ( .A(n6795), .Y(n6816) );
  INVX1 U5588 ( .A(n6772), .Y(n6793) );
  INVX1 U5589 ( .A(n6749), .Y(n6770) );
  INVX1 U5590 ( .A(n6726), .Y(n6747) );
  INVX1 U5591 ( .A(n6703), .Y(n6724) );
  INVX1 U5592 ( .A(n6680), .Y(n6701) );
  INVX1 U5593 ( .A(n6657), .Y(n6678) );
  INVX1 U5594 ( .A(n6634), .Y(n6655) );
  INVX1 U5595 ( .A(n6611), .Y(n6632) );
  INVX1 U5596 ( .A(n6957), .Y(n6978) );
  INVX1 U5597 ( .A(n6934), .Y(n6955) );
  INVX1 U5598 ( .A(n6911), .Y(n6932) );
  INVX1 U5599 ( .A(n6888), .Y(n6909) );
  INVX1 U5600 ( .A(n6864), .Y(n6886) );
  INVX1 U5601 ( .A(n6841), .Y(n6863) );
  INVX1 U5602 ( .A(n6818), .Y(n6840) );
  INVX1 U5603 ( .A(n6795), .Y(n6817) );
  INVX1 U5604 ( .A(n6772), .Y(n6794) );
  INVX1 U5605 ( .A(n6749), .Y(n6771) );
  INVX1 U5606 ( .A(n6726), .Y(n6748) );
  INVX1 U5607 ( .A(n6703), .Y(n6725) );
  INVX1 U5608 ( .A(n6680), .Y(n6702) );
  INVX1 U5609 ( .A(n6657), .Y(n6679) );
  INVX1 U5610 ( .A(n6634), .Y(n6656) );
  INVX1 U5611 ( .A(n6611), .Y(n6633) );
  INVX1 U5612 ( .A(n7001), .Y(n7000) );
  INVX1 U5613 ( .A(n7002), .Y(n7005) );
  NOR2X1 U5614 ( .A(n7015), .B(n6017), .Y(n72) );
  NOR2X1 U5615 ( .A(n7004), .B(n7006), .Y(n545) );
  NOR2X1 U5616 ( .A(n7014), .B(N23), .Y(n106) );
  NOR2X1 U5617 ( .A(n7010), .B(n7012), .Y(n544) );
  NOR2X1 U5618 ( .A(n7005), .B(n7006), .Y(n548) );
  NOR2X1 U5619 ( .A(n7011), .B(n7012), .Y(n557) );
  AND2X2 U5620 ( .A(n7006), .B(n7004), .Y(n554) );
  AND2X2 U5621 ( .A(n6018), .B(n7015), .Y(n174) );
  AND2X2 U5622 ( .A(n7012), .B(n7010), .Y(n575) );
  INVX1 U5623 ( .A(n7008), .Y(n7011) );
  INVX1 U5624 ( .A(n6048), .Y(n6049) );
  INVX1 U5625 ( .A(n7012), .Y(n6048) );
  NOR2BX1 U5626 ( .AN(n6020), .B(n7015), .Y(n140) );
  NOR2BX1 U5627 ( .AN(n7006), .B(n7002), .Y(n551) );
  INVX1 U5628 ( .A(n6958), .Y(n6956) );
  INVX1 U5629 ( .A(n6935), .Y(n6933) );
  INVX1 U5630 ( .A(n6912), .Y(n6910) );
  INVX1 U5631 ( .A(n6889), .Y(n6887) );
  INVX1 U5632 ( .A(n1), .Y(n6864) );
  INVX1 U5633 ( .A(n2), .Y(n6841) );
  INVX1 U5634 ( .A(n3), .Y(n6818) );
  INVX1 U5635 ( .A(n4), .Y(n6795) );
  INVX1 U5636 ( .A(n5), .Y(n6772) );
  INVX1 U5637 ( .A(n6), .Y(n6749) );
  INVX1 U5638 ( .A(n12), .Y(n6726) );
  INVX1 U5639 ( .A(n13), .Y(n6703) );
  INVX1 U5640 ( .A(n14), .Y(n6680) );
  INVX1 U5641 ( .A(n15), .Y(n6657) );
  INVX1 U5642 ( .A(n16), .Y(n6634) );
  INVX1 U5643 ( .A(n17), .Y(n6611) );
  INVX1 U5644 ( .A(n6958), .Y(n6957) );
  INVX1 U5645 ( .A(n6935), .Y(n6934) );
  INVX1 U5646 ( .A(n6912), .Y(n6911) );
  INVX1 U5647 ( .A(n6889), .Y(n6888) );
  INVX1 U5648 ( .A(n6979), .Y(n7001) );
  NOR2BX1 U5649 ( .AN(n7012), .B(n7008), .Y(n566) );
  MX4X1 U5650 ( .A(n4986), .B(n4976), .C(n4981), .D(n4971), .S0(n6017), .S1(
        n6021), .Y(n4987) );
  MX4X1 U5651 ( .A(n4975), .B(n4973), .C(n4974), .D(n4972), .S0(n6043), .S1(
        n6059), .Y(n4976) );
  MX4X1 U5652 ( .A(n4985), .B(n4983), .C(n4984), .D(n4982), .S0(n6047), .S1(
        n6059), .Y(n4986) );
  MX4X1 U5653 ( .A(n4970), .B(n4968), .C(n4969), .D(n4967), .S0(n6042), .S1(
        n6059), .Y(n4971) );
  MX4X1 U5654 ( .A(n4776), .B(n4766), .C(n4771), .D(n4761), .S0(n6017), .S1(
        n6021), .Y(n4777) );
  MX4X1 U5655 ( .A(n4775), .B(n4773), .C(n4774), .D(n4772), .S0(n6033), .S1(
        n6056), .Y(n4776) );
  MX4X1 U5656 ( .A(n4765), .B(n4763), .C(n4764), .D(n4762), .S0(n6033), .S1(
        n6056), .Y(n4766) );
  MX4X1 U5657 ( .A(n4770), .B(n4768), .C(n4769), .D(n4767), .S0(n6033), .S1(
        n6056), .Y(n4771) );
  MX4X1 U5658 ( .A(n4860), .B(n4850), .C(n4855), .D(n4845), .S0(n6017), .S1(
        n6021), .Y(n4861) );
  MX4X1 U5659 ( .A(n4859), .B(n4857), .C(n4858), .D(n4856), .S0(n6038), .S1(
        n6057), .Y(n4860) );
  MX4X1 U5660 ( .A(n4849), .B(n4847), .C(n4848), .D(n4846), .S0(n6042), .S1(
        n6057), .Y(n4850) );
  MX4X1 U5661 ( .A(n4854), .B(n4852), .C(n4853), .D(n4851), .S0(n6045), .S1(
        n6057), .Y(n4855) );
  MX4X1 U5662 ( .A(n5028), .B(n5018), .C(n5023), .D(n5013), .S0(n6018), .S1(
        n6022), .Y(n5029) );
  MX4X1 U5663 ( .A(n5027), .B(n5025), .C(n5026), .D(n5024), .S0(n6034), .S1(
        n6060), .Y(n5028) );
  MX4X1 U5664 ( .A(n5017), .B(n5015), .C(n5016), .D(n5014), .S0(n6034), .S1(
        n6060), .Y(n5018) );
  MX4X1 U5665 ( .A(n5022), .B(n5020), .C(n5021), .D(n5019), .S0(n6034), .S1(
        n6060), .Y(n5023) );
  MX4X1 U5666 ( .A(n5112), .B(n5102), .C(n5107), .D(n5097), .S0(n6018), .S1(
        n6022), .Y(n5113) );
  MX4X1 U5667 ( .A(n5111), .B(n5109), .C(n5110), .D(n5108), .S0(n6035), .S1(
        n6061), .Y(n5112) );
  MX4X1 U5668 ( .A(n5101), .B(n5099), .C(n5100), .D(n5098), .S0(n6041), .S1(
        n6061), .Y(n5102) );
  MX4X1 U5669 ( .A(n5106), .B(n5104), .C(n5105), .D(n5103), .S0(n6036), .S1(
        n6061), .Y(n5107) );
  MX4X1 U5670 ( .A(n5196), .B(n5186), .C(n5191), .D(n5181), .S0(n6018), .S1(
        n6022), .Y(n5197) );
  MX4X1 U5671 ( .A(n5195), .B(n5193), .C(n5194), .D(n5192), .S0(n6035), .S1(
        n6062), .Y(n5196) );
  MX4X1 U5672 ( .A(n5185), .B(n5183), .C(n5184), .D(n5182), .S0(n6035), .S1(
        n6062), .Y(n5186) );
  MX4X1 U5673 ( .A(n5190), .B(n5188), .C(n5189), .D(n5187), .S0(n6035), .S1(
        n6062), .Y(n5191) );
  MX4X1 U5674 ( .A(n5280), .B(n5270), .C(n5275), .D(n5265), .S0(n6019), .S1(
        n6022), .Y(n5281) );
  MX4X1 U5675 ( .A(n5279), .B(n5277), .C(n5278), .D(n5276), .S0(n6036), .S1(
        n6064), .Y(n5280) );
  MX4X1 U5676 ( .A(n5269), .B(n5267), .C(n5268), .D(n5266), .S0(n6036), .S1(
        n6064), .Y(n5270) );
  MX4X1 U5677 ( .A(n5274), .B(n5272), .C(n5273), .D(n5271), .S0(n6036), .S1(
        n6064), .Y(n5275) );
  MX4X1 U5678 ( .A(n5364), .B(n5354), .C(n5359), .D(n5349), .S0(n6019), .S1(
        n6022), .Y(n5365) );
  MX4X1 U5679 ( .A(n5363), .B(n5361), .C(n5362), .D(n5360), .S0(n6037), .S1(
        n6065), .Y(n5364) );
  MX4X1 U5680 ( .A(n5353), .B(n5351), .C(n5352), .D(n5350), .S0(n6037), .S1(
        n6065), .Y(n5354) );
  MX4X1 U5681 ( .A(n5358), .B(n5356), .C(n5357), .D(n5355), .S0(n6037), .S1(
        n6065), .Y(n5359) );
  MX4X1 U5682 ( .A(n5448), .B(n5438), .C(n5443), .D(n5433), .S0(n6019), .S1(
        n6022), .Y(n5449) );
  MX4X1 U5683 ( .A(n5447), .B(n5445), .C(n5446), .D(n5444), .S0(n6038), .S1(
        n6066), .Y(n5448) );
  MX4X1 U5684 ( .A(n5437), .B(n5435), .C(n5436), .D(n5434), .S0(n6038), .S1(
        n6066), .Y(n5438) );
  MX4X1 U5685 ( .A(n5442), .B(n5440), .C(n5441), .D(n5439), .S0(n6038), .S1(
        n6066), .Y(n5443) );
  MX4X1 U5686 ( .A(n5532), .B(n5522), .C(n5527), .D(n5517), .S0(n6020), .S1(
        n6023), .Y(n5533) );
  MX4X1 U5687 ( .A(n5531), .B(n5529), .C(n5530), .D(n5528), .S0(n6040), .S1(
        n6068), .Y(n5532) );
  MX4X1 U5688 ( .A(n5521), .B(n5519), .C(n5520), .D(n5518), .S0(n6040), .S1(
        n6068), .Y(n5522) );
  MX4X1 U5689 ( .A(n5526), .B(n5524), .C(n5525), .D(n5523), .S0(n6040), .S1(
        n6068), .Y(n5527) );
  MX4X1 U5690 ( .A(n5616), .B(n5606), .C(n5611), .D(n5601), .S0(n6020), .S1(
        n6023), .Y(n5617) );
  MX4X1 U5691 ( .A(n5615), .B(n5613), .C(n5614), .D(n5612), .S0(n6041), .S1(
        n6069), .Y(n5616) );
  MX4X1 U5692 ( .A(n5605), .B(n5603), .C(n5604), .D(n5602), .S0(n6041), .S1(
        n6069), .Y(n5606) );
  MX4X1 U5693 ( .A(n5610), .B(n5608), .C(n5609), .D(n5607), .S0(n6041), .S1(
        n6069), .Y(n5611) );
  MX4X1 U5694 ( .A(n5700), .B(n5690), .C(n5695), .D(n5685), .S0(n6020), .S1(
        n6023), .Y(n5701) );
  MX4X1 U5695 ( .A(n5699), .B(n5697), .C(n5698), .D(n5696), .S0(n6042), .S1(
        n6070), .Y(n5700) );
  MX4X1 U5696 ( .A(n5689), .B(n5687), .C(n5688), .D(n5686), .S0(n6042), .S1(
        n6070), .Y(n5690) );
  MX4X1 U5697 ( .A(n5694), .B(n5692), .C(n5693), .D(n5691), .S0(n6042), .S1(
        n6070), .Y(n5695) );
  MX4X1 U5698 ( .A(n5784), .B(n5774), .C(n5779), .D(n5769), .S0(n6017), .S1(
        n6021), .Y(n5785) );
  MX4X1 U5699 ( .A(n5783), .B(n5781), .C(n5782), .D(n5780), .S0(n6044), .S1(
        n6072), .Y(n5784) );
  MX4X1 U5700 ( .A(n5773), .B(n5771), .C(n5772), .D(n5770), .S0(n6044), .S1(
        n6072), .Y(n5774) );
  MX4X1 U5701 ( .A(n5778), .B(n5776), .C(n5777), .D(n5775), .S0(n6044), .S1(
        n6072), .Y(n5779) );
  MX4X1 U5702 ( .A(n5868), .B(n5858), .C(n5863), .D(n5853), .S0(n6018), .S1(
        n6023), .Y(n5869) );
  MX4X1 U5703 ( .A(n5867), .B(n5865), .C(n5866), .D(n5864), .S0(n6045), .S1(
        n6073), .Y(n5868) );
  MX4X1 U5704 ( .A(n5857), .B(n5855), .C(n5856), .D(n5854), .S0(n6045), .S1(
        n6073), .Y(n5858) );
  MX4X1 U5705 ( .A(n5862), .B(n5860), .C(n5861), .D(n5859), .S0(n6045), .S1(
        n6073), .Y(n5863) );
  MX4X1 U5706 ( .A(n5952), .B(n5942), .C(n5947), .D(n5937), .S0(n6020), .S1(
        n6021), .Y(n5953) );
  MX4X1 U5707 ( .A(n5951), .B(n5949), .C(n5950), .D(n5948), .S0(n6046), .S1(
        n6061), .Y(n5952) );
  MX4X1 U5708 ( .A(n5941), .B(n5939), .C(n5940), .D(n5938), .S0(n6046), .S1(
        n6060), .Y(n5942) );
  MX4X1 U5709 ( .A(n5946), .B(n5944), .C(n5945), .D(n5943), .S0(n6046), .S1(
        n6073), .Y(n5947) );
  MX4X1 U5710 ( .A(n4734), .B(n4724), .C(n4729), .D(n4719), .S0(n6020), .S1(
        N22), .Y(n4735) );
  MX4X1 U5711 ( .A(n4733), .B(n4731), .C(n4732), .D(n4730), .S0(n6034), .S1(
        n6071), .Y(n4734) );
  MX4X1 U5712 ( .A(n4723), .B(n4721), .C(n4722), .D(n4720), .S0(n6039), .S1(
        n6065), .Y(n4724) );
  MX4X1 U5713 ( .A(n4728), .B(n4726), .C(n4727), .D(n4725), .S0(n6045), .S1(
        n6056), .Y(n4729) );
  MX4X1 U5714 ( .A(n4756), .B(n4714), .C(n4735), .D(n4693), .S0(N25), .S1(N24), 
        .Y(mem_read_data[0]) );
  MX4X1 U5715 ( .A(n4692), .B(n4682), .C(n4687), .D(n580), .S0(n6017), .S1(N22), .Y(n4693) );
  MX4X1 U5716 ( .A(n4755), .B(n4745), .C(n4750), .D(n4740), .S0(n6019), .S1(
        n7015), .Y(n4756) );
  MX4X1 U5717 ( .A(n4713), .B(n4703), .C(n4708), .D(n4698), .S0(n6018), .S1(
        n7015), .Y(n4714) );
  MX4X1 U5718 ( .A(n4840), .B(n4798), .C(n4819), .D(n4777), .S0(N25), .S1(N24), 
        .Y(mem_read_data[1]) );
  MX4X1 U5719 ( .A(n4839), .B(n4829), .C(n4834), .D(n4824), .S0(n6017), .S1(
        n6021), .Y(n4840) );
  MX4X1 U5720 ( .A(n4797), .B(n4787), .C(n4792), .D(n4782), .S0(n6017), .S1(
        n6021), .Y(n4798) );
  MX4X1 U5721 ( .A(n4818), .B(n4808), .C(n4813), .D(n4803), .S0(n6017), .S1(
        n6021), .Y(n4819) );
  MX4X1 U5722 ( .A(n4924), .B(n4882), .C(n4903), .D(n4861), .S0(N25), .S1(N24), 
        .Y(mem_read_data[2]) );
  MX4X1 U5723 ( .A(n4923), .B(n4913), .C(n4918), .D(n4908), .S0(n6017), .S1(
        n6021), .Y(n4924) );
  MX4X1 U5724 ( .A(n4881), .B(n4871), .C(n4876), .D(n4866), .S0(n6017), .S1(
        n6021), .Y(n4882) );
  MX4X1 U5725 ( .A(n4902), .B(n4892), .C(n4897), .D(n4887), .S0(n6017), .S1(
        n6021), .Y(n4903) );
  MX4X1 U5726 ( .A(n5008), .B(n4966), .C(n4987), .D(n4945), .S0(N25), .S1(N24), 
        .Y(mem_read_data[3]) );
  MX4X1 U5727 ( .A(n4965), .B(n4955), .C(n4960), .D(n4950), .S0(n6017), .S1(
        n6021), .Y(n4966) );
  MX4X1 U5728 ( .A(n5007), .B(n4997), .C(n5002), .D(n4992), .S0(n6017), .S1(
        n6021), .Y(n5008) );
  MX4X1 U5729 ( .A(n4944), .B(n4934), .C(n4939), .D(n4929), .S0(n6017), .S1(
        n6021), .Y(n4945) );
  MX4X1 U5730 ( .A(n5092), .B(n5050), .C(n5071), .D(n5029), .S0(N25), .S1(N24), 
        .Y(mem_read_data[4]) );
  MX4X1 U5731 ( .A(n5091), .B(n5081), .C(n5086), .D(n5076), .S0(n6018), .S1(
        n6022), .Y(n5092) );
  MX4X1 U5732 ( .A(n5049), .B(n5039), .C(n5044), .D(n5034), .S0(n6018), .S1(
        n6022), .Y(n5050) );
  MX4X1 U5733 ( .A(n5070), .B(n5060), .C(n5065), .D(n5055), .S0(n6018), .S1(
        n6022), .Y(n5071) );
  MX4X1 U5734 ( .A(n5176), .B(n5134), .C(n5155), .D(n5113), .S0(N25), .S1(N24), 
        .Y(mem_read_data[5]) );
  MX4X1 U5735 ( .A(n5175), .B(n5165), .C(n5170), .D(n5160), .S0(n6018), .S1(
        n6022), .Y(n5176) );
  MX4X1 U5736 ( .A(n5133), .B(n5123), .C(n5128), .D(n5118), .S0(n6018), .S1(
        n6022), .Y(n5134) );
  MX4X1 U5737 ( .A(n5154), .B(n5144), .C(n5149), .D(n5139), .S0(n6018), .S1(
        n6022), .Y(n5155) );
  MX4X1 U5738 ( .A(n5260), .B(n5218), .C(n5239), .D(n5197), .S0(N25), .S1(N24), 
        .Y(mem_read_data[6]) );
  MX4X1 U5739 ( .A(n5259), .B(n5249), .C(n5254), .D(n5244), .S0(n6018), .S1(
        n6022), .Y(n5260) );
  MX4X1 U5740 ( .A(n5217), .B(n5207), .C(n5212), .D(n5202), .S0(n6018), .S1(
        n6022), .Y(n5218) );
  MX4X1 U5741 ( .A(n5238), .B(n5228), .C(n5233), .D(n5223), .S0(n6018), .S1(
        n6022), .Y(n5239) );
  MX4X1 U5742 ( .A(n5344), .B(n5302), .C(n5323), .D(n5281), .S0(N25), .S1(N24), 
        .Y(mem_read_data[7]) );
  MX4X1 U5743 ( .A(n5343), .B(n5333), .C(n5338), .D(n5328), .S0(n6019), .S1(
        n6023), .Y(n5344) );
  MX4X1 U5744 ( .A(n5301), .B(n5291), .C(n5296), .D(n5286), .S0(n6019), .S1(
        n6022), .Y(n5302) );
  MX4X1 U5745 ( .A(n5322), .B(n5312), .C(n5317), .D(n5307), .S0(n6019), .S1(
        n6022), .Y(n5323) );
  MX4X1 U5746 ( .A(n5428), .B(n5386), .C(n5407), .D(n5365), .S0(N25), .S1(N24), 
        .Y(mem_read_data[8]) );
  MX4X1 U5747 ( .A(n5427), .B(n5417), .C(n5422), .D(n5412), .S0(n6019), .S1(
        n6021), .Y(n5428) );
  MX4X1 U5748 ( .A(n5385), .B(n5375), .C(n5380), .D(n5370), .S0(n6019), .S1(
        N22), .Y(n5386) );
  MX4X1 U5749 ( .A(n5406), .B(n5396), .C(n5401), .D(n5391), .S0(n6019), .S1(
        n6022), .Y(n5407) );
  MX4X1 U5750 ( .A(n5512), .B(n5470), .C(n5491), .D(n5449), .S0(N25), .S1(N24), 
        .Y(mem_read_data[9]) );
  MX4X1 U5751 ( .A(n5511), .B(n5501), .C(n5506), .D(n5496), .S0(n6019), .S1(
        N22), .Y(n5512) );
  MX4X1 U5752 ( .A(n5469), .B(n5459), .C(n5464), .D(n5454), .S0(n6019), .S1(
        n6023), .Y(n5470) );
  MX4X1 U5753 ( .A(n5490), .B(n5480), .C(n5485), .D(n5475), .S0(n6019), .S1(
        n6022), .Y(n5491) );
  MX4X1 U5754 ( .A(n5596), .B(n5554), .C(n5575), .D(n5533), .S0(N25), .S1(N24), 
        .Y(mem_read_data[10]) );
  MX4X1 U5755 ( .A(n5595), .B(n5585), .C(n5590), .D(n5580), .S0(n6020), .S1(
        n6023), .Y(n5596) );
  MX4X1 U5756 ( .A(n5574), .B(n5564), .C(n5569), .D(n5559), .S0(n6020), .S1(
        n6023), .Y(n5575) );
  MX4X1 U5757 ( .A(n5553), .B(n5543), .C(n5548), .D(n5538), .S0(n6020), .S1(
        n6023), .Y(n5554) );
  MX4X1 U5758 ( .A(n5680), .B(n5638), .C(n5659), .D(n5617), .S0(N25), .S1(N24), 
        .Y(mem_read_data[11]) );
  MX4X1 U5759 ( .A(n5679), .B(n5669), .C(n5674), .D(n5664), .S0(n6020), .S1(
        n6023), .Y(n5680) );
  MX4X1 U5760 ( .A(n5637), .B(n5627), .C(n5632), .D(n5622), .S0(n6020), .S1(
        n6023), .Y(n5638) );
  MX4X1 U5761 ( .A(n5658), .B(n5648), .C(n5653), .D(n5643), .S0(n6020), .S1(
        n6023), .Y(n5659) );
  MX4X1 U5762 ( .A(n5764), .B(n5722), .C(n5743), .D(n5701), .S0(N25), .S1(N24), 
        .Y(mem_read_data[12]) );
  MX4X1 U5763 ( .A(n5763), .B(n5753), .C(n5758), .D(n5748), .S0(n6020), .S1(
        n6023), .Y(n5764) );
  MX4X1 U5764 ( .A(n5721), .B(n5711), .C(n5716), .D(n5706), .S0(n6020), .S1(
        n6023), .Y(n5722) );
  MX4X1 U5765 ( .A(n5742), .B(n5732), .C(n5737), .D(n5727), .S0(n6020), .S1(
        n6023), .Y(n5743) );
  MX4X1 U5766 ( .A(n5848), .B(n5806), .C(n5827), .D(n5785), .S0(N25), .S1(N24), 
        .Y(mem_read_data[13]) );
  MX4X1 U5767 ( .A(n5847), .B(n5837), .C(n5842), .D(n5832), .S0(n6020), .S1(
        n6021), .Y(n5848) );
  MX4X1 U5768 ( .A(n5805), .B(n5795), .C(n5800), .D(n5790), .S0(n6017), .S1(
        n7015), .Y(n5806) );
  MX4X1 U5769 ( .A(n5826), .B(n5816), .C(n5821), .D(n5811), .S0(n6017), .S1(
        n6023), .Y(n5827) );
  MX4X1 U5770 ( .A(n5932), .B(n5890), .C(n5911), .D(n5869), .S0(N25), .S1(N24), 
        .Y(mem_read_data[14]) );
  MX4X1 U5771 ( .A(n5931), .B(n5921), .C(n5926), .D(n5916), .S0(n6019), .S1(
        n6023), .Y(n5932) );
  MX4X1 U5772 ( .A(n5889), .B(n5879), .C(n5884), .D(n5874), .S0(n6018), .S1(
        n6021), .Y(n5890) );
  MX4X1 U5773 ( .A(n5910), .B(n5900), .C(n5905), .D(n5895), .S0(n6019), .S1(
        n6021), .Y(n5911) );
  MX4X1 U5774 ( .A(n6016), .B(n5974), .C(n5995), .D(n5953), .S0(N25), .S1(N24), 
        .Y(mem_read_data[15]) );
  MX4X1 U5775 ( .A(n6015), .B(n6005), .C(n6010), .D(n6000), .S0(n6018), .S1(
        n6021), .Y(n6016) );
  MX4X1 U5776 ( .A(n5973), .B(n5963), .C(n5968), .D(n5958), .S0(n6019), .S1(
        n6023), .Y(n5974) );
  MX4X1 U5777 ( .A(n5994), .B(n5984), .C(n5989), .D(n5979), .S0(n6020), .S1(
        n6023), .Y(n5995) );
  INVX1 U5778 ( .A(n7003), .Y(n7002) );
  INVX1 U5779 ( .A(N18), .Y(n7003) );
  INVX1 U5780 ( .A(n7007), .Y(n7006) );
  INVX1 U5781 ( .A(N19), .Y(n7007) );
  INVX1 U5782 ( .A(n7013), .Y(n7012) );
  INVX1 U5783 ( .A(N21), .Y(n7013) );
  INVX1 U5784 ( .A(n7009), .Y(n7008) );
  INVX1 U5785 ( .A(N20), .Y(n7009) );
  INVX1 U5786 ( .A(N22), .Y(n7014) );
  INVX1 U5787 ( .A(n7), .Y(n6958) );
  INVX1 U5788 ( .A(n9), .Y(n6935) );
  INVX1 U5789 ( .A(n10), .Y(n6912) );
  INVX1 U5790 ( .A(n11), .Y(n6889) );
  INVX1 U5791 ( .A(N23), .Y(n7016) );
  INVX1 U5792 ( .A(n6980), .Y(n6979) );
  INVX1 U5793 ( .A(mem_write_en), .Y(n6980) );
  MX4X1 U5794 ( .A(\ram[84][0] ), .B(\ram[85][0] ), .C(\ram[86][0] ), .D(
        \ram[87][0] ), .S0(n6271), .S1(n6137), .Y(n4727) );
  MX4X1 U5795 ( .A(\ram[100][0] ), .B(\ram[101][0] ), .C(\ram[102][0] ), .D(
        \ram[103][0] ), .S0(n6270), .S1(n6136), .Y(n4722) );
  MX4X1 U5796 ( .A(\ram[68][0] ), .B(\ram[69][0] ), .C(\ram[70][0] ), .D(
        \ram[71][0] ), .S0(n6271), .S1(n6137), .Y(n4732) );
  MX4X1 U5797 ( .A(\ram[212][1] ), .B(\ram[213][1] ), .C(\ram[214][1] ), .D(
        \ram[215][1] ), .S0(n6273), .S1(n6139), .Y(n4769) );
  MX4X1 U5798 ( .A(\ram[228][1] ), .B(\ram[229][1] ), .C(\ram[230][1] ), .D(
        \ram[231][1] ), .S0(n6273), .S1(n6139), .Y(n4764) );
  MX4X1 U5799 ( .A(\ram[196][1] ), .B(\ram[197][1] ), .C(\ram[198][1] ), .D(
        \ram[199][1] ), .S0(n6274), .S1(n6140), .Y(n4774) );
  MX4X1 U5800 ( .A(\ram[212][2] ), .B(\ram[213][2] ), .C(\ram[214][2] ), .D(
        \ram[215][2] ), .S0(n6279), .S1(n6145), .Y(n4853) );
  MX4X1 U5801 ( .A(\ram[228][2] ), .B(\ram[229][2] ), .C(\ram[230][2] ), .D(
        \ram[231][2] ), .S0(n6278), .S1(n6144), .Y(n4848) );
  MX4X1 U5802 ( .A(\ram[196][2] ), .B(\ram[197][2] ), .C(\ram[198][2] ), .D(
        \ram[199][2] ), .S0(n6279), .S1(n6145), .Y(n4858) );
  MX4X1 U5803 ( .A(\ram[116][3] ), .B(\ram[117][3] ), .C(\ram[118][3] ), .D(
        \ram[119][3] ), .S0(n6286), .S1(n6152), .Y(n4969) );
  MX4X1 U5804 ( .A(\ram[68][3] ), .B(\ram[69][3] ), .C(\ram[70][3] ), .D(
        \ram[71][3] ), .S0(n6287), .S1(n6153), .Y(n4984) );
  MX4X1 U5805 ( .A(\ram[100][3] ), .B(\ram[101][3] ), .C(\ram[102][3] ), .D(
        \ram[103][3] ), .S0(n6286), .S1(n6152), .Y(n4974) );
  MX4X1 U5806 ( .A(\ram[212][4] ), .B(\ram[213][4] ), .C(\ram[214][4] ), .D(
        \ram[215][4] ), .S0(n6289), .S1(n6155), .Y(n5021) );
  MX4X1 U5807 ( .A(\ram[228][4] ), .B(\ram[229][4] ), .C(\ram[230][4] ), .D(
        \ram[231][4] ), .S0(n6289), .S1(n6155), .Y(n5016) );
  MX4X1 U5808 ( .A(\ram[196][4] ), .B(\ram[197][4] ), .C(\ram[198][4] ), .D(
        \ram[199][4] ), .S0(n6290), .S1(n6156), .Y(n5026) );
  MX4X1 U5809 ( .A(\ram[212][5] ), .B(\ram[213][5] ), .C(\ram[214][5] ), .D(
        \ram[215][5] ), .S0(n6295), .S1(n6161), .Y(n5105) );
  MX4X1 U5810 ( .A(\ram[228][5] ), .B(\ram[229][5] ), .C(\ram[230][5] ), .D(
        \ram[231][5] ), .S0(n6294), .S1(n6160), .Y(n5100) );
  MX4X1 U5811 ( .A(\ram[196][5] ), .B(\ram[197][5] ), .C(\ram[198][5] ), .D(
        \ram[199][5] ), .S0(n6295), .S1(n6161), .Y(n5110) );
  MX4X1 U5812 ( .A(\ram[212][6] ), .B(\ram[213][6] ), .C(\ram[214][6] ), .D(
        \ram[215][6] ), .S0(n6300), .S1(n6166), .Y(n5189) );
  MX4X1 U5813 ( .A(\ram[228][6] ), .B(\ram[229][6] ), .C(\ram[230][6] ), .D(
        \ram[231][6] ), .S0(n6300), .S1(n6166), .Y(n5184) );
  MX4X1 U5814 ( .A(\ram[196][6] ), .B(\ram[197][6] ), .C(\ram[198][6] ), .D(
        \ram[199][6] ), .S0(n6300), .S1(n6166), .Y(n5194) );
  MX4X1 U5815 ( .A(\ram[212][7] ), .B(\ram[213][7] ), .C(\ram[214][7] ), .D(
        \ram[215][7] ), .S0(n6305), .S1(n6171), .Y(n5273) );
  MX4X1 U5816 ( .A(\ram[228][7] ), .B(\ram[229][7] ), .C(\ram[230][7] ), .D(
        \ram[231][7] ), .S0(n6305), .S1(n6171), .Y(n5268) );
  MX4X1 U5817 ( .A(\ram[196][7] ), .B(\ram[197][7] ), .C(\ram[198][7] ), .D(
        \ram[199][7] ), .S0(n6306), .S1(n6172), .Y(n5278) );
  MX4X1 U5818 ( .A(\ram[212][8] ), .B(\ram[213][8] ), .C(\ram[214][8] ), .D(
        \ram[215][8] ), .S0(n6311), .S1(n6177), .Y(n5357) );
  MX4X1 U5819 ( .A(\ram[228][8] ), .B(\ram[229][8] ), .C(\ram[230][8] ), .D(
        \ram[231][8] ), .S0(n6310), .S1(n6176), .Y(n5352) );
  MX4X1 U5820 ( .A(\ram[196][8] ), .B(\ram[197][8] ), .C(\ram[198][8] ), .D(
        \ram[199][8] ), .S0(n6311), .S1(n6177), .Y(n5362) );
  MX4X1 U5821 ( .A(\ram[212][9] ), .B(\ram[213][9] ), .C(\ram[214][9] ), .D(
        \ram[215][9] ), .S0(n6316), .S1(n6182), .Y(n5441) );
  MX4X1 U5822 ( .A(\ram[228][9] ), .B(\ram[229][9] ), .C(\ram[230][9] ), .D(
        \ram[231][9] ), .S0(n6316), .S1(n6182), .Y(n5436) );
  MX4X1 U5823 ( .A(\ram[196][9] ), .B(\ram[197][9] ), .C(\ram[198][9] ), .D(
        \ram[199][9] ), .S0(n6316), .S1(n6182), .Y(n5446) );
  MX4X1 U5824 ( .A(\ram[212][10] ), .B(\ram[213][10] ), .C(\ram[214][10] ), 
        .D(\ram[215][10] ), .S0(n6321), .S1(n6187), .Y(n5525) );
  MX4X1 U5825 ( .A(\ram[228][10] ), .B(\ram[229][10] ), .C(\ram[230][10] ), 
        .D(\ram[231][10] ), .S0(n6321), .S1(n6187), .Y(n5520) );
  MX4X1 U5826 ( .A(\ram[196][10] ), .B(\ram[197][10] ), .C(\ram[198][10] ), 
        .D(\ram[199][10] ), .S0(n6322), .S1(n6188), .Y(n5530) );
  MX4X1 U5827 ( .A(\ram[212][11] ), .B(\ram[213][11] ), .C(\ram[214][11] ), 
        .D(\ram[215][11] ), .S0(n6327), .S1(n6193), .Y(n5609) );
  MX4X1 U5828 ( .A(\ram[228][11] ), .B(\ram[229][11] ), .C(\ram[230][11] ), 
        .D(\ram[231][11] ), .S0(n6326), .S1(n6192), .Y(n5604) );
  MX4X1 U5829 ( .A(\ram[196][11] ), .B(\ram[197][11] ), .C(\ram[198][11] ), 
        .D(\ram[199][11] ), .S0(n6327), .S1(n6193), .Y(n5614) );
  MX4X1 U5830 ( .A(\ram[212][12] ), .B(\ram[213][12] ), .C(\ram[214][12] ), 
        .D(\ram[215][12] ), .S0(n6332), .S1(n6198), .Y(n5693) );
  MX4X1 U5831 ( .A(\ram[228][12] ), .B(\ram[229][12] ), .C(\ram[230][12] ), 
        .D(\ram[231][12] ), .S0(n6332), .S1(n6198), .Y(n5688) );
  MX4X1 U5832 ( .A(\ram[196][12] ), .B(\ram[197][12] ), .C(\ram[198][12] ), 
        .D(\ram[199][12] ), .S0(n6332), .S1(n6198), .Y(n5698) );
  MX4X1 U5833 ( .A(\ram[212][13] ), .B(\ram[213][13] ), .C(\ram[214][13] ), 
        .D(\ram[215][13] ), .S0(n6337), .S1(n6203), .Y(n5777) );
  MX4X1 U5834 ( .A(\ram[228][13] ), .B(\ram[229][13] ), .C(\ram[230][13] ), 
        .D(\ram[231][13] ), .S0(n6337), .S1(n6203), .Y(n5772) );
  MX4X1 U5835 ( .A(\ram[196][13] ), .B(\ram[197][13] ), .C(\ram[198][13] ), 
        .D(\ram[199][13] ), .S0(n6338), .S1(n6204), .Y(n5782) );
  MX4X1 U5836 ( .A(\ram[212][14] ), .B(\ram[213][14] ), .C(\ram[214][14] ), 
        .D(\ram[215][14] ), .S0(n6343), .S1(n6209), .Y(n5861) );
  MX4X1 U5837 ( .A(\ram[228][14] ), .B(\ram[229][14] ), .C(\ram[230][14] ), 
        .D(\ram[231][14] ), .S0(n6342), .S1(n6208), .Y(n5856) );
  MX4X1 U5838 ( .A(\ram[196][14] ), .B(\ram[197][14] ), .C(\ram[198][14] ), 
        .D(\ram[199][14] ), .S0(n6343), .S1(n6209), .Y(n5866) );
  MX4X1 U5839 ( .A(\ram[212][15] ), .B(\ram[213][15] ), .C(\ram[214][15] ), 
        .D(\ram[215][15] ), .S0(n6348), .S1(n6213), .Y(n5945) );
  MX4X1 U5840 ( .A(\ram[228][15] ), .B(\ram[229][15] ), .C(\ram[230][15] ), 
        .D(\ram[231][15] ), .S0(n6348), .S1(n6213), .Y(n5940) );
  MX4X1 U5841 ( .A(\ram[196][15] ), .B(\ram[197][15] ), .C(\ram[198][15] ), 
        .D(\ram[199][15] ), .S0(n6348), .S1(n6213), .Y(n5950) );
  MX4X1 U5842 ( .A(n4707), .B(n4705), .C(n4706), .D(n4704), .S0(n6047), .S1(
        n6057), .Y(n4708) );
  MX4X1 U5843 ( .A(\ram[144][0] ), .B(\ram[145][0] ), .C(\ram[146][0] ), .D(
        \ram[147][0] ), .S0(n6269), .S1(n6135), .Y(n4707) );
  MX4X1 U5844 ( .A(\ram[152][0] ), .B(\ram[153][0] ), .C(\ram[154][0] ), .D(
        \ram[155][0] ), .S0(n6269), .S1(n6135), .Y(n4705) );
  MX4X1 U5845 ( .A(\ram[148][0] ), .B(\ram[149][0] ), .C(\ram[150][0] ), .D(
        \ram[151][0] ), .S0(n6269), .S1(n6135), .Y(n4706) );
  MX4X1 U5846 ( .A(n4749), .B(n4747), .C(n4748), .D(n4746), .S0(n6034), .S1(
        n6067), .Y(n4750) );
  MX4X1 U5847 ( .A(\ram[16][0] ), .B(\ram[17][0] ), .C(\ram[18][0] ), .D(
        \ram[19][0] ), .S0(n6272), .S1(n6138), .Y(n4749) );
  MX4X1 U5848 ( .A(\ram[24][0] ), .B(\ram[25][0] ), .C(\ram[26][0] ), .D(
        \ram[27][0] ), .S0(n6272), .S1(n6138), .Y(n4747) );
  MX4X1 U5849 ( .A(\ram[20][0] ), .B(\ram[21][0] ), .C(\ram[22][0] ), .D(
        \ram[23][0] ), .S0(n6272), .S1(n6138), .Y(n4748) );
  MX4X1 U5850 ( .A(n4812), .B(n4810), .C(n4811), .D(n4809), .S0(n6033), .S1(
        n6056), .Y(n4813) );
  MX4X1 U5851 ( .A(\ram[80][1] ), .B(\ram[81][1] ), .C(\ram[82][1] ), .D(
        \ram[83][1] ), .S0(n6276), .S1(n6142), .Y(n4812) );
  MX4X1 U5852 ( .A(\ram[88][1] ), .B(\ram[89][1] ), .C(\ram[90][1] ), .D(
        \ram[91][1] ), .S0(n6276), .S1(n6142), .Y(n4810) );
  MX4X1 U5853 ( .A(\ram[84][1] ), .B(\ram[85][1] ), .C(\ram[86][1] ), .D(
        \ram[87][1] ), .S0(n6276), .S1(n6142), .Y(n4811) );
  MX4X1 U5854 ( .A(n4791), .B(n4789), .C(n4790), .D(n4788), .S0(n6033), .S1(
        n6056), .Y(n4792) );
  MX4X1 U5855 ( .A(\ram[144][1] ), .B(\ram[145][1] ), .C(\ram[146][1] ), .D(
        \ram[147][1] ), .S0(n6275), .S1(n6141), .Y(n4791) );
  MX4X1 U5856 ( .A(\ram[152][1] ), .B(\ram[153][1] ), .C(\ram[154][1] ), .D(
        \ram[155][1] ), .S0(n6275), .S1(n6141), .Y(n4789) );
  MX4X1 U5857 ( .A(\ram[148][1] ), .B(\ram[149][1] ), .C(\ram[150][1] ), .D(
        \ram[151][1] ), .S0(n6275), .S1(n6141), .Y(n4790) );
  MX4X1 U5858 ( .A(n4833), .B(n4831), .C(n4832), .D(n4830), .S0(n6039), .S1(
        n6057), .Y(n4834) );
  MX4X1 U5859 ( .A(\ram[16][1] ), .B(\ram[17][1] ), .C(\ram[18][1] ), .D(
        \ram[19][1] ), .S0(n6277), .S1(n6143), .Y(n4833) );
  MX4X1 U5860 ( .A(\ram[24][1] ), .B(\ram[25][1] ), .C(\ram[26][1] ), .D(
        \ram[27][1] ), .S0(n6277), .S1(n6143), .Y(n4831) );
  MX4X1 U5861 ( .A(\ram[20][1] ), .B(\ram[21][1] ), .C(\ram[22][1] ), .D(
        \ram[23][1] ), .S0(n6277), .S1(n6143), .Y(n4832) );
  MX4X1 U5862 ( .A(n4896), .B(n4894), .C(n4895), .D(n4893), .S0(n6040), .S1(
        n6058), .Y(n4897) );
  MX4X1 U5863 ( .A(\ram[80][2] ), .B(\ram[81][2] ), .C(\ram[82][2] ), .D(
        \ram[83][2] ), .S0(n6281), .S1(n6147), .Y(n4896) );
  MX4X1 U5864 ( .A(\ram[88][2] ), .B(\ram[89][2] ), .C(\ram[90][2] ), .D(
        \ram[91][2] ), .S0(n6281), .S1(n6147), .Y(n4894) );
  MX4X1 U5865 ( .A(\ram[84][2] ), .B(\ram[85][2] ), .C(\ram[86][2] ), .D(
        \ram[87][2] ), .S0(n6281), .S1(n6147), .Y(n4895) );
  MX4X1 U5866 ( .A(n4875), .B(n4873), .C(n4874), .D(n4872), .S0(n6043), .S1(
        n6057), .Y(n4876) );
  MX4X1 U5867 ( .A(\ram[144][2] ), .B(\ram[145][2] ), .C(\ram[146][2] ), .D(
        \ram[147][2] ), .S0(n6280), .S1(n6146), .Y(n4875) );
  MX4X1 U5868 ( .A(\ram[152][2] ), .B(\ram[153][2] ), .C(\ram[154][2] ), .D(
        \ram[155][2] ), .S0(n6280), .S1(n6146), .Y(n4873) );
  MX4X1 U5869 ( .A(\ram[148][2] ), .B(\ram[149][2] ), .C(\ram[150][2] ), .D(
        \ram[151][2] ), .S0(n6280), .S1(n6146), .Y(n4874) );
  MX4X1 U5870 ( .A(n4917), .B(n4915), .C(n4916), .D(n4914), .S0(n6047), .S1(
        n6058), .Y(n4918) );
  MX4X1 U5871 ( .A(\ram[16][2] ), .B(\ram[17][2] ), .C(\ram[18][2] ), .D(
        \ram[19][2] ), .S0(n6283), .S1(n6149), .Y(n4917) );
  MX4X1 U5872 ( .A(\ram[24][2] ), .B(\ram[25][2] ), .C(\ram[26][2] ), .D(
        \ram[27][2] ), .S0(n6283), .S1(n6149), .Y(n4915) );
  MX4X1 U5873 ( .A(\ram[20][2] ), .B(\ram[21][2] ), .C(\ram[22][2] ), .D(
        \ram[23][2] ), .S0(n6283), .S1(n6149), .Y(n4916) );
  MX4X1 U5874 ( .A(n4980), .B(n4978), .C(n4979), .D(n4977), .S0(n6044), .S1(
        n6059), .Y(n4981) );
  MX4X1 U5875 ( .A(\ram[80][3] ), .B(\ram[81][3] ), .C(\ram[82][3] ), .D(
        \ram[83][3] ), .S0(n6287), .S1(n6153), .Y(n4980) );
  MX4X1 U5876 ( .A(\ram[88][3] ), .B(\ram[89][3] ), .C(\ram[90][3] ), .D(
        \ram[91][3] ), .S0(n6287), .S1(n6153), .Y(n4978) );
  MX4X1 U5877 ( .A(\ram[84][3] ), .B(\ram[85][3] ), .C(\ram[86][3] ), .D(
        \ram[87][3] ), .S0(n6287), .S1(n6153), .Y(n4979) );
  MX4X1 U5878 ( .A(n4938), .B(n4936), .C(n4937), .D(n4935), .S0(n6045), .S1(
        n6058), .Y(n4939) );
  MX4X1 U5879 ( .A(\ram[208][3] ), .B(\ram[209][3] ), .C(\ram[210][3] ), .D(
        \ram[211][3] ), .S0(n6284), .S1(n6150), .Y(n4938) );
  MX4X1 U5880 ( .A(\ram[216][3] ), .B(\ram[217][3] ), .C(\ram[218][3] ), .D(
        \ram[219][3] ), .S0(n6284), .S1(n6150), .Y(n4936) );
  MX4X1 U5881 ( .A(\ram[212][3] ), .B(\ram[213][3] ), .C(\ram[214][3] ), .D(
        \ram[215][3] ), .S0(n6284), .S1(n6150), .Y(n4937) );
  MX4X1 U5882 ( .A(n5001), .B(n4999), .C(n5000), .D(n4998), .S0(n6039), .S1(
        n6059), .Y(n5002) );
  MX4X1 U5883 ( .A(\ram[16][3] ), .B(\ram[17][3] ), .C(\ram[18][3] ), .D(
        \ram[19][3] ), .S0(n6288), .S1(n6154), .Y(n5001) );
  MX4X1 U5884 ( .A(\ram[24][3] ), .B(\ram[25][3] ), .C(\ram[26][3] ), .D(
        \ram[27][3] ), .S0(n6288), .S1(n6154), .Y(n4999) );
  MX4X1 U5885 ( .A(\ram[20][3] ), .B(\ram[21][3] ), .C(\ram[22][3] ), .D(
        \ram[23][3] ), .S0(n6288), .S1(n6154), .Y(n5000) );
  MX4X1 U5886 ( .A(n4959), .B(n4957), .C(n4958), .D(n4956), .S0(n6038), .S1(
        n6059), .Y(n4960) );
  MX4X1 U5887 ( .A(\ram[144][3] ), .B(\ram[145][3] ), .C(\ram[146][3] ), .D(
        \ram[147][3] ), .S0(n6285), .S1(n6151), .Y(n4959) );
  MX4X1 U5888 ( .A(\ram[152][3] ), .B(\ram[153][3] ), .C(\ram[154][3] ), .D(
        \ram[155][3] ), .S0(n6285), .S1(n6151), .Y(n4957) );
  MX4X1 U5889 ( .A(\ram[148][3] ), .B(\ram[149][3] ), .C(\ram[150][3] ), .D(
        \ram[151][3] ), .S0(n6285), .S1(n6151), .Y(n4958) );
  MX4X1 U5890 ( .A(n5064), .B(n5062), .C(n5063), .D(n5061), .S0(n6034), .S1(
        n6060), .Y(n5065) );
  MX4X1 U5891 ( .A(\ram[80][4] ), .B(\ram[81][4] ), .C(\ram[82][4] ), .D(
        \ram[83][4] ), .S0(n6292), .S1(n6158), .Y(n5064) );
  MX4X1 U5892 ( .A(\ram[88][4] ), .B(\ram[89][4] ), .C(\ram[90][4] ), .D(
        \ram[91][4] ), .S0(n6292), .S1(n6158), .Y(n5062) );
  MX4X1 U5893 ( .A(\ram[84][4] ), .B(\ram[85][4] ), .C(\ram[86][4] ), .D(
        \ram[87][4] ), .S0(n6292), .S1(n6158), .Y(n5063) );
  MX4X1 U5894 ( .A(n5043), .B(n5041), .C(n5042), .D(n5040), .S0(n6034), .S1(
        n6060), .Y(n5044) );
  MX4X1 U5895 ( .A(\ram[144][4] ), .B(\ram[145][4] ), .C(\ram[146][4] ), .D(
        \ram[147][4] ), .S0(n6291), .S1(n6157), .Y(n5043) );
  MX4X1 U5896 ( .A(\ram[152][4] ), .B(\ram[153][4] ), .C(\ram[154][4] ), .D(
        \ram[155][4] ), .S0(n6291), .S1(n6157), .Y(n5041) );
  MX4X1 U5897 ( .A(\ram[148][4] ), .B(\ram[149][4] ), .C(\ram[150][4] ), .D(
        \ram[151][4] ), .S0(n6291), .S1(n6157), .Y(n5042) );
  MX4X1 U5898 ( .A(n5085), .B(n5083), .C(n5084), .D(n5082), .S0(n6033), .S1(
        n6061), .Y(n5086) );
  MX4X1 U5899 ( .A(\ram[16][4] ), .B(\ram[17][4] ), .C(\ram[18][4] ), .D(
        \ram[19][4] ), .S0(n6293), .S1(n6159), .Y(n5085) );
  MX4X1 U5900 ( .A(\ram[24][4] ), .B(\ram[25][4] ), .C(\ram[26][4] ), .D(
        \ram[27][4] ), .S0(n6293), .S1(n6159), .Y(n5083) );
  MX4X1 U5901 ( .A(\ram[20][4] ), .B(\ram[21][4] ), .C(\ram[22][4] ), .D(
        \ram[23][4] ), .S0(n6293), .S1(n6159), .Y(n5084) );
  MX4X1 U5902 ( .A(n5148), .B(n5146), .C(n5147), .D(n5145), .S0(n6035), .S1(
        n6062), .Y(n5149) );
  MX4X1 U5903 ( .A(\ram[80][5] ), .B(\ram[81][5] ), .C(\ram[82][5] ), .D(
        \ram[83][5] ), .S0(n6297), .S1(n6163), .Y(n5148) );
  MX4X1 U5904 ( .A(\ram[88][5] ), .B(\ram[89][5] ), .C(\ram[90][5] ), .D(
        \ram[91][5] ), .S0(n6297), .S1(n6163), .Y(n5146) );
  MX4X1 U5905 ( .A(\ram[84][5] ), .B(\ram[85][5] ), .C(\ram[86][5] ), .D(
        \ram[87][5] ), .S0(n6297), .S1(n6163), .Y(n5147) );
  MX4X1 U5906 ( .A(n5127), .B(n5125), .C(n5126), .D(n5124), .S0(n6035), .S1(
        n6061), .Y(n5128) );
  MX4X1 U5907 ( .A(\ram[144][5] ), .B(\ram[145][5] ), .C(\ram[146][5] ), .D(
        \ram[147][5] ), .S0(n6296), .S1(n6162), .Y(n5127) );
  MX4X1 U5908 ( .A(\ram[152][5] ), .B(\ram[153][5] ), .C(\ram[154][5] ), .D(
        \ram[155][5] ), .S0(n6296), .S1(n6162), .Y(n5125) );
  MX4X1 U5909 ( .A(\ram[148][5] ), .B(\ram[149][5] ), .C(\ram[150][5] ), .D(
        \ram[151][5] ), .S0(n6296), .S1(n6162), .Y(n5126) );
  MX4X1 U5910 ( .A(n5169), .B(n5167), .C(n5168), .D(n5166), .S0(n6035), .S1(
        n6062), .Y(n5170) );
  MX4X1 U5911 ( .A(\ram[16][5] ), .B(\ram[17][5] ), .C(\ram[18][5] ), .D(
        \ram[19][5] ), .S0(n6299), .S1(n6165), .Y(n5169) );
  MX4X1 U5912 ( .A(\ram[24][5] ), .B(\ram[25][5] ), .C(\ram[26][5] ), .D(
        \ram[27][5] ), .S0(n6299), .S1(n6165), .Y(n5167) );
  MX4X1 U5913 ( .A(\ram[20][5] ), .B(\ram[21][5] ), .C(\ram[22][5] ), .D(
        \ram[23][5] ), .S0(n6299), .S1(n6165), .Y(n5168) );
  MX4X1 U5914 ( .A(n5232), .B(n5230), .C(n5231), .D(n5229), .S0(n6033), .S1(
        n6063), .Y(n5233) );
  MX4X1 U5915 ( .A(\ram[80][6] ), .B(\ram[81][6] ), .C(\ram[82][6] ), .D(
        \ram[83][6] ), .S0(n6303), .S1(n6169), .Y(n5232) );
  MX4X1 U5916 ( .A(\ram[88][6] ), .B(\ram[89][6] ), .C(\ram[90][6] ), .D(
        \ram[91][6] ), .S0(n6303), .S1(n6169), .Y(n5230) );
  MX4X1 U5917 ( .A(\ram[84][6] ), .B(\ram[85][6] ), .C(\ram[86][6] ), .D(
        \ram[87][6] ), .S0(n6303), .S1(n6169), .Y(n5231) );
  MX4X1 U5918 ( .A(n5211), .B(n5209), .C(n5210), .D(n5208), .S0(n6034), .S1(
        n6063), .Y(n5212) );
  MX4X1 U5919 ( .A(\ram[144][6] ), .B(\ram[145][6] ), .C(\ram[146][6] ), .D(
        \ram[147][6] ), .S0(n6301), .S1(n6167), .Y(n5211) );
  MX4X1 U5920 ( .A(\ram[152][6] ), .B(\ram[153][6] ), .C(\ram[154][6] ), .D(
        \ram[155][6] ), .S0(n6301), .S1(n6167), .Y(n5209) );
  MX4X1 U5921 ( .A(\ram[148][6] ), .B(\ram[149][6] ), .C(\ram[150][6] ), .D(
        \ram[151][6] ), .S0(n6301), .S1(n6167), .Y(n5210) );
  MX4X1 U5922 ( .A(n5253), .B(n5251), .C(n5252), .D(n5250), .S0(n6033), .S1(
        n6063), .Y(n5254) );
  MX4X1 U5923 ( .A(\ram[16][6] ), .B(\ram[17][6] ), .C(\ram[18][6] ), .D(
        \ram[19][6] ), .S0(n6304), .S1(n6170), .Y(n5253) );
  MX4X1 U5924 ( .A(\ram[24][6] ), .B(\ram[25][6] ), .C(\ram[26][6] ), .D(
        \ram[27][6] ), .S0(n6304), .S1(n6170), .Y(n5251) );
  MX4X1 U5925 ( .A(\ram[20][6] ), .B(\ram[21][6] ), .C(\ram[22][6] ), .D(
        \ram[23][6] ), .S0(n6304), .S1(n6170), .Y(n5252) );
  MX4X1 U5926 ( .A(n5316), .B(n5314), .C(n5315), .D(n5313), .S0(n6036), .S1(
        n6064), .Y(n5317) );
  MX4X1 U5927 ( .A(\ram[80][7] ), .B(\ram[81][7] ), .C(\ram[82][7] ), .D(
        \ram[83][7] ), .S0(n6308), .S1(n6174), .Y(n5316) );
  MX4X1 U5928 ( .A(\ram[88][7] ), .B(\ram[89][7] ), .C(\ram[90][7] ), .D(
        \ram[91][7] ), .S0(n6308), .S1(n6174), .Y(n5314) );
  MX4X1 U5929 ( .A(\ram[84][7] ), .B(\ram[85][7] ), .C(\ram[86][7] ), .D(
        \ram[87][7] ), .S0(n6308), .S1(n6174), .Y(n5315) );
  MX4X1 U5930 ( .A(n5295), .B(n5293), .C(n5294), .D(n5292), .S0(n6036), .S1(
        n6064), .Y(n5296) );
  MX4X1 U5931 ( .A(\ram[144][7] ), .B(\ram[145][7] ), .C(\ram[146][7] ), .D(
        \ram[147][7] ), .S0(n6307), .S1(n6173), .Y(n5295) );
  MX4X1 U5932 ( .A(\ram[152][7] ), .B(\ram[153][7] ), .C(\ram[154][7] ), .D(
        \ram[155][7] ), .S0(n6307), .S1(n6173), .Y(n5293) );
  MX4X1 U5933 ( .A(\ram[148][7] ), .B(\ram[149][7] ), .C(\ram[150][7] ), .D(
        \ram[151][7] ), .S0(n6307), .S1(n6173), .Y(n5294) );
  MX4X1 U5934 ( .A(n5337), .B(n5335), .C(n5336), .D(n5334), .S0(n6037), .S1(
        n6065), .Y(n5338) );
  MX4X1 U5935 ( .A(\ram[16][7] ), .B(\ram[17][7] ), .C(\ram[18][7] ), .D(
        \ram[19][7] ), .S0(n6309), .S1(n6175), .Y(n5337) );
  MX4X1 U5936 ( .A(\ram[24][7] ), .B(\ram[25][7] ), .C(\ram[26][7] ), .D(
        \ram[27][7] ), .S0(n6309), .S1(n6175), .Y(n5335) );
  MX4X1 U5937 ( .A(\ram[20][7] ), .B(\ram[21][7] ), .C(\ram[22][7] ), .D(
        \ram[23][7] ), .S0(n6309), .S1(n6175), .Y(n5336) );
  MX4X1 U5938 ( .A(n5400), .B(n5398), .C(n5399), .D(n5397), .S0(n6038), .S1(
        n6066), .Y(n5401) );
  MX4X1 U5939 ( .A(\ram[80][8] ), .B(\ram[81][8] ), .C(\ram[82][8] ), .D(
        \ram[83][8] ), .S0(n6313), .S1(n6179), .Y(n5400) );
  MX4X1 U5940 ( .A(\ram[88][8] ), .B(\ram[89][8] ), .C(\ram[90][8] ), .D(
        \ram[91][8] ), .S0(n6313), .S1(n6179), .Y(n5398) );
  MX4X1 U5941 ( .A(\ram[84][8] ), .B(\ram[85][8] ), .C(\ram[86][8] ), .D(
        \ram[87][8] ), .S0(n6313), .S1(n6179), .Y(n5399) );
  MX4X1 U5942 ( .A(n5379), .B(n5377), .C(n5378), .D(n5376), .S0(n6037), .S1(
        n6065), .Y(n5380) );
  MX4X1 U5943 ( .A(\ram[144][8] ), .B(\ram[145][8] ), .C(\ram[146][8] ), .D(
        \ram[147][8] ), .S0(n6312), .S1(n6178), .Y(n5379) );
  MX4X1 U5944 ( .A(\ram[152][8] ), .B(\ram[153][8] ), .C(\ram[154][8] ), .D(
        \ram[155][8] ), .S0(n6312), .S1(n6178), .Y(n5377) );
  MX4X1 U5945 ( .A(\ram[148][8] ), .B(\ram[149][8] ), .C(\ram[150][8] ), .D(
        \ram[151][8] ), .S0(n6312), .S1(n6178), .Y(n5378) );
  MX4X1 U5946 ( .A(n5421), .B(n5419), .C(n5420), .D(n5418), .S0(n6038), .S1(
        n6066), .Y(n5422) );
  MX4X1 U5947 ( .A(\ram[16][8] ), .B(\ram[17][8] ), .C(\ram[18][8] ), .D(
        \ram[19][8] ), .S0(n6315), .S1(n6181), .Y(n5421) );
  MX4X1 U5948 ( .A(\ram[24][8] ), .B(\ram[25][8] ), .C(\ram[26][8] ), .D(
        \ram[27][8] ), .S0(n6315), .S1(n6181), .Y(n5419) );
  MX4X1 U5949 ( .A(\ram[20][8] ), .B(\ram[21][8] ), .C(\ram[22][8] ), .D(
        \ram[23][8] ), .S0(n6315), .S1(n6181), .Y(n5420) );
  MX4X1 U5950 ( .A(n5484), .B(n5482), .C(n5483), .D(n5481), .S0(n6039), .S1(
        n6067), .Y(n5485) );
  MX4X1 U5951 ( .A(\ram[80][9] ), .B(\ram[81][9] ), .C(\ram[82][9] ), .D(
        \ram[83][9] ), .S0(n6319), .S1(n6185), .Y(n5484) );
  MX4X1 U5952 ( .A(\ram[88][9] ), .B(\ram[89][9] ), .C(\ram[90][9] ), .D(
        \ram[91][9] ), .S0(n6319), .S1(n6185), .Y(n5482) );
  MX4X1 U5953 ( .A(\ram[84][9] ), .B(\ram[85][9] ), .C(\ram[86][9] ), .D(
        \ram[87][9] ), .S0(n6319), .S1(n6185), .Y(n5483) );
  MX4X1 U5954 ( .A(n5463), .B(n5461), .C(n5462), .D(n5460), .S0(n6039), .S1(
        n6067), .Y(n5464) );
  MX4X1 U5955 ( .A(\ram[144][9] ), .B(\ram[145][9] ), .C(\ram[146][9] ), .D(
        \ram[147][9] ), .S0(n6317), .S1(n6183), .Y(n5463) );
  MX4X1 U5956 ( .A(\ram[152][9] ), .B(\ram[153][9] ), .C(\ram[154][9] ), .D(
        \ram[155][9] ), .S0(n6317), .S1(n6183), .Y(n5461) );
  MX4X1 U5957 ( .A(\ram[148][9] ), .B(\ram[149][9] ), .C(\ram[150][9] ), .D(
        \ram[151][9] ), .S0(n6317), .S1(n6183), .Y(n5462) );
  MX4X1 U5958 ( .A(n5505), .B(n5503), .C(n5504), .D(n5502), .S0(n6039), .S1(
        n6067), .Y(n5506) );
  MX4X1 U5959 ( .A(\ram[16][9] ), .B(\ram[17][9] ), .C(\ram[18][9] ), .D(
        \ram[19][9] ), .S0(n6320), .S1(n6186), .Y(n5505) );
  MX4X1 U5960 ( .A(\ram[24][9] ), .B(\ram[25][9] ), .C(\ram[26][9] ), .D(
        \ram[27][9] ), .S0(n6320), .S1(n6186), .Y(n5503) );
  MX4X1 U5961 ( .A(\ram[20][9] ), .B(\ram[21][9] ), .C(\ram[22][9] ), .D(
        \ram[23][9] ), .S0(n6320), .S1(n6186), .Y(n5504) );
  MX4X1 U5962 ( .A(n5547), .B(n5545), .C(n5546), .D(n5544), .S0(n6040), .S1(
        n6068), .Y(n5548) );
  MX4X1 U5963 ( .A(\ram[144][10] ), .B(\ram[145][10] ), .C(\ram[146][10] ), 
        .D(\ram[147][10] ), .S0(n6323), .S1(n6189), .Y(n5547) );
  MX4X1 U5964 ( .A(\ram[152][10] ), .B(\ram[153][10] ), .C(\ram[154][10] ), 
        .D(\ram[155][10] ), .S0(n6323), .S1(n6189), .Y(n5545) );
  MX4X1 U5965 ( .A(\ram[148][10] ), .B(\ram[149][10] ), .C(\ram[150][10] ), 
        .D(\ram[151][10] ), .S0(n6323), .S1(n6189), .Y(n5546) );
  MX4X1 U5966 ( .A(n5568), .B(n5566), .C(n5567), .D(n5565), .S0(n6040), .S1(
        n6068), .Y(n5569) );
  MX4X1 U5967 ( .A(\ram[80][10] ), .B(\ram[81][10] ), .C(\ram[82][10] ), .D(
        \ram[83][10] ), .S0(n6324), .S1(n6190), .Y(n5568) );
  MX4X1 U5968 ( .A(\ram[88][10] ), .B(\ram[89][10] ), .C(\ram[90][10] ), .D(
        \ram[91][10] ), .S0(n6324), .S1(n6190), .Y(n5566) );
  MX4X1 U5969 ( .A(\ram[84][10] ), .B(\ram[85][10] ), .C(\ram[86][10] ), .D(
        \ram[87][10] ), .S0(n6324), .S1(n6190), .Y(n5567) );
  MX4X1 U5970 ( .A(n5589), .B(n5587), .C(n5588), .D(n5586), .S0(n6041), .S1(
        n6069), .Y(n5590) );
  MX4X1 U5971 ( .A(\ram[16][10] ), .B(\ram[17][10] ), .C(\ram[18][10] ), .D(
        \ram[19][10] ), .S0(n6325), .S1(n6191), .Y(n5589) );
  MX4X1 U5972 ( .A(\ram[24][10] ), .B(\ram[25][10] ), .C(\ram[26][10] ), .D(
        \ram[27][10] ), .S0(n6325), .S1(n6191), .Y(n5587) );
  MX4X1 U5973 ( .A(\ram[20][10] ), .B(\ram[21][10] ), .C(\ram[22][10] ), .D(
        \ram[23][10] ), .S0(n6325), .S1(n6191), .Y(n5588) );
  MX4X1 U5974 ( .A(n5652), .B(n5650), .C(n5651), .D(n5649), .S0(n6042), .S1(
        n6070), .Y(n5653) );
  MX4X1 U5975 ( .A(\ram[80][11] ), .B(\ram[81][11] ), .C(\ram[82][11] ), .D(
        \ram[83][11] ), .S0(n6329), .S1(n6195), .Y(n5652) );
  MX4X1 U5976 ( .A(\ram[88][11] ), .B(\ram[89][11] ), .C(\ram[90][11] ), .D(
        \ram[91][11] ), .S0(n6329), .S1(n6195), .Y(n5650) );
  MX4X1 U5977 ( .A(\ram[84][11] ), .B(\ram[85][11] ), .C(\ram[86][11] ), .D(
        \ram[87][11] ), .S0(n6329), .S1(n6195), .Y(n5651) );
  MX4X1 U5978 ( .A(n5631), .B(n5629), .C(n5630), .D(n5628), .S0(n6041), .S1(
        n6069), .Y(n5632) );
  MX4X1 U5979 ( .A(\ram[144][11] ), .B(\ram[145][11] ), .C(\ram[146][11] ), 
        .D(\ram[147][11] ), .S0(n6328), .S1(n6194), .Y(n5631) );
  MX4X1 U5980 ( .A(\ram[152][11] ), .B(\ram[153][11] ), .C(\ram[154][11] ), 
        .D(\ram[155][11] ), .S0(n6328), .S1(n6194), .Y(n5629) );
  MX4X1 U5981 ( .A(\ram[148][11] ), .B(\ram[149][11] ), .C(\ram[150][11] ), 
        .D(\ram[151][11] ), .S0(n6328), .S1(n6194), .Y(n5630) );
  MX4X1 U5982 ( .A(n5673), .B(n5671), .C(n5672), .D(n5670), .S0(n6042), .S1(
        n6070), .Y(n5674) );
  MX4X1 U5983 ( .A(\ram[16][11] ), .B(\ram[17][11] ), .C(\ram[18][11] ), .D(
        \ram[19][11] ), .S0(n6331), .S1(n6197), .Y(n5673) );
  MX4X1 U5984 ( .A(\ram[24][11] ), .B(\ram[25][11] ), .C(\ram[26][11] ), .D(
        \ram[27][11] ), .S0(n6331), .S1(n6197), .Y(n5671) );
  MX4X1 U5985 ( .A(\ram[20][11] ), .B(\ram[21][11] ), .C(\ram[22][11] ), .D(
        \ram[23][11] ), .S0(n6331), .S1(n6197), .Y(n5672) );
  MX4X1 U5986 ( .A(n5736), .B(n5734), .C(n5735), .D(n5733), .S0(n6043), .S1(
        n6071), .Y(n5737) );
  MX4X1 U5987 ( .A(\ram[80][12] ), .B(\ram[81][12] ), .C(\ram[82][12] ), .D(
        \ram[83][12] ), .S0(n6335), .S1(n6201), .Y(n5736) );
  MX4X1 U5988 ( .A(\ram[88][12] ), .B(\ram[89][12] ), .C(\ram[90][12] ), .D(
        \ram[91][12] ), .S0(n6335), .S1(n6201), .Y(n5734) );
  MX4X1 U5989 ( .A(\ram[84][12] ), .B(\ram[85][12] ), .C(\ram[86][12] ), .D(
        \ram[87][12] ), .S0(n6335), .S1(n6201), .Y(n5735) );
  MX4X1 U5990 ( .A(n5715), .B(n5713), .C(n5714), .D(n5712), .S0(n6043), .S1(
        n6071), .Y(n5716) );
  MX4X1 U5991 ( .A(\ram[144][12] ), .B(\ram[145][12] ), .C(\ram[146][12] ), 
        .D(\ram[147][12] ), .S0(n6333), .S1(n6199), .Y(n5715) );
  MX4X1 U5992 ( .A(\ram[152][12] ), .B(\ram[153][12] ), .C(\ram[154][12] ), 
        .D(\ram[155][12] ), .S0(n6333), .S1(n6199), .Y(n5713) );
  MX4X1 U5993 ( .A(\ram[148][12] ), .B(\ram[149][12] ), .C(\ram[150][12] ), 
        .D(\ram[151][12] ), .S0(n6333), .S1(n6199), .Y(n5714) );
  MX4X1 U5994 ( .A(n5757), .B(n5755), .C(n5756), .D(n5754), .S0(n6043), .S1(
        n6071), .Y(n5758) );
  MX4X1 U5995 ( .A(\ram[16][12] ), .B(\ram[17][12] ), .C(\ram[18][12] ), .D(
        \ram[19][12] ), .S0(n6336), .S1(n6202), .Y(n5757) );
  MX4X1 U5996 ( .A(\ram[24][12] ), .B(\ram[25][12] ), .C(\ram[26][12] ), .D(
        \ram[27][12] ), .S0(n6336), .S1(n6202), .Y(n5755) );
  MX4X1 U5997 ( .A(\ram[20][12] ), .B(\ram[21][12] ), .C(\ram[22][12] ), .D(
        \ram[23][12] ), .S0(n6336), .S1(n6202), .Y(n5756) );
  MX4X1 U5998 ( .A(n5820), .B(n5818), .C(n5819), .D(n5817), .S0(n6044), .S1(
        n6072), .Y(n5821) );
  MX4X1 U5999 ( .A(\ram[80][13] ), .B(\ram[81][13] ), .C(\ram[82][13] ), .D(
        \ram[83][13] ), .S0(n6340), .S1(n6206), .Y(n5820) );
  MX4X1 U6000 ( .A(\ram[88][13] ), .B(\ram[89][13] ), .C(\ram[90][13] ), .D(
        \ram[91][13] ), .S0(n6340), .S1(n6206), .Y(n5818) );
  MX4X1 U6001 ( .A(\ram[84][13] ), .B(\ram[85][13] ), .C(\ram[86][13] ), .D(
        \ram[87][13] ), .S0(n6340), .S1(n6206), .Y(n5819) );
  MX4X1 U6002 ( .A(n5799), .B(n5797), .C(n5798), .D(n5796), .S0(n6044), .S1(
        n6072), .Y(n5800) );
  MX4X1 U6003 ( .A(\ram[144][13] ), .B(\ram[145][13] ), .C(\ram[146][13] ), 
        .D(\ram[147][13] ), .S0(n6339), .S1(n6205), .Y(n5799) );
  MX4X1 U6004 ( .A(\ram[152][13] ), .B(\ram[153][13] ), .C(\ram[154][13] ), 
        .D(\ram[155][13] ), .S0(n6339), .S1(n6205), .Y(n5797) );
  MX4X1 U6005 ( .A(\ram[148][13] ), .B(\ram[149][13] ), .C(\ram[150][13] ), 
        .D(\ram[151][13] ), .S0(n6339), .S1(n6205), .Y(n5798) );
  MX4X1 U6006 ( .A(n5841), .B(n5839), .C(n5840), .D(n5838), .S0(n6045), .S1(
        n6073), .Y(n5842) );
  MX4X1 U6007 ( .A(\ram[16][13] ), .B(\ram[17][13] ), .C(\ram[18][13] ), .D(
        \ram[19][13] ), .S0(n6341), .S1(n6207), .Y(n5841) );
  MX4X1 U6008 ( .A(\ram[24][13] ), .B(\ram[25][13] ), .C(\ram[26][13] ), .D(
        \ram[27][13] ), .S0(n6341), .S1(n6207), .Y(n5839) );
  MX4X1 U6009 ( .A(\ram[20][13] ), .B(\ram[21][13] ), .C(\ram[22][13] ), .D(
        \ram[23][13] ), .S0(n6341), .S1(n6207), .Y(n5840) );
  MX4X1 U6010 ( .A(n5904), .B(n5902), .C(n5903), .D(n5901), .S0(n6046), .S1(
        n6063), .Y(n5905) );
  MX4X1 U6011 ( .A(\ram[80][14] ), .B(\ram[81][14] ), .C(\ram[82][14] ), .D(
        \ram[83][14] ), .S0(n6345), .S1(n6211), .Y(n5904) );
  MX4X1 U6012 ( .A(\ram[88][14] ), .B(\ram[89][14] ), .C(\ram[90][14] ), .D(
        \ram[91][14] ), .S0(n6345), .S1(n6211), .Y(n5902) );
  MX4X1 U6013 ( .A(\ram[84][14] ), .B(\ram[85][14] ), .C(\ram[86][14] ), .D(
        \ram[87][14] ), .S0(n6345), .S1(n6211), .Y(n5903) );
  MX4X1 U6014 ( .A(n5883), .B(n5881), .C(n5882), .D(n5880), .S0(n6045), .S1(
        n6073), .Y(n5884) );
  MX4X1 U6015 ( .A(\ram[144][14] ), .B(\ram[145][14] ), .C(\ram[146][14] ), 
        .D(\ram[147][14] ), .S0(n6344), .S1(n6210), .Y(n5883) );
  MX4X1 U6016 ( .A(\ram[152][14] ), .B(\ram[153][14] ), .C(\ram[154][14] ), 
        .D(\ram[155][14] ), .S0(n6344), .S1(n6210), .Y(n5881) );
  MX4X1 U6017 ( .A(\ram[148][14] ), .B(\ram[149][14] ), .C(\ram[150][14] ), 
        .D(\ram[151][14] ), .S0(n6344), .S1(n6210), .Y(n5882) );
  MX4X1 U6018 ( .A(n5925), .B(n5923), .C(n5924), .D(n5922), .S0(n6046), .S1(
        n6063), .Y(n5926) );
  MX4X1 U6019 ( .A(\ram[16][14] ), .B(\ram[17][14] ), .C(\ram[18][14] ), .D(
        \ram[19][14] ), .S0(n6347), .S1(n6213), .Y(n5925) );
  MX4X1 U6020 ( .A(\ram[24][14] ), .B(\ram[25][14] ), .C(\ram[26][14] ), .D(
        \ram[27][14] ), .S0(n6347), .S1(n6214), .Y(n5923) );
  MX4X1 U6021 ( .A(\ram[20][14] ), .B(\ram[21][14] ), .C(\ram[22][14] ), .D(
        \ram[23][14] ), .S0(n6347), .S1(n6213), .Y(n5924) );
  MX4X1 U6022 ( .A(n5988), .B(n5986), .C(n5987), .D(n5985), .S0(n6047), .S1(
        n6061), .Y(n5989) );
  MX4X1 U6023 ( .A(\ram[80][15] ), .B(\ram[81][15] ), .C(\ram[82][15] ), .D(
        \ram[83][15] ), .S0(n6351), .S1(n6194), .Y(n5988) );
  MX4X1 U6024 ( .A(\ram[88][15] ), .B(\ram[89][15] ), .C(\ram[90][15] ), .D(
        \ram[91][15] ), .S0(n6351), .S1(n6191), .Y(n5986) );
  MX4X1 U6025 ( .A(\ram[84][15] ), .B(\ram[85][15] ), .C(\ram[86][15] ), .D(
        \ram[87][15] ), .S0(n6351), .S1(n6193), .Y(n5987) );
  MX4X1 U6026 ( .A(n5967), .B(n5965), .C(n5966), .D(n5964), .S0(n6047), .S1(
        n6073), .Y(n5968) );
  MX4X1 U6027 ( .A(\ram[144][15] ), .B(\ram[145][15] ), .C(\ram[146][15] ), 
        .D(\ram[147][15] ), .S0(n6349), .S1(n6214), .Y(n5967) );
  MX4X1 U6028 ( .A(\ram[152][15] ), .B(\ram[153][15] ), .C(\ram[154][15] ), 
        .D(\ram[155][15] ), .S0(n6349), .S1(n6214), .Y(n5965) );
  MX4X1 U6029 ( .A(\ram[148][15] ), .B(\ram[149][15] ), .C(\ram[150][15] ), 
        .D(\ram[151][15] ), .S0(n6349), .S1(n6214), .Y(n5966) );
  MX4X1 U6030 ( .A(n6009), .B(n6007), .C(n6008), .D(n6006), .S0(n6047), .S1(
        n6060), .Y(n6010) );
  MX4X1 U6031 ( .A(\ram[16][15] ), .B(\ram[17][15] ), .C(\ram[18][15] ), .D(
        \ram[19][15] ), .S0(n6352), .S1(n6214), .Y(n6009) );
  MX4X1 U6032 ( .A(\ram[24][15] ), .B(\ram[25][15] ), .C(\ram[26][15] ), .D(
        \ram[27][15] ), .S0(n6352), .S1(n6140), .Y(n6007) );
  MX4X1 U6033 ( .A(\ram[20][15] ), .B(\ram[21][15] ), .C(\ram[22][15] ), .D(
        \ram[23][15] ), .S0(n6352), .S1(n6213), .Y(n6008) );
  MX4X1 U6034 ( .A(\ram[80][0] ), .B(\ram[81][0] ), .C(\ram[82][0] ), .D(
        \ram[83][0] ), .S0(n6271), .S1(n6137), .Y(n4728) );
  MX4X1 U6035 ( .A(\ram[96][0] ), .B(\ram[97][0] ), .C(\ram[98][0] ), .D(
        \ram[99][0] ), .S0(n6270), .S1(n6136), .Y(n4723) );
  MX4X1 U6036 ( .A(\ram[64][0] ), .B(\ram[65][0] ), .C(\ram[66][0] ), .D(
        \ram[67][0] ), .S0(n6271), .S1(n6137), .Y(n4733) );
  MX4X1 U6037 ( .A(\ram[208][1] ), .B(\ram[209][1] ), .C(\ram[210][1] ), .D(
        \ram[211][1] ), .S0(n6273), .S1(n6139), .Y(n4770) );
  MX4X1 U6038 ( .A(\ram[224][1] ), .B(\ram[225][1] ), .C(\ram[226][1] ), .D(
        \ram[227][1] ), .S0(n6273), .S1(n6139), .Y(n4765) );
  MX4X1 U6039 ( .A(\ram[192][1] ), .B(\ram[193][1] ), .C(\ram[194][1] ), .D(
        \ram[195][1] ), .S0(n6274), .S1(n6140), .Y(n4775) );
  MX4X1 U6040 ( .A(\ram[208][2] ), .B(\ram[209][2] ), .C(\ram[210][2] ), .D(
        \ram[211][2] ), .S0(n6279), .S1(n6145), .Y(n4854) );
  MX4X1 U6041 ( .A(\ram[224][2] ), .B(\ram[225][2] ), .C(\ram[226][2] ), .D(
        \ram[227][2] ), .S0(n6278), .S1(n6144), .Y(n4849) );
  MX4X1 U6042 ( .A(\ram[192][2] ), .B(\ram[193][2] ), .C(\ram[194][2] ), .D(
        \ram[195][2] ), .S0(n6279), .S1(n6145), .Y(n4859) );
  MX4X1 U6043 ( .A(\ram[112][3] ), .B(\ram[113][3] ), .C(\ram[114][3] ), .D(
        \ram[115][3] ), .S0(n6286), .S1(n6152), .Y(n4970) );
  MX4X1 U6044 ( .A(\ram[64][3] ), .B(\ram[65][3] ), .C(\ram[66][3] ), .D(
        \ram[67][3] ), .S0(n6287), .S1(n6153), .Y(n4985) );
  MX4X1 U6045 ( .A(\ram[96][3] ), .B(\ram[97][3] ), .C(\ram[98][3] ), .D(
        \ram[99][3] ), .S0(n6286), .S1(n6152), .Y(n4975) );
  MX4X1 U6046 ( .A(\ram[208][4] ), .B(\ram[209][4] ), .C(\ram[210][4] ), .D(
        \ram[211][4] ), .S0(n6289), .S1(n6155), .Y(n5022) );
  MX4X1 U6047 ( .A(\ram[224][4] ), .B(\ram[225][4] ), .C(\ram[226][4] ), .D(
        \ram[227][4] ), .S0(n6289), .S1(n6155), .Y(n5017) );
  MX4X1 U6048 ( .A(\ram[192][4] ), .B(\ram[193][4] ), .C(\ram[194][4] ), .D(
        \ram[195][4] ), .S0(n6290), .S1(n6156), .Y(n5027) );
  MX4X1 U6049 ( .A(\ram[208][5] ), .B(\ram[209][5] ), .C(\ram[210][5] ), .D(
        \ram[211][5] ), .S0(n6295), .S1(n6161), .Y(n5106) );
  MX4X1 U6050 ( .A(\ram[224][5] ), .B(\ram[225][5] ), .C(\ram[226][5] ), .D(
        \ram[227][5] ), .S0(n6294), .S1(n6160), .Y(n5101) );
  MX4X1 U6051 ( .A(\ram[192][5] ), .B(\ram[193][5] ), .C(\ram[194][5] ), .D(
        \ram[195][5] ), .S0(n6295), .S1(n6161), .Y(n5111) );
  MX4X1 U6052 ( .A(\ram[208][6] ), .B(\ram[209][6] ), .C(\ram[210][6] ), .D(
        \ram[211][6] ), .S0(n6300), .S1(n6166), .Y(n5190) );
  MX4X1 U6053 ( .A(\ram[224][6] ), .B(\ram[225][6] ), .C(\ram[226][6] ), .D(
        \ram[227][6] ), .S0(n6300), .S1(n6166), .Y(n5185) );
  MX4X1 U6054 ( .A(\ram[192][6] ), .B(\ram[193][6] ), .C(\ram[194][6] ), .D(
        \ram[195][6] ), .S0(n6300), .S1(n6166), .Y(n5195) );
  MX4X1 U6055 ( .A(\ram[208][7] ), .B(\ram[209][7] ), .C(\ram[210][7] ), .D(
        \ram[211][7] ), .S0(n6305), .S1(n6171), .Y(n5274) );
  MX4X1 U6056 ( .A(\ram[224][7] ), .B(\ram[225][7] ), .C(\ram[226][7] ), .D(
        \ram[227][7] ), .S0(n6305), .S1(n6171), .Y(n5269) );
  MX4X1 U6057 ( .A(\ram[192][7] ), .B(\ram[193][7] ), .C(\ram[194][7] ), .D(
        \ram[195][7] ), .S0(n6306), .S1(n6172), .Y(n5279) );
  MX4X1 U6058 ( .A(\ram[208][8] ), .B(\ram[209][8] ), .C(\ram[210][8] ), .D(
        \ram[211][8] ), .S0(n6311), .S1(n6177), .Y(n5358) );
  MX4X1 U6059 ( .A(\ram[224][8] ), .B(\ram[225][8] ), .C(\ram[226][8] ), .D(
        \ram[227][8] ), .S0(n6310), .S1(n6176), .Y(n5353) );
  MX4X1 U6060 ( .A(\ram[192][8] ), .B(\ram[193][8] ), .C(\ram[194][8] ), .D(
        \ram[195][8] ), .S0(n6311), .S1(n6177), .Y(n5363) );
  MX4X1 U6061 ( .A(\ram[208][9] ), .B(\ram[209][9] ), .C(\ram[210][9] ), .D(
        \ram[211][9] ), .S0(n6316), .S1(n6182), .Y(n5442) );
  MX4X1 U6062 ( .A(\ram[224][9] ), .B(\ram[225][9] ), .C(\ram[226][9] ), .D(
        \ram[227][9] ), .S0(n6316), .S1(n6182), .Y(n5437) );
  MX4X1 U6063 ( .A(\ram[192][9] ), .B(\ram[193][9] ), .C(\ram[194][9] ), .D(
        \ram[195][9] ), .S0(n6316), .S1(n6182), .Y(n5447) );
  MX4X1 U6064 ( .A(\ram[208][10] ), .B(\ram[209][10] ), .C(\ram[210][10] ), 
        .D(\ram[211][10] ), .S0(n6321), .S1(n6187), .Y(n5526) );
  MX4X1 U6065 ( .A(\ram[224][10] ), .B(\ram[225][10] ), .C(\ram[226][10] ), 
        .D(\ram[227][10] ), .S0(n6321), .S1(n6187), .Y(n5521) );
  MX4X1 U6066 ( .A(\ram[192][10] ), .B(\ram[193][10] ), .C(\ram[194][10] ), 
        .D(\ram[195][10] ), .S0(n6322), .S1(n6188), .Y(n5531) );
  MX4X1 U6067 ( .A(\ram[208][11] ), .B(\ram[209][11] ), .C(\ram[210][11] ), 
        .D(\ram[211][11] ), .S0(n6327), .S1(n6193), .Y(n5610) );
  MX4X1 U6068 ( .A(\ram[224][11] ), .B(\ram[225][11] ), .C(\ram[226][11] ), 
        .D(\ram[227][11] ), .S0(n6326), .S1(n6192), .Y(n5605) );
  MX4X1 U6069 ( .A(\ram[192][11] ), .B(\ram[193][11] ), .C(\ram[194][11] ), 
        .D(\ram[195][11] ), .S0(n6327), .S1(n6193), .Y(n5615) );
  MX4X1 U6070 ( .A(\ram[208][12] ), .B(\ram[209][12] ), .C(\ram[210][12] ), 
        .D(\ram[211][12] ), .S0(n6332), .S1(n6198), .Y(n5694) );
  MX4X1 U6071 ( .A(\ram[224][12] ), .B(\ram[225][12] ), .C(\ram[226][12] ), 
        .D(\ram[227][12] ), .S0(n6332), .S1(n6198), .Y(n5689) );
  MX4X1 U6072 ( .A(\ram[192][12] ), .B(\ram[193][12] ), .C(\ram[194][12] ), 
        .D(\ram[195][12] ), .S0(n6332), .S1(n6198), .Y(n5699) );
  MX4X1 U6073 ( .A(\ram[208][13] ), .B(\ram[209][13] ), .C(\ram[210][13] ), 
        .D(\ram[211][13] ), .S0(n6337), .S1(n6203), .Y(n5778) );
  MX4X1 U6074 ( .A(\ram[224][13] ), .B(\ram[225][13] ), .C(\ram[226][13] ), 
        .D(\ram[227][13] ), .S0(n6337), .S1(n6203), .Y(n5773) );
  MX4X1 U6075 ( .A(\ram[192][13] ), .B(\ram[193][13] ), .C(\ram[194][13] ), 
        .D(\ram[195][13] ), .S0(n6338), .S1(n6204), .Y(n5783) );
  MX4X1 U6076 ( .A(\ram[208][14] ), .B(\ram[209][14] ), .C(\ram[210][14] ), 
        .D(\ram[211][14] ), .S0(n6343), .S1(n6209), .Y(n5862) );
  MX4X1 U6077 ( .A(\ram[224][14] ), .B(\ram[225][14] ), .C(\ram[226][14] ), 
        .D(\ram[227][14] ), .S0(n6342), .S1(n6208), .Y(n5857) );
  MX4X1 U6078 ( .A(\ram[192][14] ), .B(\ram[193][14] ), .C(\ram[194][14] ), 
        .D(\ram[195][14] ), .S0(n6343), .S1(n6209), .Y(n5867) );
  MX4X1 U6079 ( .A(\ram[208][15] ), .B(\ram[209][15] ), .C(\ram[210][15] ), 
        .D(\ram[211][15] ), .S0(n6348), .S1(n6213), .Y(n5946) );
  MX4X1 U6080 ( .A(\ram[224][15] ), .B(\ram[225][15] ), .C(\ram[226][15] ), 
        .D(\ram[227][15] ), .S0(n6348), .S1(n6213), .Y(n5941) );
  MX4X1 U6081 ( .A(\ram[192][15] ), .B(\ram[193][15] ), .C(\ram[194][15] ), 
        .D(\ram[195][15] ), .S0(n6348), .S1(n6213), .Y(n5951) );
  MX4X1 U6082 ( .A(n4712), .B(n4710), .C(n4711), .D(n4709), .S0(n6039), .S1(
        n6063), .Y(n4713) );
  MX4X1 U6083 ( .A(\ram[128][0] ), .B(\ram[129][0] ), .C(\ram[130][0] ), .D(
        \ram[131][0] ), .S0(n6270), .S1(n6136), .Y(n4712) );
  MX4X1 U6084 ( .A(\ram[136][0] ), .B(\ram[137][0] ), .C(\ram[138][0] ), .D(
        \ram[139][0] ), .S0(n6270), .S1(n6136), .Y(n4710) );
  MX4X1 U6085 ( .A(\ram[132][0] ), .B(\ram[133][0] ), .C(\ram[134][0] ), .D(
        \ram[135][0] ), .S0(n6270), .S1(n6136), .Y(n4711) );
  MX4X1 U6086 ( .A(n4754), .B(n4752), .C(n4753), .D(n4751), .S0(n6047), .S1(
        n6064), .Y(n4755) );
  MX4X1 U6087 ( .A(\ram[0][0] ), .B(\ram[1][0] ), .C(\ram[2][0] ), .D(
        \ram[3][0] ), .S0(n6272), .S1(n6138), .Y(n4754) );
  MX4X1 U6088 ( .A(\ram[8][0] ), .B(\ram[9][0] ), .C(\ram[10][0] ), .D(
        \ram[11][0] ), .S0(n6272), .S1(n6138), .Y(n4752) );
  MX4X1 U6089 ( .A(\ram[4][0] ), .B(\ram[5][0] ), .C(\ram[6][0] ), .D(
        \ram[7][0] ), .S0(n6272), .S1(n6138), .Y(n4753) );
  MX4X1 U6090 ( .A(n4817), .B(n4815), .C(n4816), .D(n4814), .S0(n6033), .S1(
        n6056), .Y(n4818) );
  MX4X1 U6091 ( .A(\ram[64][1] ), .B(\ram[65][1] ), .C(\ram[66][1] ), .D(
        \ram[67][1] ), .S0(n6276), .S1(n6142), .Y(n4817) );
  MX4X1 U6092 ( .A(\ram[72][1] ), .B(\ram[73][1] ), .C(\ram[74][1] ), .D(
        \ram[75][1] ), .S0(n6276), .S1(n6142), .Y(n4815) );
  MX4X1 U6093 ( .A(\ram[68][1] ), .B(\ram[69][1] ), .C(\ram[70][1] ), .D(
        \ram[71][1] ), .S0(n6276), .S1(n6142), .Y(n4816) );
  MX4X1 U6094 ( .A(n4796), .B(n4794), .C(n4795), .D(n4793), .S0(n6033), .S1(
        n6056), .Y(n4797) );
  MX4X1 U6095 ( .A(\ram[128][1] ), .B(\ram[129][1] ), .C(\ram[130][1] ), .D(
        \ram[131][1] ), .S0(n6275), .S1(n6141), .Y(n4796) );
  MX4X1 U6096 ( .A(\ram[136][1] ), .B(\ram[137][1] ), .C(\ram[138][1] ), .D(
        \ram[139][1] ), .S0(n6275), .S1(n6141), .Y(n4794) );
  MX4X1 U6097 ( .A(\ram[132][1] ), .B(\ram[133][1] ), .C(\ram[134][1] ), .D(
        \ram[135][1] ), .S0(n6275), .S1(n6141), .Y(n4795) );
  MX4X1 U6098 ( .A(n4838), .B(n4836), .C(n4837), .D(n4835), .S0(n6045), .S1(
        n6057), .Y(n4839) );
  MX4X1 U6099 ( .A(\ram[0][1] ), .B(\ram[1][1] ), .C(\ram[2][1] ), .D(
        \ram[3][1] ), .S0(n6278), .S1(n6144), .Y(n4838) );
  MX4X1 U6100 ( .A(\ram[8][1] ), .B(\ram[9][1] ), .C(\ram[10][1] ), .D(
        \ram[11][1] ), .S0(n6278), .S1(n6144), .Y(n4836) );
  MX4X1 U6101 ( .A(\ram[4][1] ), .B(\ram[5][1] ), .C(\ram[6][1] ), .D(
        \ram[7][1] ), .S0(n6278), .S1(n6144), .Y(n4837) );
  MX4X1 U6102 ( .A(n4901), .B(n4899), .C(n4900), .D(n4898), .S0(n6039), .S1(
        n6058), .Y(n4902) );
  MX4X1 U6103 ( .A(\ram[64][2] ), .B(\ram[65][2] ), .C(\ram[66][2] ), .D(
        \ram[67][2] ), .S0(n6282), .S1(n6148), .Y(n4901) );
  MX4X1 U6104 ( .A(\ram[72][2] ), .B(\ram[73][2] ), .C(\ram[74][2] ), .D(
        \ram[75][2] ), .S0(n6282), .S1(n6148), .Y(n4899) );
  MX4X1 U6105 ( .A(\ram[68][2] ), .B(\ram[69][2] ), .C(\ram[70][2] ), .D(
        \ram[71][2] ), .S0(n6282), .S1(n6148), .Y(n4900) );
  MX4X1 U6106 ( .A(n4880), .B(n4878), .C(n4879), .D(n4877), .S0(n6041), .S1(
        n6057), .Y(n4881) );
  MX4X1 U6107 ( .A(\ram[128][2] ), .B(\ram[129][2] ), .C(\ram[130][2] ), .D(
        \ram[131][2] ), .S0(n6280), .S1(n6146), .Y(n4880) );
  MX4X1 U6108 ( .A(\ram[136][2] ), .B(\ram[137][2] ), .C(\ram[138][2] ), .D(
        \ram[139][2] ), .S0(n6280), .S1(n6146), .Y(n4878) );
  MX4X1 U6109 ( .A(\ram[132][2] ), .B(\ram[133][2] ), .C(\ram[134][2] ), .D(
        \ram[135][2] ), .S0(n6280), .S1(n6146), .Y(n4879) );
  MX4X1 U6110 ( .A(n4922), .B(n4920), .C(n4921), .D(n4919), .S0(n6043), .S1(
        n6058), .Y(n4923) );
  MX4X1 U6111 ( .A(\ram[0][2] ), .B(\ram[1][2] ), .C(\ram[2][2] ), .D(
        \ram[3][2] ), .S0(n6283), .S1(n6149), .Y(n4922) );
  MX4X1 U6112 ( .A(\ram[8][2] ), .B(\ram[9][2] ), .C(\ram[10][2] ), .D(
        \ram[11][2] ), .S0(n6283), .S1(n6149), .Y(n4920) );
  MX4X1 U6113 ( .A(\ram[4][2] ), .B(\ram[5][2] ), .C(\ram[6][2] ), .D(
        \ram[7][2] ), .S0(n6283), .S1(n6149), .Y(n4921) );
  MX4X1 U6114 ( .A(n4943), .B(n4941), .C(n4942), .D(n4940), .S0(n6043), .S1(
        n6058), .Y(n4944) );
  MX4X1 U6115 ( .A(\ram[192][3] ), .B(\ram[193][3] ), .C(\ram[194][3] ), .D(
        \ram[195][3] ), .S0(n6284), .S1(n6150), .Y(n4943) );
  MX4X1 U6116 ( .A(\ram[200][3] ), .B(\ram[201][3] ), .C(\ram[202][3] ), .D(
        \ram[203][3] ), .S0(n6284), .S1(n6150), .Y(n4941) );
  MX4X1 U6117 ( .A(\ram[196][3] ), .B(\ram[197][3] ), .C(\ram[198][3] ), .D(
        \ram[199][3] ), .S0(n6284), .S1(n6150), .Y(n4942) );
  MX4X1 U6118 ( .A(n5006), .B(n5004), .C(n5005), .D(n5003), .S0(n6049), .S1(
        n6059), .Y(n5007) );
  MX4X1 U6119 ( .A(\ram[0][3] ), .B(\ram[1][3] ), .C(\ram[2][3] ), .D(
        \ram[3][3] ), .S0(n6288), .S1(n6154), .Y(n5006) );
  MX4X1 U6120 ( .A(\ram[8][3] ), .B(\ram[9][3] ), .C(\ram[10][3] ), .D(
        \ram[11][3] ), .S0(n6288), .S1(n6154), .Y(n5004) );
  MX4X1 U6121 ( .A(\ram[4][3] ), .B(\ram[5][3] ), .C(\ram[6][3] ), .D(
        \ram[7][3] ), .S0(n6288), .S1(n6154), .Y(n5005) );
  MX4X1 U6122 ( .A(n4964), .B(n4962), .C(n4963), .D(n4961), .S0(n6025), .S1(
        n6059), .Y(n4965) );
  MX4X1 U6123 ( .A(\ram[128][3] ), .B(\ram[129][3] ), .C(\ram[130][3] ), .D(
        \ram[131][3] ), .S0(n6286), .S1(n6152), .Y(n4964) );
  MX4X1 U6124 ( .A(\ram[136][3] ), .B(\ram[137][3] ), .C(\ram[138][3] ), .D(
        \ram[139][3] ), .S0(n6286), .S1(n6152), .Y(n4962) );
  MX4X1 U6125 ( .A(\ram[132][3] ), .B(\ram[133][3] ), .C(\ram[134][3] ), .D(
        \ram[135][3] ), .S0(n6286), .S1(n6152), .Y(n4963) );
  MX4X1 U6126 ( .A(n5069), .B(n5067), .C(n5068), .D(n5066), .S0(n6034), .S1(
        n6060), .Y(n5070) );
  MX4X1 U6127 ( .A(\ram[64][4] ), .B(\ram[65][4] ), .C(\ram[66][4] ), .D(
        \ram[67][4] ), .S0(n6292), .S1(n6158), .Y(n5069) );
  MX4X1 U6128 ( .A(\ram[72][4] ), .B(\ram[73][4] ), .C(\ram[74][4] ), .D(
        \ram[75][4] ), .S0(n6292), .S1(n6158), .Y(n5067) );
  MX4X1 U6129 ( .A(\ram[68][4] ), .B(\ram[69][4] ), .C(\ram[70][4] ), .D(
        \ram[71][4] ), .S0(n6292), .S1(n6158), .Y(n5068) );
  MX4X1 U6130 ( .A(n5048), .B(n5046), .C(n5047), .D(n5045), .S0(n6034), .S1(
        n6060), .Y(n5049) );
  MX4X1 U6131 ( .A(\ram[128][4] ), .B(\ram[129][4] ), .C(\ram[130][4] ), .D(
        \ram[131][4] ), .S0(n6291), .S1(n6157), .Y(n5048) );
  MX4X1 U6132 ( .A(\ram[136][4] ), .B(\ram[137][4] ), .C(\ram[138][4] ), .D(
        \ram[139][4] ), .S0(n6291), .S1(n6157), .Y(n5046) );
  MX4X1 U6133 ( .A(\ram[132][4] ), .B(\ram[133][4] ), .C(\ram[134][4] ), .D(
        \ram[135][4] ), .S0(n6291), .S1(n6157), .Y(n5047) );
  MX4X1 U6134 ( .A(n5090), .B(n5088), .C(n5089), .D(n5087), .S0(n6045), .S1(
        n6061), .Y(n5091) );
  MX4X1 U6135 ( .A(\ram[0][4] ), .B(\ram[1][4] ), .C(\ram[2][4] ), .D(
        \ram[3][4] ), .S0(n6294), .S1(n6160), .Y(n5090) );
  MX4X1 U6136 ( .A(\ram[8][4] ), .B(\ram[9][4] ), .C(\ram[10][4] ), .D(
        \ram[11][4] ), .S0(n6294), .S1(n6160), .Y(n5088) );
  MX4X1 U6137 ( .A(\ram[4][4] ), .B(\ram[5][4] ), .C(\ram[6][4] ), .D(
        \ram[7][4] ), .S0(n6294), .S1(n6160), .Y(n5089) );
  MX4X1 U6138 ( .A(n5153), .B(n5151), .C(n5152), .D(n5150), .S0(n6035), .S1(
        n6062), .Y(n5154) );
  MX4X1 U6139 ( .A(\ram[64][5] ), .B(\ram[65][5] ), .C(\ram[66][5] ), .D(
        \ram[67][5] ), .S0(n6298), .S1(n6164), .Y(n5153) );
  MX4X1 U6140 ( .A(\ram[72][5] ), .B(\ram[73][5] ), .C(\ram[74][5] ), .D(
        \ram[75][5] ), .S0(n6298), .S1(n6164), .Y(n5151) );
  MX4X1 U6141 ( .A(\ram[68][5] ), .B(\ram[69][5] ), .C(\ram[70][5] ), .D(
        \ram[71][5] ), .S0(n6298), .S1(n6164), .Y(n5152) );
  MX4X1 U6142 ( .A(n5132), .B(n5130), .C(n5131), .D(n5129), .S0(n6033), .S1(
        n6061), .Y(n5133) );
  MX4X1 U6143 ( .A(\ram[128][5] ), .B(\ram[129][5] ), .C(\ram[130][5] ), .D(
        \ram[131][5] ), .S0(n6296), .S1(n6162), .Y(n5132) );
  MX4X1 U6144 ( .A(\ram[136][5] ), .B(\ram[137][5] ), .C(\ram[138][5] ), .D(
        \ram[139][5] ), .S0(n6296), .S1(n6162), .Y(n5130) );
  MX4X1 U6145 ( .A(\ram[132][5] ), .B(\ram[133][5] ), .C(\ram[134][5] ), .D(
        \ram[135][5] ), .S0(n6296), .S1(n6162), .Y(n5131) );
  MX4X1 U6146 ( .A(n5174), .B(n5172), .C(n5173), .D(n5171), .S0(n6035), .S1(
        n6062), .Y(n5175) );
  MX4X1 U6147 ( .A(\ram[0][5] ), .B(\ram[1][5] ), .C(\ram[2][5] ), .D(
        \ram[3][5] ), .S0(n6299), .S1(n6165), .Y(n5174) );
  MX4X1 U6148 ( .A(\ram[8][5] ), .B(\ram[9][5] ), .C(\ram[10][5] ), .D(
        \ram[11][5] ), .S0(n6299), .S1(n6165), .Y(n5172) );
  MX4X1 U6149 ( .A(\ram[4][5] ), .B(\ram[5][5] ), .C(\ram[6][5] ), .D(
        \ram[7][5] ), .S0(n6299), .S1(n6165), .Y(n5173) );
  MX4X1 U6150 ( .A(n5237), .B(n5235), .C(n5236), .D(n5234), .S0(n6042), .S1(
        n6063), .Y(n5238) );
  MX4X1 U6151 ( .A(\ram[64][6] ), .B(\ram[65][6] ), .C(\ram[66][6] ), .D(
        \ram[67][6] ), .S0(n6303), .S1(n6169), .Y(n5237) );
  MX4X1 U6152 ( .A(\ram[72][6] ), .B(\ram[73][6] ), .C(\ram[74][6] ), .D(
        \ram[75][6] ), .S0(n6303), .S1(n6169), .Y(n5235) );
  MX4X1 U6153 ( .A(\ram[68][6] ), .B(\ram[69][6] ), .C(\ram[70][6] ), .D(
        \ram[71][6] ), .S0(n6303), .S1(n6169), .Y(n5236) );
  MX4X1 U6154 ( .A(n5216), .B(n5214), .C(n5215), .D(n5213), .S0(n6037), .S1(
        n6063), .Y(n5217) );
  MX4X1 U6155 ( .A(\ram[128][6] ), .B(\ram[129][6] ), .C(\ram[130][6] ), .D(
        \ram[131][6] ), .S0(n6302), .S1(n6168), .Y(n5216) );
  MX4X1 U6156 ( .A(\ram[136][6] ), .B(\ram[137][6] ), .C(\ram[138][6] ), .D(
        \ram[139][6] ), .S0(n6302), .S1(n6168), .Y(n5214) );
  MX4X1 U6157 ( .A(\ram[132][6] ), .B(\ram[133][6] ), .C(\ram[134][6] ), .D(
        \ram[135][6] ), .S0(n6302), .S1(n6168), .Y(n5215) );
  MX4X1 U6158 ( .A(n5258), .B(n5256), .C(n5257), .D(n5255), .S0(n6034), .S1(
        n6063), .Y(n5259) );
  MX4X1 U6159 ( .A(\ram[0][6] ), .B(\ram[1][6] ), .C(\ram[2][6] ), .D(
        \ram[3][6] ), .S0(n6304), .S1(n6170), .Y(n5258) );
  MX4X1 U6160 ( .A(\ram[8][6] ), .B(\ram[9][6] ), .C(\ram[10][6] ), .D(
        \ram[11][6] ), .S0(n6304), .S1(n6170), .Y(n5256) );
  MX4X1 U6161 ( .A(\ram[4][6] ), .B(\ram[5][6] ), .C(\ram[6][6] ), .D(
        \ram[7][6] ), .S0(n6304), .S1(n6170), .Y(n5257) );
  MX4X1 U6162 ( .A(n5321), .B(n5319), .C(n5320), .D(n5318), .S0(n6036), .S1(
        n6064), .Y(n5322) );
  MX4X1 U6163 ( .A(\ram[64][7] ), .B(\ram[65][7] ), .C(\ram[66][7] ), .D(
        \ram[67][7] ), .S0(n6308), .S1(n6174), .Y(n5321) );
  MX4X1 U6164 ( .A(\ram[72][7] ), .B(\ram[73][7] ), .C(\ram[74][7] ), .D(
        \ram[75][7] ), .S0(n6308), .S1(n6174), .Y(n5319) );
  MX4X1 U6165 ( .A(\ram[68][7] ), .B(\ram[69][7] ), .C(\ram[70][7] ), .D(
        \ram[71][7] ), .S0(n6308), .S1(n6174), .Y(n5320) );
  MX4X1 U6166 ( .A(n5300), .B(n5298), .C(n5299), .D(n5297), .S0(n6036), .S1(
        n6064), .Y(n5301) );
  MX4X1 U6167 ( .A(\ram[128][7] ), .B(\ram[129][7] ), .C(\ram[130][7] ), .D(
        \ram[131][7] ), .S0(n6307), .S1(n6173), .Y(n5300) );
  MX4X1 U6168 ( .A(\ram[136][7] ), .B(\ram[137][7] ), .C(\ram[138][7] ), .D(
        \ram[139][7] ), .S0(n6307), .S1(n6173), .Y(n5298) );
  MX4X1 U6169 ( .A(\ram[132][7] ), .B(\ram[133][7] ), .C(\ram[134][7] ), .D(
        \ram[135][7] ), .S0(n6307), .S1(n6173), .Y(n5299) );
  MX4X1 U6170 ( .A(n5342), .B(n5340), .C(n5341), .D(n5339), .S0(n6037), .S1(
        n6065), .Y(n5343) );
  MX4X1 U6171 ( .A(\ram[0][7] ), .B(\ram[1][7] ), .C(\ram[2][7] ), .D(
        \ram[3][7] ), .S0(n6310), .S1(n6176), .Y(n5342) );
  MX4X1 U6172 ( .A(\ram[8][7] ), .B(\ram[9][7] ), .C(\ram[10][7] ), .D(
        \ram[11][7] ), .S0(n6310), .S1(n6176), .Y(n5340) );
  MX4X1 U6173 ( .A(\ram[4][7] ), .B(\ram[5][7] ), .C(\ram[6][7] ), .D(
        \ram[7][7] ), .S0(n6310), .S1(n6176), .Y(n5341) );
  MX4X1 U6174 ( .A(n5405), .B(n5403), .C(n5404), .D(n5402), .S0(n6038), .S1(
        n6066), .Y(n5406) );
  MX4X1 U6175 ( .A(\ram[64][8] ), .B(\ram[65][8] ), .C(\ram[66][8] ), .D(
        \ram[67][8] ), .S0(n6314), .S1(n6180), .Y(n5405) );
  MX4X1 U6176 ( .A(\ram[72][8] ), .B(\ram[73][8] ), .C(\ram[74][8] ), .D(
        \ram[75][8] ), .S0(n6314), .S1(n6180), .Y(n5403) );
  MX4X1 U6177 ( .A(\ram[68][8] ), .B(\ram[69][8] ), .C(\ram[70][8] ), .D(
        \ram[71][8] ), .S0(n6314), .S1(n6180), .Y(n5404) );
  MX4X1 U6178 ( .A(n5384), .B(n5382), .C(n5383), .D(n5381), .S0(n6037), .S1(
        n6065), .Y(n5385) );
  MX4X1 U6179 ( .A(\ram[128][8] ), .B(\ram[129][8] ), .C(\ram[130][8] ), .D(
        \ram[131][8] ), .S0(n6312), .S1(n6178), .Y(n5384) );
  MX4X1 U6180 ( .A(\ram[136][8] ), .B(\ram[137][8] ), .C(\ram[138][8] ), .D(
        \ram[139][8] ), .S0(n6312), .S1(n6178), .Y(n5382) );
  MX4X1 U6181 ( .A(\ram[132][8] ), .B(\ram[133][8] ), .C(\ram[134][8] ), .D(
        \ram[135][8] ), .S0(n6312), .S1(n6178), .Y(n5383) );
  MX4X1 U6182 ( .A(n5426), .B(n5424), .C(n5425), .D(n5423), .S0(n6038), .S1(
        n6066), .Y(n5427) );
  MX4X1 U6183 ( .A(\ram[0][8] ), .B(\ram[1][8] ), .C(\ram[2][8] ), .D(
        \ram[3][8] ), .S0(n6315), .S1(n6181), .Y(n5426) );
  MX4X1 U6184 ( .A(\ram[8][8] ), .B(\ram[9][8] ), .C(\ram[10][8] ), .D(
        \ram[11][8] ), .S0(n6315), .S1(n6181), .Y(n5424) );
  MX4X1 U6185 ( .A(\ram[4][8] ), .B(\ram[5][8] ), .C(\ram[6][8] ), .D(
        \ram[7][8] ), .S0(n6315), .S1(n6181), .Y(n5425) );
  MX4X1 U6186 ( .A(n5489), .B(n5487), .C(n5488), .D(n5486), .S0(n6039), .S1(
        n6067), .Y(n5490) );
  MX4X1 U6187 ( .A(\ram[64][9] ), .B(\ram[65][9] ), .C(\ram[66][9] ), .D(
        \ram[67][9] ), .S0(n6319), .S1(n6185), .Y(n5489) );
  MX4X1 U6188 ( .A(\ram[72][9] ), .B(\ram[73][9] ), .C(\ram[74][9] ), .D(
        \ram[75][9] ), .S0(n6319), .S1(n6185), .Y(n5487) );
  MX4X1 U6189 ( .A(\ram[68][9] ), .B(\ram[69][9] ), .C(\ram[70][9] ), .D(
        \ram[71][9] ), .S0(n6319), .S1(n6185), .Y(n5488) );
  MX4X1 U6190 ( .A(n5468), .B(n5466), .C(n5467), .D(n5465), .S0(n6039), .S1(
        n6067), .Y(n5469) );
  MX4X1 U6191 ( .A(\ram[128][9] ), .B(\ram[129][9] ), .C(\ram[130][9] ), .D(
        \ram[131][9] ), .S0(n6318), .S1(n6184), .Y(n5468) );
  MX4X1 U6192 ( .A(\ram[136][9] ), .B(\ram[137][9] ), .C(\ram[138][9] ), .D(
        \ram[139][9] ), .S0(n6318), .S1(n6184), .Y(n5466) );
  MX4X1 U6193 ( .A(\ram[132][9] ), .B(\ram[133][9] ), .C(\ram[134][9] ), .D(
        \ram[135][9] ), .S0(n6318), .S1(n6184), .Y(n5467) );
  MX4X1 U6194 ( .A(n5510), .B(n5508), .C(n5509), .D(n5507), .S0(n6039), .S1(
        n6067), .Y(n5511) );
  MX4X1 U6195 ( .A(\ram[0][9] ), .B(\ram[1][9] ), .C(\ram[2][9] ), .D(
        \ram[3][9] ), .S0(n6320), .S1(n6186), .Y(n5510) );
  MX4X1 U6196 ( .A(\ram[8][9] ), .B(\ram[9][9] ), .C(\ram[10][9] ), .D(
        \ram[11][9] ), .S0(n6320), .S1(n6186), .Y(n5508) );
  MX4X1 U6197 ( .A(\ram[4][9] ), .B(\ram[5][9] ), .C(\ram[6][9] ), .D(
        \ram[7][9] ), .S0(n6320), .S1(n6186), .Y(n5509) );
  MX4X1 U6198 ( .A(n5552), .B(n5550), .C(n5551), .D(n5549), .S0(n6040), .S1(
        n6068), .Y(n5553) );
  MX4X1 U6199 ( .A(\ram[128][10] ), .B(\ram[129][10] ), .C(\ram[130][10] ), 
        .D(\ram[131][10] ), .S0(n6323), .S1(n6189), .Y(n5552) );
  MX4X1 U6200 ( .A(\ram[136][10] ), .B(\ram[137][10] ), .C(\ram[138][10] ), 
        .D(\ram[139][10] ), .S0(n6323), .S1(n6189), .Y(n5550) );
  MX4X1 U6201 ( .A(\ram[132][10] ), .B(\ram[133][10] ), .C(\ram[134][10] ), 
        .D(\ram[135][10] ), .S0(n6323), .S1(n6189), .Y(n5551) );
  MX4X1 U6202 ( .A(n5573), .B(n5571), .C(n5572), .D(n5570), .S0(n6040), .S1(
        n6068), .Y(n5574) );
  MX4X1 U6203 ( .A(\ram[64][10] ), .B(\ram[65][10] ), .C(\ram[66][10] ), .D(
        \ram[67][10] ), .S0(n6324), .S1(n6190), .Y(n5573) );
  MX4X1 U6204 ( .A(\ram[72][10] ), .B(\ram[73][10] ), .C(\ram[74][10] ), .D(
        \ram[75][10] ), .S0(n6324), .S1(n6190), .Y(n5571) );
  MX4X1 U6205 ( .A(\ram[68][10] ), .B(\ram[69][10] ), .C(\ram[70][10] ), .D(
        \ram[71][10] ), .S0(n6324), .S1(n6190), .Y(n5572) );
  MX4X1 U6206 ( .A(n5594), .B(n5592), .C(n5593), .D(n5591), .S0(n6041), .S1(
        n6069), .Y(n5595) );
  MX4X1 U6207 ( .A(\ram[0][10] ), .B(\ram[1][10] ), .C(\ram[2][10] ), .D(
        \ram[3][10] ), .S0(n6326), .S1(n6192), .Y(n5594) );
  MX4X1 U6208 ( .A(\ram[8][10] ), .B(\ram[9][10] ), .C(\ram[10][10] ), .D(
        \ram[11][10] ), .S0(n6326), .S1(n6192), .Y(n5592) );
  MX4X1 U6209 ( .A(\ram[4][10] ), .B(\ram[5][10] ), .C(\ram[6][10] ), .D(
        \ram[7][10] ), .S0(n6326), .S1(n6192), .Y(n5593) );
  MX4X1 U6210 ( .A(n5657), .B(n5655), .C(n5656), .D(n5654), .S0(n6042), .S1(
        n6070), .Y(n5658) );
  MX4X1 U6211 ( .A(\ram[64][11] ), .B(\ram[65][11] ), .C(\ram[66][11] ), .D(
        \ram[67][11] ), .S0(n6330), .S1(n6196), .Y(n5657) );
  MX4X1 U6212 ( .A(\ram[72][11] ), .B(\ram[73][11] ), .C(\ram[74][11] ), .D(
        \ram[75][11] ), .S0(n6330), .S1(n6196), .Y(n5655) );
  MX4X1 U6213 ( .A(\ram[68][11] ), .B(\ram[69][11] ), .C(\ram[70][11] ), .D(
        \ram[71][11] ), .S0(n6330), .S1(n6196), .Y(n5656) );
  MX4X1 U6214 ( .A(n5636), .B(n5634), .C(n5635), .D(n5633), .S0(n6041), .S1(
        n6069), .Y(n5637) );
  MX4X1 U6215 ( .A(\ram[128][11] ), .B(\ram[129][11] ), .C(\ram[130][11] ), 
        .D(\ram[131][11] ), .S0(n6328), .S1(n6194), .Y(n5636) );
  MX4X1 U6216 ( .A(\ram[136][11] ), .B(\ram[137][11] ), .C(\ram[138][11] ), 
        .D(\ram[139][11] ), .S0(n6328), .S1(n6194), .Y(n5634) );
  MX4X1 U6217 ( .A(\ram[132][11] ), .B(\ram[133][11] ), .C(\ram[134][11] ), 
        .D(\ram[135][11] ), .S0(n6328), .S1(n6194), .Y(n5635) );
  MX4X1 U6218 ( .A(n5678), .B(n5676), .C(n5677), .D(n5675), .S0(n6042), .S1(
        n6070), .Y(n5679) );
  MX4X1 U6219 ( .A(\ram[0][11] ), .B(\ram[1][11] ), .C(\ram[2][11] ), .D(
        \ram[3][11] ), .S0(n6331), .S1(n6197), .Y(n5678) );
  MX4X1 U6220 ( .A(\ram[8][11] ), .B(\ram[9][11] ), .C(\ram[10][11] ), .D(
        \ram[11][11] ), .S0(n6331), .S1(n6197), .Y(n5676) );
  MX4X1 U6221 ( .A(\ram[4][11] ), .B(\ram[5][11] ), .C(\ram[6][11] ), .D(
        \ram[7][11] ), .S0(n6331), .S1(n6197), .Y(n5677) );
  MX4X1 U6222 ( .A(n5741), .B(n5739), .C(n5740), .D(n5738), .S0(n6043), .S1(
        n6071), .Y(n5742) );
  MX4X1 U6223 ( .A(\ram[64][12] ), .B(\ram[65][12] ), .C(\ram[66][12] ), .D(
        \ram[67][12] ), .S0(n6335), .S1(n6201), .Y(n5741) );
  MX4X1 U6224 ( .A(\ram[72][12] ), .B(\ram[73][12] ), .C(\ram[74][12] ), .D(
        \ram[75][12] ), .S0(n6335), .S1(n6201), .Y(n5739) );
  MX4X1 U6225 ( .A(\ram[68][12] ), .B(\ram[69][12] ), .C(\ram[70][12] ), .D(
        \ram[71][12] ), .S0(n6335), .S1(n6201), .Y(n5740) );
  MX4X1 U6226 ( .A(n5720), .B(n5718), .C(n5719), .D(n5717), .S0(n6043), .S1(
        n6071), .Y(n5721) );
  MX4X1 U6227 ( .A(\ram[128][12] ), .B(\ram[129][12] ), .C(\ram[130][12] ), 
        .D(\ram[131][12] ), .S0(n6334), .S1(n6200), .Y(n5720) );
  MX4X1 U6228 ( .A(\ram[136][12] ), .B(\ram[137][12] ), .C(\ram[138][12] ), 
        .D(\ram[139][12] ), .S0(n6334), .S1(n6200), .Y(n5718) );
  MX4X1 U6229 ( .A(\ram[132][12] ), .B(\ram[133][12] ), .C(\ram[134][12] ), 
        .D(\ram[135][12] ), .S0(n6334), .S1(n6200), .Y(n5719) );
  MX4X1 U6230 ( .A(n5762), .B(n5760), .C(n5761), .D(n5759), .S0(n6043), .S1(
        n6071), .Y(n5763) );
  MX4X1 U6231 ( .A(\ram[0][12] ), .B(\ram[1][12] ), .C(\ram[2][12] ), .D(
        \ram[3][12] ), .S0(n6336), .S1(n6202), .Y(n5762) );
  MX4X1 U6232 ( .A(\ram[8][12] ), .B(\ram[9][12] ), .C(\ram[10][12] ), .D(
        \ram[11][12] ), .S0(n6336), .S1(n6202), .Y(n5760) );
  MX4X1 U6233 ( .A(\ram[4][12] ), .B(\ram[5][12] ), .C(\ram[6][12] ), .D(
        \ram[7][12] ), .S0(n6336), .S1(n6202), .Y(n5761) );
  MX4X1 U6234 ( .A(n5825), .B(n5823), .C(n5824), .D(n5822), .S0(n6044), .S1(
        n6072), .Y(n5826) );
  MX4X1 U6235 ( .A(\ram[64][13] ), .B(\ram[65][13] ), .C(\ram[66][13] ), .D(
        \ram[67][13] ), .S0(n6340), .S1(n6206), .Y(n5825) );
  MX4X1 U6236 ( .A(\ram[72][13] ), .B(\ram[73][13] ), .C(\ram[74][13] ), .D(
        \ram[75][13] ), .S0(n6340), .S1(n6206), .Y(n5823) );
  MX4X1 U6237 ( .A(\ram[68][13] ), .B(\ram[69][13] ), .C(\ram[70][13] ), .D(
        \ram[71][13] ), .S0(n6340), .S1(n6206), .Y(n5824) );
  MX4X1 U6238 ( .A(n5804), .B(n5802), .C(n5803), .D(n5801), .S0(n6044), .S1(
        n6072), .Y(n5805) );
  MX4X1 U6239 ( .A(\ram[128][13] ), .B(\ram[129][13] ), .C(\ram[130][13] ), 
        .D(\ram[131][13] ), .S0(n6339), .S1(n6205), .Y(n5804) );
  MX4X1 U6240 ( .A(\ram[136][13] ), .B(\ram[137][13] ), .C(\ram[138][13] ), 
        .D(\ram[139][13] ), .S0(n6339), .S1(n6205), .Y(n5802) );
  MX4X1 U6241 ( .A(\ram[132][13] ), .B(\ram[133][13] ), .C(\ram[134][13] ), 
        .D(\ram[135][13] ), .S0(n6339), .S1(n6205), .Y(n5803) );
  MX4X1 U6242 ( .A(n5846), .B(n5844), .C(n5845), .D(n5843), .S0(n6045), .S1(
        n6073), .Y(n5847) );
  MX4X1 U6243 ( .A(\ram[0][13] ), .B(\ram[1][13] ), .C(\ram[2][13] ), .D(
        \ram[3][13] ), .S0(n6342), .S1(n6208), .Y(n5846) );
  MX4X1 U6244 ( .A(\ram[8][13] ), .B(\ram[9][13] ), .C(\ram[10][13] ), .D(
        \ram[11][13] ), .S0(n6342), .S1(n6208), .Y(n5844) );
  MX4X1 U6245 ( .A(\ram[4][13] ), .B(\ram[5][13] ), .C(\ram[6][13] ), .D(
        \ram[7][13] ), .S0(n6342), .S1(n6208), .Y(n5845) );
  MX4X1 U6246 ( .A(n5909), .B(n5907), .C(n5908), .D(n5906), .S0(n6046), .S1(
        n6060), .Y(n5910) );
  MX4X1 U6247 ( .A(\ram[64][14] ), .B(\ram[65][14] ), .C(\ram[66][14] ), .D(
        \ram[67][14] ), .S0(n6346), .S1(n6212), .Y(n5909) );
  MX4X1 U6248 ( .A(\ram[72][14] ), .B(\ram[73][14] ), .C(\ram[74][14] ), .D(
        \ram[75][14] ), .S0(n6346), .S1(n6212), .Y(n5907) );
  MX4X1 U6249 ( .A(\ram[68][14] ), .B(\ram[69][14] ), .C(\ram[70][14] ), .D(
        \ram[71][14] ), .S0(n6346), .S1(n6212), .Y(n5908) );
  MX4X1 U6250 ( .A(n5888), .B(n5886), .C(n5887), .D(n5885), .S0(n6045), .S1(
        n6073), .Y(n5889) );
  MX4X1 U6251 ( .A(\ram[128][14] ), .B(\ram[129][14] ), .C(\ram[130][14] ), 
        .D(\ram[131][14] ), .S0(n6344), .S1(n6210), .Y(n5888) );
  MX4X1 U6252 ( .A(\ram[136][14] ), .B(\ram[137][14] ), .C(\ram[138][14] ), 
        .D(\ram[139][14] ), .S0(n6344), .S1(n6210), .Y(n5886) );
  MX4X1 U6253 ( .A(\ram[132][14] ), .B(\ram[133][14] ), .C(\ram[134][14] ), 
        .D(\ram[135][14] ), .S0(n6344), .S1(n6210), .Y(n5887) );
  MX4X1 U6254 ( .A(n5930), .B(n5928), .C(n5929), .D(n5927), .S0(n6046), .S1(
        n6073), .Y(n5931) );
  MX4X1 U6255 ( .A(\ram[0][14] ), .B(\ram[1][14] ), .C(\ram[2][14] ), .D(
        \ram[3][14] ), .S0(n6347), .S1(n6140), .Y(n5930) );
  MX4X1 U6256 ( .A(\ram[8][14] ), .B(\ram[9][14] ), .C(\ram[10][14] ), .D(
        \ram[11][14] ), .S0(n6347), .S1(n6214), .Y(n5928) );
  MX4X1 U6257 ( .A(\ram[4][14] ), .B(\ram[5][14] ), .C(\ram[6][14] ), .D(
        \ram[7][14] ), .S0(n6347), .S1(n6140), .Y(n5929) );
  MX4X1 U6258 ( .A(n5993), .B(n5991), .C(n5992), .D(n5990), .S0(n6047), .S1(
        n6061), .Y(n5994) );
  MX4X1 U6259 ( .A(\ram[64][15] ), .B(\ram[65][15] ), .C(\ram[66][15] ), .D(
        \ram[67][15] ), .S0(n6351), .S1(n6165), .Y(n5993) );
  MX4X1 U6260 ( .A(\ram[72][15] ), .B(\ram[73][15] ), .C(\ram[74][15] ), .D(
        \ram[75][15] ), .S0(n6351), .S1(n6076), .Y(n5991) );
  MX4X1 U6261 ( .A(\ram[68][15] ), .B(\ram[69][15] ), .C(\ram[70][15] ), .D(
        \ram[71][15] ), .S0(n6351), .S1(n6190), .Y(n5992) );
  MX4X1 U6262 ( .A(n5972), .B(n5970), .C(n5971), .D(n5969), .S0(n6047), .S1(
        n6061), .Y(n5973) );
  MX4X1 U6263 ( .A(\ram[128][15] ), .B(\ram[129][15] ), .C(\ram[130][15] ), 
        .D(\ram[131][15] ), .S0(n6350), .S1(n6192), .Y(n5972) );
  MX4X1 U6264 ( .A(\ram[136][15] ), .B(\ram[137][15] ), .C(\ram[138][15] ), 
        .D(\ram[139][15] ), .S0(n6350), .S1(n6140), .Y(n5970) );
  MX4X1 U6265 ( .A(\ram[132][15] ), .B(\ram[133][15] ), .C(\ram[134][15] ), 
        .D(\ram[135][15] ), .S0(n6350), .S1(n6139), .Y(n5971) );
  MX4X1 U6266 ( .A(n6014), .B(n6012), .C(n6013), .D(n6011), .S0(n6047), .S1(
        n6073), .Y(n6015) );
  MX4X1 U6267 ( .A(\ram[0][15] ), .B(\ram[1][15] ), .C(\ram[2][15] ), .D(
        \ram[3][15] ), .S0(n6352), .S1(n6213), .Y(n6014) );
  MX4X1 U6268 ( .A(\ram[8][15] ), .B(\ram[9][15] ), .C(\ram[10][15] ), .D(
        \ram[11][15] ), .S0(n6352), .S1(n6140), .Y(n6012) );
  MX4X1 U6269 ( .A(\ram[4][15] ), .B(\ram[5][15] ), .C(\ram[6][15] ), .D(
        \ram[7][15] ), .S0(n6352), .S1(n6160), .Y(n6013) );
  MX4X1 U6270 ( .A(\ram[124][0] ), .B(\ram[125][0] ), .C(\ram[126][0] ), .D(
        \ram[127][0] ), .S0(n6270), .S1(n6136), .Y(n4715) );
  MX4X1 U6271 ( .A(\ram[92][0] ), .B(\ram[93][0] ), .C(\ram[94][0] ), .D(
        \ram[95][0] ), .S0(n6271), .S1(n6137), .Y(n4725) );
  MX4X1 U6272 ( .A(\ram[108][0] ), .B(\ram[109][0] ), .C(\ram[110][0] ), .D(
        \ram[111][0] ), .S0(n6270), .S1(n6136), .Y(n4720) );
  MX4X1 U6273 ( .A(\ram[76][0] ), .B(\ram[77][0] ), .C(\ram[78][0] ), .D(
        \ram[79][0] ), .S0(n6271), .S1(n6137), .Y(n4730) );
  MX4X1 U6274 ( .A(\ram[188][0] ), .B(\ram[189][0] ), .C(\ram[190][0] ), .D(
        \ram[191][0] ), .S0(n6269), .S1(n6135), .Y(n4694) );
  MX4X1 U6275 ( .A(\ram[156][0] ), .B(\ram[157][0] ), .C(\ram[158][0] ), .D(
        \ram[159][0] ), .S0(n6269), .S1(n6135), .Y(n4704) );
  MX4X1 U6276 ( .A(\ram[172][0] ), .B(\ram[173][0] ), .C(\ram[174][0] ), .D(
        \ram[175][0] ), .S0(n6269), .S1(n6135), .Y(n4699) );
  MX4X1 U6277 ( .A(\ram[140][0] ), .B(\ram[141][0] ), .C(\ram[142][0] ), .D(
        \ram[143][0] ), .S0(n6270), .S1(n6136), .Y(n4709) );
  MX4X1 U6278 ( .A(\ram[60][0] ), .B(\ram[61][0] ), .C(\ram[62][0] ), .D(
        \ram[63][0] ), .S0(n6271), .S1(n6137), .Y(n4736) );
  MX4X1 U6279 ( .A(\ram[28][0] ), .B(\ram[29][0] ), .C(\ram[30][0] ), .D(
        \ram[31][0] ), .S0(n6272), .S1(n6138), .Y(n4746) );
  MX4X1 U6280 ( .A(\ram[44][0] ), .B(\ram[45][0] ), .C(\ram[46][0] ), .D(
        \ram[47][0] ), .S0(n6272), .S1(n6138), .Y(n4741) );
  MX4X1 U6281 ( .A(\ram[12][0] ), .B(\ram[13][0] ), .C(\ram[14][0] ), .D(
        \ram[15][0] ), .S0(n6272), .S1(n6138), .Y(n4751) );
  MX4X1 U6282 ( .A(\ram[220][0] ), .B(\ram[221][0] ), .C(\ram[222][0] ), .D(
        \ram[223][0] ), .S0(n6268), .S1(n6134), .Y(n4683) );
  MX4X1 U6283 ( .A(\ram[236][0] ), .B(\ram[237][0] ), .C(\ram[238][0] ), .D(
        \ram[239][0] ), .S0(n6268), .S1(n6134), .Y(n4678) );
  MX4X1 U6284 ( .A(\ram[204][0] ), .B(\ram[205][0] ), .C(\ram[206][0] ), .D(
        \ram[207][0] ), .S0(n6268), .S1(n6134), .Y(n4688) );
  MX4X1 U6285 ( .A(\ram[252][1] ), .B(\ram[253][1] ), .C(\ram[254][1] ), .D(
        \ram[255][1] ), .S0(n6273), .S1(n6139), .Y(n4757) );
  MX4X1 U6286 ( .A(\ram[220][1] ), .B(\ram[221][1] ), .C(\ram[222][1] ), .D(
        \ram[223][1] ), .S0(n6273), .S1(n6139), .Y(n4767) );
  MX4X1 U6287 ( .A(\ram[236][1] ), .B(\ram[237][1] ), .C(\ram[238][1] ), .D(
        \ram[239][1] ), .S0(n6273), .S1(n6139), .Y(n4762) );
  MX4X1 U6288 ( .A(\ram[204][1] ), .B(\ram[205][1] ), .C(\ram[206][1] ), .D(
        \ram[207][1] ), .S0(n6274), .S1(n6140), .Y(n4772) );
  MX4X1 U6289 ( .A(\ram[124][1] ), .B(\ram[125][1] ), .C(\ram[126][1] ), .D(
        \ram[127][1] ), .S0(n6275), .S1(n6141), .Y(n4799) );
  MX4X1 U6290 ( .A(\ram[92][1] ), .B(\ram[93][1] ), .C(\ram[94][1] ), .D(
        \ram[95][1] ), .S0(n6276), .S1(n6142), .Y(n4809) );
  MX4X1 U6291 ( .A(\ram[108][1] ), .B(\ram[109][1] ), .C(\ram[110][1] ), .D(
        \ram[111][1] ), .S0(n6276), .S1(n6142), .Y(n4804) );
  MX4X1 U6292 ( .A(\ram[76][1] ), .B(\ram[77][1] ), .C(\ram[78][1] ), .D(
        \ram[79][1] ), .S0(n6276), .S1(n6142), .Y(n4814) );
  MX4X1 U6293 ( .A(\ram[188][1] ), .B(\ram[189][1] ), .C(\ram[190][1] ), .D(
        \ram[191][1] ), .S0(n6274), .S1(n6140), .Y(n4778) );
  MX4X1 U6294 ( .A(\ram[156][1] ), .B(\ram[157][1] ), .C(\ram[158][1] ), .D(
        \ram[159][1] ), .S0(n6275), .S1(n6141), .Y(n4788) );
  MX4X1 U6295 ( .A(\ram[172][1] ), .B(\ram[173][1] ), .C(\ram[174][1] ), .D(
        \ram[175][1] ), .S0(n6274), .S1(n6140), .Y(n4783) );
  MX4X1 U6296 ( .A(\ram[140][1] ), .B(\ram[141][1] ), .C(\ram[142][1] ), .D(
        \ram[143][1] ), .S0(n6275), .S1(n6141), .Y(n4793) );
  MX4X1 U6297 ( .A(\ram[60][1] ), .B(\ram[61][1] ), .C(\ram[62][1] ), .D(
        \ram[63][1] ), .S0(n6277), .S1(n6143), .Y(n4820) );
  MX4X1 U6298 ( .A(\ram[28][1] ), .B(\ram[29][1] ), .C(\ram[30][1] ), .D(
        \ram[31][1] ), .S0(n6277), .S1(n6143), .Y(n4830) );
  MX4X1 U6299 ( .A(\ram[44][1] ), .B(\ram[45][1] ), .C(\ram[46][1] ), .D(
        \ram[47][1] ), .S0(n6277), .S1(n6143), .Y(n4825) );
  MX4X1 U6300 ( .A(\ram[12][1] ), .B(\ram[13][1] ), .C(\ram[14][1] ), .D(
        \ram[15][1] ), .S0(n6278), .S1(n6144), .Y(n4835) );
  MX4X1 U6301 ( .A(\ram[252][2] ), .B(\ram[253][2] ), .C(\ram[254][2] ), .D(
        \ram[255][2] ), .S0(n6278), .S1(n6144), .Y(n4841) );
  MX4X1 U6302 ( .A(\ram[220][2] ), .B(\ram[221][2] ), .C(\ram[222][2] ), .D(
        \ram[223][2] ), .S0(n6279), .S1(n6145), .Y(n4851) );
  MX4X1 U6303 ( .A(\ram[236][2] ), .B(\ram[237][2] ), .C(\ram[238][2] ), .D(
        \ram[239][2] ), .S0(n6278), .S1(n6144), .Y(n4846) );
  MX4X1 U6304 ( .A(\ram[204][2] ), .B(\ram[205][2] ), .C(\ram[206][2] ), .D(
        \ram[207][2] ), .S0(n6279), .S1(n6145), .Y(n4856) );
  MX4X1 U6305 ( .A(\ram[124][2] ), .B(\ram[125][2] ), .C(\ram[126][2] ), .D(
        \ram[127][2] ), .S0(n6281), .S1(n6147), .Y(n4883) );
  MX4X1 U6306 ( .A(\ram[92][2] ), .B(\ram[93][2] ), .C(\ram[94][2] ), .D(
        \ram[95][2] ), .S0(n6281), .S1(n6147), .Y(n4893) );
  MX4X1 U6307 ( .A(\ram[108][2] ), .B(\ram[109][2] ), .C(\ram[110][2] ), .D(
        \ram[111][2] ), .S0(n6281), .S1(n6147), .Y(n4888) );
  MX4X1 U6308 ( .A(\ram[76][2] ), .B(\ram[77][2] ), .C(\ram[78][2] ), .D(
        \ram[79][2] ), .S0(n6282), .S1(n6148), .Y(n4898) );
  MX4X1 U6309 ( .A(\ram[188][2] ), .B(\ram[189][2] ), .C(\ram[190][2] ), .D(
        \ram[191][2] ), .S0(n6279), .S1(n6145), .Y(n4862) );
  MX4X1 U6310 ( .A(\ram[156][2] ), .B(\ram[157][2] ), .C(\ram[158][2] ), .D(
        \ram[159][2] ), .S0(n6280), .S1(n6146), .Y(n4872) );
  MX4X1 U6311 ( .A(\ram[172][2] ), .B(\ram[173][2] ), .C(\ram[174][2] ), .D(
        \ram[175][2] ), .S0(n6280), .S1(n6146), .Y(n4867) );
  MX4X1 U6312 ( .A(\ram[140][2] ), .B(\ram[141][2] ), .C(\ram[142][2] ), .D(
        \ram[143][2] ), .S0(n6280), .S1(n6146), .Y(n4877) );
  MX4X1 U6313 ( .A(\ram[60][2] ), .B(\ram[61][2] ), .C(\ram[62][2] ), .D(
        \ram[63][2] ), .S0(n6282), .S1(n6148), .Y(n4904) );
  MX4X1 U6314 ( .A(\ram[28][2] ), .B(\ram[29][2] ), .C(\ram[30][2] ), .D(
        \ram[31][2] ), .S0(n6283), .S1(n6149), .Y(n4914) );
  MX4X1 U6315 ( .A(\ram[44][2] ), .B(\ram[45][2] ), .C(\ram[46][2] ), .D(
        \ram[47][2] ), .S0(n6282), .S1(n6148), .Y(n4909) );
  MX4X1 U6316 ( .A(\ram[12][2] ), .B(\ram[13][2] ), .C(\ram[14][2] ), .D(
        \ram[15][2] ), .S0(n6283), .S1(n6149), .Y(n4919) );
  MX4X1 U6317 ( .A(\ram[92][3] ), .B(\ram[93][3] ), .C(\ram[94][3] ), .D(
        \ram[95][3] ), .S0(n6287), .S1(n6153), .Y(n4977) );
  MX4X1 U6318 ( .A(\ram[124][3] ), .B(\ram[125][3] ), .C(\ram[126][3] ), .D(
        \ram[127][3] ), .S0(n6286), .S1(n6152), .Y(n4967) );
  MX4X1 U6319 ( .A(\ram[76][3] ), .B(\ram[77][3] ), .C(\ram[78][3] ), .D(
        \ram[79][3] ), .S0(n6287), .S1(n6153), .Y(n4982) );
  MX4X1 U6320 ( .A(\ram[108][3] ), .B(\ram[109][3] ), .C(\ram[110][3] ), .D(
        \ram[111][3] ), .S0(n6286), .S1(n6152), .Y(n4972) );
  MX4X1 U6321 ( .A(\ram[252][3] ), .B(\ram[253][3] ), .C(\ram[254][3] ), .D(
        \ram[255][3] ), .S0(n6283), .S1(n6149), .Y(n4925) );
  MX4X1 U6322 ( .A(\ram[220][3] ), .B(\ram[221][3] ), .C(\ram[222][3] ), .D(
        \ram[223][3] ), .S0(n6284), .S1(n6150), .Y(n4935) );
  MX4X1 U6323 ( .A(\ram[236][3] ), .B(\ram[237][3] ), .C(\ram[238][3] ), .D(
        \ram[239][3] ), .S0(n6284), .S1(n6150), .Y(n4930) );
  MX4X1 U6324 ( .A(\ram[204][3] ), .B(\ram[205][3] ), .C(\ram[206][3] ), .D(
        \ram[207][3] ), .S0(n6284), .S1(n6150), .Y(n4940) );
  MX4X1 U6325 ( .A(\ram[60][3] ), .B(\ram[61][3] ), .C(\ram[62][3] ), .D(
        \ram[63][3] ), .S0(n6287), .S1(n6153), .Y(n4988) );
  MX4X1 U6326 ( .A(\ram[28][3] ), .B(\ram[29][3] ), .C(\ram[30][3] ), .D(
        \ram[31][3] ), .S0(n6288), .S1(n6154), .Y(n4998) );
  MX4X1 U6327 ( .A(\ram[44][3] ), .B(\ram[45][3] ), .C(\ram[46][3] ), .D(
        \ram[47][3] ), .S0(n6288), .S1(n6154), .Y(n4993) );
  MX4X1 U6328 ( .A(\ram[12][3] ), .B(\ram[13][3] ), .C(\ram[14][3] ), .D(
        \ram[15][3] ), .S0(n6288), .S1(n6154), .Y(n5003) );
  MX4X1 U6329 ( .A(\ram[188][3] ), .B(\ram[189][3] ), .C(\ram[190][3] ), .D(
        \ram[191][3] ), .S0(n6285), .S1(n6151), .Y(n4946) );
  MX4X1 U6330 ( .A(\ram[156][3] ), .B(\ram[157][3] ), .C(\ram[158][3] ), .D(
        \ram[159][3] ), .S0(n6285), .S1(n6151), .Y(n4956) );
  MX4X1 U6331 ( .A(\ram[172][3] ), .B(\ram[173][3] ), .C(\ram[174][3] ), .D(
        \ram[175][3] ), .S0(n6285), .S1(n6151), .Y(n4951) );
  MX4X1 U6332 ( .A(\ram[140][3] ), .B(\ram[141][3] ), .C(\ram[142][3] ), .D(
        \ram[143][3] ), .S0(n6286), .S1(n6152), .Y(n4961) );
  MX4X1 U6333 ( .A(\ram[252][4] ), .B(\ram[253][4] ), .C(\ram[254][4] ), .D(
        \ram[255][4] ), .S0(n6289), .S1(n6155), .Y(n5009) );
  MX4X1 U6334 ( .A(\ram[220][4] ), .B(\ram[221][4] ), .C(\ram[222][4] ), .D(
        \ram[223][4] ), .S0(n6289), .S1(n6155), .Y(n5019) );
  MX4X1 U6335 ( .A(\ram[236][4] ), .B(\ram[237][4] ), .C(\ram[238][4] ), .D(
        \ram[239][4] ), .S0(n6289), .S1(n6155), .Y(n5014) );
  MX4X1 U6336 ( .A(\ram[204][4] ), .B(\ram[205][4] ), .C(\ram[206][4] ), .D(
        \ram[207][4] ), .S0(n6290), .S1(n6156), .Y(n5024) );
  MX4X1 U6337 ( .A(\ram[124][4] ), .B(\ram[125][4] ), .C(\ram[126][4] ), .D(
        \ram[127][4] ), .S0(n6291), .S1(n6157), .Y(n5051) );
  MX4X1 U6338 ( .A(\ram[92][4] ), .B(\ram[93][4] ), .C(\ram[94][4] ), .D(
        \ram[95][4] ), .S0(n6292), .S1(n6158), .Y(n5061) );
  MX4X1 U6339 ( .A(\ram[108][4] ), .B(\ram[109][4] ), .C(\ram[110][4] ), .D(
        \ram[111][4] ), .S0(n6292), .S1(n6158), .Y(n5056) );
  MX4X1 U6340 ( .A(\ram[76][4] ), .B(\ram[77][4] ), .C(\ram[78][4] ), .D(
        \ram[79][4] ), .S0(n6292), .S1(n6158), .Y(n5066) );
  MX4X1 U6341 ( .A(\ram[188][4] ), .B(\ram[189][4] ), .C(\ram[190][4] ), .D(
        \ram[191][4] ), .S0(n6290), .S1(n6156), .Y(n5030) );
  MX4X1 U6342 ( .A(\ram[156][4] ), .B(\ram[157][4] ), .C(\ram[158][4] ), .D(
        \ram[159][4] ), .S0(n6291), .S1(n6157), .Y(n5040) );
  MX4X1 U6343 ( .A(\ram[172][4] ), .B(\ram[173][4] ), .C(\ram[174][4] ), .D(
        \ram[175][4] ), .S0(n6290), .S1(n6156), .Y(n5035) );
  MX4X1 U6344 ( .A(\ram[140][4] ), .B(\ram[141][4] ), .C(\ram[142][4] ), .D(
        \ram[143][4] ), .S0(n6291), .S1(n6157), .Y(n5045) );
  MX4X1 U6345 ( .A(\ram[60][4] ), .B(\ram[61][4] ), .C(\ram[62][4] ), .D(
        \ram[63][4] ), .S0(n6293), .S1(n6159), .Y(n5072) );
  MX4X1 U6346 ( .A(\ram[28][4] ), .B(\ram[29][4] ), .C(\ram[30][4] ), .D(
        \ram[31][4] ), .S0(n6293), .S1(n6159), .Y(n5082) );
  MX4X1 U6347 ( .A(\ram[44][4] ), .B(\ram[45][4] ), .C(\ram[46][4] ), .D(
        \ram[47][4] ), .S0(n6293), .S1(n6159), .Y(n5077) );
  MX4X1 U6348 ( .A(\ram[12][4] ), .B(\ram[13][4] ), .C(\ram[14][4] ), .D(
        \ram[15][4] ), .S0(n6294), .S1(n6160), .Y(n5087) );
  MX4X1 U6349 ( .A(\ram[252][5] ), .B(\ram[253][5] ), .C(\ram[254][5] ), .D(
        \ram[255][5] ), .S0(n6294), .S1(n6160), .Y(n5093) );
  MX4X1 U6350 ( .A(\ram[220][5] ), .B(\ram[221][5] ), .C(\ram[222][5] ), .D(
        \ram[223][5] ), .S0(n6295), .S1(n6161), .Y(n5103) );
  MX4X1 U6351 ( .A(\ram[236][5] ), .B(\ram[237][5] ), .C(\ram[238][5] ), .D(
        \ram[239][5] ), .S0(n6294), .S1(n6160), .Y(n5098) );
  MX4X1 U6352 ( .A(\ram[204][5] ), .B(\ram[205][5] ), .C(\ram[206][5] ), .D(
        \ram[207][5] ), .S0(n6295), .S1(n6161), .Y(n5108) );
  MX4X1 U6353 ( .A(\ram[124][5] ), .B(\ram[125][5] ), .C(\ram[126][5] ), .D(
        \ram[127][5] ), .S0(n6297), .S1(n6163), .Y(n5135) );
  MX4X1 U6354 ( .A(\ram[92][5] ), .B(\ram[93][5] ), .C(\ram[94][5] ), .D(
        \ram[95][5] ), .S0(n6297), .S1(n6163), .Y(n5145) );
  MX4X1 U6355 ( .A(\ram[108][5] ), .B(\ram[109][5] ), .C(\ram[110][5] ), .D(
        \ram[111][5] ), .S0(n6297), .S1(n6163), .Y(n5140) );
  MX4X1 U6356 ( .A(\ram[76][5] ), .B(\ram[77][5] ), .C(\ram[78][5] ), .D(
        \ram[79][5] ), .S0(n6298), .S1(n6164), .Y(n5150) );
  MX4X1 U6357 ( .A(\ram[188][5] ), .B(\ram[189][5] ), .C(\ram[190][5] ), .D(
        \ram[191][5] ), .S0(n6295), .S1(n6161), .Y(n5114) );
  MX4X1 U6358 ( .A(\ram[156][5] ), .B(\ram[157][5] ), .C(\ram[158][5] ), .D(
        \ram[159][5] ), .S0(n6296), .S1(n6162), .Y(n5124) );
  MX4X1 U6359 ( .A(\ram[172][5] ), .B(\ram[173][5] ), .C(\ram[174][5] ), .D(
        \ram[175][5] ), .S0(n6296), .S1(n6162), .Y(n5119) );
  MX4X1 U6360 ( .A(\ram[140][5] ), .B(\ram[141][5] ), .C(\ram[142][5] ), .D(
        \ram[143][5] ), .S0(n6296), .S1(n6162), .Y(n5129) );
  MX4X1 U6361 ( .A(\ram[60][5] ), .B(\ram[61][5] ), .C(\ram[62][5] ), .D(
        \ram[63][5] ), .S0(n6298), .S1(n6164), .Y(n5156) );
  MX4X1 U6362 ( .A(\ram[28][5] ), .B(\ram[29][5] ), .C(\ram[30][5] ), .D(
        \ram[31][5] ), .S0(n6299), .S1(n6165), .Y(n5166) );
  MX4X1 U6363 ( .A(\ram[44][5] ), .B(\ram[45][5] ), .C(\ram[46][5] ), .D(
        \ram[47][5] ), .S0(n6298), .S1(n6164), .Y(n5161) );
  MX4X1 U6364 ( .A(\ram[12][5] ), .B(\ram[13][5] ), .C(\ram[14][5] ), .D(
        \ram[15][5] ), .S0(n6299), .S1(n6165), .Y(n5171) );
  MX4X1 U6365 ( .A(\ram[252][6] ), .B(\ram[253][6] ), .C(\ram[254][6] ), .D(
        \ram[255][6] ), .S0(n6299), .S1(n6165), .Y(n5177) );
  MX4X1 U6366 ( .A(\ram[220][6] ), .B(\ram[221][6] ), .C(\ram[222][6] ), .D(
        \ram[223][6] ), .S0(n6300), .S1(n6166), .Y(n5187) );
  MX4X1 U6367 ( .A(\ram[236][6] ), .B(\ram[237][6] ), .C(\ram[238][6] ), .D(
        \ram[239][6] ), .S0(n6300), .S1(n6166), .Y(n5182) );
  MX4X1 U6368 ( .A(\ram[204][6] ), .B(\ram[205][6] ), .C(\ram[206][6] ), .D(
        \ram[207][6] ), .S0(n6300), .S1(n6166), .Y(n5192) );
  MX4X1 U6369 ( .A(\ram[124][6] ), .B(\ram[125][6] ), .C(\ram[126][6] ), .D(
        \ram[127][6] ), .S0(n6302), .S1(n6168), .Y(n5219) );
  MX4X1 U6370 ( .A(\ram[92][6] ), .B(\ram[93][6] ), .C(\ram[94][6] ), .D(
        \ram[95][6] ), .S0(n6303), .S1(n6169), .Y(n5229) );
  MX4X1 U6371 ( .A(\ram[108][6] ), .B(\ram[109][6] ), .C(\ram[110][6] ), .D(
        \ram[111][6] ), .S0(n6302), .S1(n6168), .Y(n5224) );
  MX4X1 U6372 ( .A(\ram[76][6] ), .B(\ram[77][6] ), .C(\ram[78][6] ), .D(
        \ram[79][6] ), .S0(n6303), .S1(n6169), .Y(n5234) );
  MX4X1 U6373 ( .A(\ram[188][6] ), .B(\ram[189][6] ), .C(\ram[190][6] ), .D(
        \ram[191][6] ), .S0(n6301), .S1(n6167), .Y(n5198) );
  MX4X1 U6374 ( .A(\ram[156][6] ), .B(\ram[157][6] ), .C(\ram[158][6] ), .D(
        \ram[159][6] ), .S0(n6301), .S1(n6167), .Y(n5208) );
  MX4X1 U6375 ( .A(\ram[172][6] ), .B(\ram[173][6] ), .C(\ram[174][6] ), .D(
        \ram[175][6] ), .S0(n6301), .S1(n6167), .Y(n5203) );
  MX4X1 U6376 ( .A(\ram[140][6] ), .B(\ram[141][6] ), .C(\ram[142][6] ), .D(
        \ram[143][6] ), .S0(n6302), .S1(n6168), .Y(n5213) );
  MX4X1 U6377 ( .A(\ram[60][6] ), .B(\ram[61][6] ), .C(\ram[62][6] ), .D(
        \ram[63][6] ), .S0(n6303), .S1(n6169), .Y(n5240) );
  MX4X1 U6378 ( .A(\ram[28][6] ), .B(\ram[29][6] ), .C(\ram[30][6] ), .D(
        \ram[31][6] ), .S0(n6304), .S1(n6170), .Y(n5250) );
  MX4X1 U6379 ( .A(\ram[44][6] ), .B(\ram[45][6] ), .C(\ram[46][6] ), .D(
        \ram[47][6] ), .S0(n6304), .S1(n6170), .Y(n5245) );
  MX4X1 U6380 ( .A(\ram[12][6] ), .B(\ram[13][6] ), .C(\ram[14][6] ), .D(
        \ram[15][6] ), .S0(n6304), .S1(n6170), .Y(n5255) );
  MX4X1 U6381 ( .A(\ram[252][7] ), .B(\ram[253][7] ), .C(\ram[254][7] ), .D(
        \ram[255][7] ), .S0(n6305), .S1(n6171), .Y(n5261) );
  MX4X1 U6382 ( .A(\ram[220][7] ), .B(\ram[221][7] ), .C(\ram[222][7] ), .D(
        \ram[223][7] ), .S0(n6305), .S1(n6171), .Y(n5271) );
  MX4X1 U6383 ( .A(\ram[236][7] ), .B(\ram[237][7] ), .C(\ram[238][7] ), .D(
        \ram[239][7] ), .S0(n6305), .S1(n6171), .Y(n5266) );
  MX4X1 U6384 ( .A(\ram[204][7] ), .B(\ram[205][7] ), .C(\ram[206][7] ), .D(
        \ram[207][7] ), .S0(n6306), .S1(n6172), .Y(n5276) );
  MX4X1 U6385 ( .A(\ram[124][7] ), .B(\ram[125][7] ), .C(\ram[126][7] ), .D(
        \ram[127][7] ), .S0(n6307), .S1(n6173), .Y(n5303) );
  MX4X1 U6386 ( .A(\ram[92][7] ), .B(\ram[93][7] ), .C(\ram[94][7] ), .D(
        \ram[95][7] ), .S0(n6308), .S1(n6174), .Y(n5313) );
  MX4X1 U6387 ( .A(\ram[108][7] ), .B(\ram[109][7] ), .C(\ram[110][7] ), .D(
        \ram[111][7] ), .S0(n6308), .S1(n6174), .Y(n5308) );
  MX4X1 U6388 ( .A(\ram[76][7] ), .B(\ram[77][7] ), .C(\ram[78][7] ), .D(
        \ram[79][7] ), .S0(n6308), .S1(n6174), .Y(n5318) );
  MX4X1 U6389 ( .A(\ram[188][7] ), .B(\ram[189][7] ), .C(\ram[190][7] ), .D(
        \ram[191][7] ), .S0(n6306), .S1(n6172), .Y(n5282) );
  MX4X1 U6390 ( .A(\ram[156][7] ), .B(\ram[157][7] ), .C(\ram[158][7] ), .D(
        \ram[159][7] ), .S0(n6307), .S1(n6173), .Y(n5292) );
  MX4X1 U6391 ( .A(\ram[172][7] ), .B(\ram[173][7] ), .C(\ram[174][7] ), .D(
        \ram[175][7] ), .S0(n6306), .S1(n6172), .Y(n5287) );
  MX4X1 U6392 ( .A(\ram[140][7] ), .B(\ram[141][7] ), .C(\ram[142][7] ), .D(
        \ram[143][7] ), .S0(n6307), .S1(n6173), .Y(n5297) );
  MX4X1 U6393 ( .A(\ram[60][7] ), .B(\ram[61][7] ), .C(\ram[62][7] ), .D(
        \ram[63][7] ), .S0(n6309), .S1(n6175), .Y(n5324) );
  MX4X1 U6394 ( .A(\ram[28][7] ), .B(\ram[29][7] ), .C(\ram[30][7] ), .D(
        \ram[31][7] ), .S0(n6309), .S1(n6175), .Y(n5334) );
  MX4X1 U6395 ( .A(\ram[44][7] ), .B(\ram[45][7] ), .C(\ram[46][7] ), .D(
        \ram[47][7] ), .S0(n6309), .S1(n6175), .Y(n5329) );
  MX4X1 U6396 ( .A(\ram[12][7] ), .B(\ram[13][7] ), .C(\ram[14][7] ), .D(
        \ram[15][7] ), .S0(n6310), .S1(n6176), .Y(n5339) );
  MX4X1 U6397 ( .A(\ram[252][8] ), .B(\ram[253][8] ), .C(\ram[254][8] ), .D(
        \ram[255][8] ), .S0(n6310), .S1(n6176), .Y(n5345) );
  MX4X1 U6398 ( .A(\ram[220][8] ), .B(\ram[221][8] ), .C(\ram[222][8] ), .D(
        \ram[223][8] ), .S0(n6311), .S1(n6177), .Y(n5355) );
  MX4X1 U6399 ( .A(\ram[236][8] ), .B(\ram[237][8] ), .C(\ram[238][8] ), .D(
        \ram[239][8] ), .S0(n6310), .S1(n6176), .Y(n5350) );
  MX4X1 U6400 ( .A(\ram[204][8] ), .B(\ram[205][8] ), .C(\ram[206][8] ), .D(
        \ram[207][8] ), .S0(n6311), .S1(n6177), .Y(n5360) );
  MX4X1 U6401 ( .A(\ram[124][8] ), .B(\ram[125][8] ), .C(\ram[126][8] ), .D(
        \ram[127][8] ), .S0(n6313), .S1(n6179), .Y(n5387) );
  MX4X1 U6402 ( .A(\ram[92][8] ), .B(\ram[93][8] ), .C(\ram[94][8] ), .D(
        \ram[95][8] ), .S0(n6313), .S1(n6179), .Y(n5397) );
  MX4X1 U6403 ( .A(\ram[108][8] ), .B(\ram[109][8] ), .C(\ram[110][8] ), .D(
        \ram[111][8] ), .S0(n6313), .S1(n6179), .Y(n5392) );
  MX4X1 U6404 ( .A(\ram[76][8] ), .B(\ram[77][8] ), .C(\ram[78][8] ), .D(
        \ram[79][8] ), .S0(n6314), .S1(n6180), .Y(n5402) );
  MX4X1 U6405 ( .A(\ram[188][8] ), .B(\ram[189][8] ), .C(\ram[190][8] ), .D(
        \ram[191][8] ), .S0(n6311), .S1(n6177), .Y(n5366) );
  MX4X1 U6406 ( .A(\ram[156][8] ), .B(\ram[157][8] ), .C(\ram[158][8] ), .D(
        \ram[159][8] ), .S0(n6312), .S1(n6178), .Y(n5376) );
  MX4X1 U6407 ( .A(\ram[172][8] ), .B(\ram[173][8] ), .C(\ram[174][8] ), .D(
        \ram[175][8] ), .S0(n6312), .S1(n6178), .Y(n5371) );
  MX4X1 U6408 ( .A(\ram[140][8] ), .B(\ram[141][8] ), .C(\ram[142][8] ), .D(
        \ram[143][8] ), .S0(n6312), .S1(n6178), .Y(n5381) );
  MX4X1 U6409 ( .A(\ram[60][8] ), .B(\ram[61][8] ), .C(\ram[62][8] ), .D(
        \ram[63][8] ), .S0(n6314), .S1(n6180), .Y(n5408) );
  MX4X1 U6410 ( .A(\ram[28][8] ), .B(\ram[29][8] ), .C(\ram[30][8] ), .D(
        \ram[31][8] ), .S0(n6315), .S1(n6181), .Y(n5418) );
  MX4X1 U6411 ( .A(\ram[44][8] ), .B(\ram[45][8] ), .C(\ram[46][8] ), .D(
        \ram[47][8] ), .S0(n6314), .S1(n6180), .Y(n5413) );
  MX4X1 U6412 ( .A(\ram[12][8] ), .B(\ram[13][8] ), .C(\ram[14][8] ), .D(
        \ram[15][8] ), .S0(n6315), .S1(n6181), .Y(n5423) );
  MX4X1 U6413 ( .A(\ram[252][9] ), .B(\ram[253][9] ), .C(\ram[254][9] ), .D(
        \ram[255][9] ), .S0(n6315), .S1(n6181), .Y(n5429) );
  MX4X1 U6414 ( .A(\ram[220][9] ), .B(\ram[221][9] ), .C(\ram[222][9] ), .D(
        \ram[223][9] ), .S0(n6316), .S1(n6182), .Y(n5439) );
  MX4X1 U6415 ( .A(\ram[236][9] ), .B(\ram[237][9] ), .C(\ram[238][9] ), .D(
        \ram[239][9] ), .S0(n6316), .S1(n6182), .Y(n5434) );
  MX4X1 U6416 ( .A(\ram[204][9] ), .B(\ram[205][9] ), .C(\ram[206][9] ), .D(
        \ram[207][9] ), .S0(n6316), .S1(n6182), .Y(n5444) );
  MX4X1 U6417 ( .A(\ram[124][9] ), .B(\ram[125][9] ), .C(\ram[126][9] ), .D(
        \ram[127][9] ), .S0(n6318), .S1(n6184), .Y(n5471) );
  MX4X1 U6418 ( .A(\ram[92][9] ), .B(\ram[93][9] ), .C(\ram[94][9] ), .D(
        \ram[95][9] ), .S0(n6319), .S1(n6185), .Y(n5481) );
  MX4X1 U6419 ( .A(\ram[108][9] ), .B(\ram[109][9] ), .C(\ram[110][9] ), .D(
        \ram[111][9] ), .S0(n6318), .S1(n6184), .Y(n5476) );
  MX4X1 U6420 ( .A(\ram[76][9] ), .B(\ram[77][9] ), .C(\ram[78][9] ), .D(
        \ram[79][9] ), .S0(n6319), .S1(n6185), .Y(n5486) );
  MX4X1 U6421 ( .A(\ram[188][9] ), .B(\ram[189][9] ), .C(\ram[190][9] ), .D(
        \ram[191][9] ), .S0(n6317), .S1(n6183), .Y(n5450) );
  MX4X1 U6422 ( .A(\ram[156][9] ), .B(\ram[157][9] ), .C(\ram[158][9] ), .D(
        \ram[159][9] ), .S0(n6317), .S1(n6183), .Y(n5460) );
  MX4X1 U6423 ( .A(\ram[172][9] ), .B(\ram[173][9] ), .C(\ram[174][9] ), .D(
        \ram[175][9] ), .S0(n6317), .S1(n6183), .Y(n5455) );
  MX4X1 U6424 ( .A(\ram[140][9] ), .B(\ram[141][9] ), .C(\ram[142][9] ), .D(
        \ram[143][9] ), .S0(n6318), .S1(n6184), .Y(n5465) );
  MX4X1 U6425 ( .A(\ram[60][9] ), .B(\ram[61][9] ), .C(\ram[62][9] ), .D(
        \ram[63][9] ), .S0(n6319), .S1(n6185), .Y(n5492) );
  MX4X1 U6426 ( .A(\ram[28][9] ), .B(\ram[29][9] ), .C(\ram[30][9] ), .D(
        \ram[31][9] ), .S0(n6320), .S1(n6186), .Y(n5502) );
  MX4X1 U6427 ( .A(\ram[44][9] ), .B(\ram[45][9] ), .C(\ram[46][9] ), .D(
        \ram[47][9] ), .S0(n6320), .S1(n6186), .Y(n5497) );
  MX4X1 U6428 ( .A(\ram[12][9] ), .B(\ram[13][9] ), .C(\ram[14][9] ), .D(
        \ram[15][9] ), .S0(n6320), .S1(n6186), .Y(n5507) );
  MX4X1 U6429 ( .A(\ram[252][10] ), .B(\ram[253][10] ), .C(\ram[254][10] ), 
        .D(\ram[255][10] ), .S0(n6321), .S1(n6187), .Y(n5513) );
  MX4X1 U6430 ( .A(\ram[220][10] ), .B(\ram[221][10] ), .C(\ram[222][10] ), 
        .D(\ram[223][10] ), .S0(n6321), .S1(n6187), .Y(n5523) );
  MX4X1 U6431 ( .A(\ram[236][10] ), .B(\ram[237][10] ), .C(\ram[238][10] ), 
        .D(\ram[239][10] ), .S0(n6321), .S1(n6187), .Y(n5518) );
  MX4X1 U6432 ( .A(\ram[204][10] ), .B(\ram[205][10] ), .C(\ram[206][10] ), 
        .D(\ram[207][10] ), .S0(n6322), .S1(n6188), .Y(n5528) );
  MX4X1 U6433 ( .A(\ram[188][10] ), .B(\ram[189][10] ), .C(\ram[190][10] ), 
        .D(\ram[191][10] ), .S0(n6322), .S1(n6188), .Y(n5534) );
  MX4X1 U6434 ( .A(\ram[172][10] ), .B(\ram[173][10] ), .C(\ram[174][10] ), 
        .D(\ram[175][10] ), .S0(n6322), .S1(n6188), .Y(n5539) );
  MX4X1 U6435 ( .A(\ram[156][10] ), .B(\ram[157][10] ), .C(\ram[158][10] ), 
        .D(\ram[159][10] ), .S0(n6323), .S1(n6189), .Y(n5544) );
  MX4X1 U6436 ( .A(\ram[140][10] ), .B(\ram[141][10] ), .C(\ram[142][10] ), 
        .D(\ram[143][10] ), .S0(n6323), .S1(n6189), .Y(n5549) );
  MX4X1 U6437 ( .A(\ram[124][10] ), .B(\ram[125][10] ), .C(\ram[126][10] ), 
        .D(\ram[127][10] ), .S0(n6323), .S1(n6189), .Y(n5555) );
  MX4X1 U6438 ( .A(\ram[92][10] ), .B(\ram[93][10] ), .C(\ram[94][10] ), .D(
        \ram[95][10] ), .S0(n6324), .S1(n6190), .Y(n5565) );
  MX4X1 U6439 ( .A(\ram[108][10] ), .B(\ram[109][10] ), .C(\ram[110][10] ), 
        .D(\ram[111][10] ), .S0(n6324), .S1(n6190), .Y(n5560) );
  MX4X1 U6440 ( .A(\ram[76][10] ), .B(\ram[77][10] ), .C(\ram[78][10] ), .D(
        \ram[79][10] ), .S0(n6324), .S1(n6190), .Y(n5570) );
  MX4X1 U6441 ( .A(\ram[60][10] ), .B(\ram[61][10] ), .C(\ram[62][10] ), .D(
        \ram[63][10] ), .S0(n6325), .S1(n6191), .Y(n5576) );
  MX4X1 U6442 ( .A(\ram[28][10] ), .B(\ram[29][10] ), .C(\ram[30][10] ), .D(
        \ram[31][10] ), .S0(n6325), .S1(n6191), .Y(n5586) );
  MX4X1 U6443 ( .A(\ram[44][10] ), .B(\ram[45][10] ), .C(\ram[46][10] ), .D(
        \ram[47][10] ), .S0(n6325), .S1(n6191), .Y(n5581) );
  MX4X1 U6444 ( .A(\ram[12][10] ), .B(\ram[13][10] ), .C(\ram[14][10] ), .D(
        \ram[15][10] ), .S0(n6326), .S1(n6192), .Y(n5591) );
  MX4X1 U6445 ( .A(\ram[252][11] ), .B(\ram[253][11] ), .C(\ram[254][11] ), 
        .D(\ram[255][11] ), .S0(n6326), .S1(n6192), .Y(n5597) );
  MX4X1 U6446 ( .A(\ram[220][11] ), .B(\ram[221][11] ), .C(\ram[222][11] ), 
        .D(\ram[223][11] ), .S0(n6327), .S1(n6193), .Y(n5607) );
  MX4X1 U6447 ( .A(\ram[236][11] ), .B(\ram[237][11] ), .C(\ram[238][11] ), 
        .D(\ram[239][11] ), .S0(n6326), .S1(n6192), .Y(n5602) );
  MX4X1 U6448 ( .A(\ram[204][11] ), .B(\ram[205][11] ), .C(\ram[206][11] ), 
        .D(\ram[207][11] ), .S0(n6327), .S1(n6193), .Y(n5612) );
  MX4X1 U6449 ( .A(\ram[124][11] ), .B(\ram[125][11] ), .C(\ram[126][11] ), 
        .D(\ram[127][11] ), .S0(n6329), .S1(n6195), .Y(n5639) );
  MX4X1 U6450 ( .A(\ram[92][11] ), .B(\ram[93][11] ), .C(\ram[94][11] ), .D(
        \ram[95][11] ), .S0(n6329), .S1(n6195), .Y(n5649) );
  MX4X1 U6451 ( .A(\ram[108][11] ), .B(\ram[109][11] ), .C(\ram[110][11] ), 
        .D(\ram[111][11] ), .S0(n6329), .S1(n6195), .Y(n5644) );
  MX4X1 U6452 ( .A(\ram[76][11] ), .B(\ram[77][11] ), .C(\ram[78][11] ), .D(
        \ram[79][11] ), .S0(n6330), .S1(n6196), .Y(n5654) );
  MX4X1 U6453 ( .A(\ram[188][11] ), .B(\ram[189][11] ), .C(\ram[190][11] ), 
        .D(\ram[191][11] ), .S0(n6327), .S1(n6193), .Y(n5618) );
  MX4X1 U6454 ( .A(\ram[156][11] ), .B(\ram[157][11] ), .C(\ram[158][11] ), 
        .D(\ram[159][11] ), .S0(n6328), .S1(n6194), .Y(n5628) );
  MX4X1 U6455 ( .A(\ram[172][11] ), .B(\ram[173][11] ), .C(\ram[174][11] ), 
        .D(\ram[175][11] ), .S0(n6328), .S1(n6194), .Y(n5623) );
  MX4X1 U6456 ( .A(\ram[140][11] ), .B(\ram[141][11] ), .C(\ram[142][11] ), 
        .D(\ram[143][11] ), .S0(n6328), .S1(n6194), .Y(n5633) );
  MX4X1 U6457 ( .A(\ram[60][11] ), .B(\ram[61][11] ), .C(\ram[62][11] ), .D(
        \ram[63][11] ), .S0(n6330), .S1(n6196), .Y(n5660) );
  MX4X1 U6458 ( .A(\ram[28][11] ), .B(\ram[29][11] ), .C(\ram[30][11] ), .D(
        \ram[31][11] ), .S0(n6331), .S1(n6197), .Y(n5670) );
  MX4X1 U6459 ( .A(\ram[44][11] ), .B(\ram[45][11] ), .C(\ram[46][11] ), .D(
        \ram[47][11] ), .S0(n6330), .S1(n6196), .Y(n5665) );
  MX4X1 U6460 ( .A(\ram[12][11] ), .B(\ram[13][11] ), .C(\ram[14][11] ), .D(
        \ram[15][11] ), .S0(n6331), .S1(n6197), .Y(n5675) );
  MX4X1 U6461 ( .A(\ram[252][12] ), .B(\ram[253][12] ), .C(\ram[254][12] ), 
        .D(\ram[255][12] ), .S0(n6331), .S1(n6197), .Y(n5681) );
  MX4X1 U6462 ( .A(\ram[220][12] ), .B(\ram[221][12] ), .C(\ram[222][12] ), 
        .D(\ram[223][12] ), .S0(n6332), .S1(n6198), .Y(n5691) );
  MX4X1 U6463 ( .A(\ram[236][12] ), .B(\ram[237][12] ), .C(\ram[238][12] ), 
        .D(\ram[239][12] ), .S0(n6332), .S1(n6198), .Y(n5686) );
  MX4X1 U6464 ( .A(\ram[204][12] ), .B(\ram[205][12] ), .C(\ram[206][12] ), 
        .D(\ram[207][12] ), .S0(n6332), .S1(n6198), .Y(n5696) );
  MX4X1 U6465 ( .A(\ram[124][12] ), .B(\ram[125][12] ), .C(\ram[126][12] ), 
        .D(\ram[127][12] ), .S0(n6334), .S1(n6200), .Y(n5723) );
  MX4X1 U6466 ( .A(\ram[92][12] ), .B(\ram[93][12] ), .C(\ram[94][12] ), .D(
        \ram[95][12] ), .S0(n6335), .S1(n6201), .Y(n5733) );
  MX4X1 U6467 ( .A(\ram[108][12] ), .B(\ram[109][12] ), .C(\ram[110][12] ), 
        .D(\ram[111][12] ), .S0(n6334), .S1(n6200), .Y(n5728) );
  MX4X1 U6468 ( .A(\ram[76][12] ), .B(\ram[77][12] ), .C(\ram[78][12] ), .D(
        \ram[79][12] ), .S0(n6335), .S1(n6201), .Y(n5738) );
  MX4X1 U6469 ( .A(\ram[188][12] ), .B(\ram[189][12] ), .C(\ram[190][12] ), 
        .D(\ram[191][12] ), .S0(n6333), .S1(n6199), .Y(n5702) );
  MX4X1 U6470 ( .A(\ram[156][12] ), .B(\ram[157][12] ), .C(\ram[158][12] ), 
        .D(\ram[159][12] ), .S0(n6333), .S1(n6199), .Y(n5712) );
  MX4X1 U6471 ( .A(\ram[172][12] ), .B(\ram[173][12] ), .C(\ram[174][12] ), 
        .D(\ram[175][12] ), .S0(n6333), .S1(n6199), .Y(n5707) );
  MX4X1 U6472 ( .A(\ram[140][12] ), .B(\ram[141][12] ), .C(\ram[142][12] ), 
        .D(\ram[143][12] ), .S0(n6334), .S1(n6200), .Y(n5717) );
  MX4X1 U6473 ( .A(\ram[60][12] ), .B(\ram[61][12] ), .C(\ram[62][12] ), .D(
        \ram[63][12] ), .S0(n6335), .S1(n6201), .Y(n5744) );
  MX4X1 U6474 ( .A(\ram[28][12] ), .B(\ram[29][12] ), .C(\ram[30][12] ), .D(
        \ram[31][12] ), .S0(n6336), .S1(n6202), .Y(n5754) );
  MX4X1 U6475 ( .A(\ram[44][12] ), .B(\ram[45][12] ), .C(\ram[46][12] ), .D(
        \ram[47][12] ), .S0(n6336), .S1(n6202), .Y(n5749) );
  MX4X1 U6476 ( .A(\ram[12][12] ), .B(\ram[13][12] ), .C(\ram[14][12] ), .D(
        \ram[15][12] ), .S0(n6336), .S1(n6202), .Y(n5759) );
  MX4X1 U6477 ( .A(\ram[252][13] ), .B(\ram[253][13] ), .C(\ram[254][13] ), 
        .D(\ram[255][13] ), .S0(n6337), .S1(n6203), .Y(n5765) );
  MX4X1 U6478 ( .A(\ram[220][13] ), .B(\ram[221][13] ), .C(\ram[222][13] ), 
        .D(\ram[223][13] ), .S0(n6337), .S1(n6203), .Y(n5775) );
  MX4X1 U6479 ( .A(\ram[236][13] ), .B(\ram[237][13] ), .C(\ram[238][13] ), 
        .D(\ram[239][13] ), .S0(n6337), .S1(n6203), .Y(n5770) );
  MX4X1 U6480 ( .A(\ram[204][13] ), .B(\ram[205][13] ), .C(\ram[206][13] ), 
        .D(\ram[207][13] ), .S0(n6338), .S1(n6204), .Y(n5780) );
  MX4X1 U6481 ( .A(\ram[124][13] ), .B(\ram[125][13] ), .C(\ram[126][13] ), 
        .D(\ram[127][13] ), .S0(n6339), .S1(n6205), .Y(n5807) );
  MX4X1 U6482 ( .A(\ram[92][13] ), .B(\ram[93][13] ), .C(\ram[94][13] ), .D(
        \ram[95][13] ), .S0(n6340), .S1(n6206), .Y(n5817) );
  MX4X1 U6483 ( .A(\ram[108][13] ), .B(\ram[109][13] ), .C(\ram[110][13] ), 
        .D(\ram[111][13] ), .S0(n6340), .S1(n6206), .Y(n5812) );
  MX4X1 U6484 ( .A(\ram[76][13] ), .B(\ram[77][13] ), .C(\ram[78][13] ), .D(
        \ram[79][13] ), .S0(n6340), .S1(n6206), .Y(n5822) );
  MX4X1 U6485 ( .A(\ram[188][13] ), .B(\ram[189][13] ), .C(\ram[190][13] ), 
        .D(\ram[191][13] ), .S0(n6338), .S1(n6204), .Y(n5786) );
  MX4X1 U6486 ( .A(\ram[156][13] ), .B(\ram[157][13] ), .C(\ram[158][13] ), 
        .D(\ram[159][13] ), .S0(n6339), .S1(n6205), .Y(n5796) );
  MX4X1 U6487 ( .A(\ram[172][13] ), .B(\ram[173][13] ), .C(\ram[174][13] ), 
        .D(\ram[175][13] ), .S0(n6338), .S1(n6204), .Y(n5791) );
  MX4X1 U6488 ( .A(\ram[140][13] ), .B(\ram[141][13] ), .C(\ram[142][13] ), 
        .D(\ram[143][13] ), .S0(n6339), .S1(n6205), .Y(n5801) );
  MX4X1 U6489 ( .A(\ram[60][13] ), .B(\ram[61][13] ), .C(\ram[62][13] ), .D(
        \ram[63][13] ), .S0(n6341), .S1(n6207), .Y(n5828) );
  MX4X1 U6490 ( .A(\ram[28][13] ), .B(\ram[29][13] ), .C(\ram[30][13] ), .D(
        \ram[31][13] ), .S0(n6341), .S1(n6207), .Y(n5838) );
  MX4X1 U6491 ( .A(\ram[44][13] ), .B(\ram[45][13] ), .C(\ram[46][13] ), .D(
        \ram[47][13] ), .S0(n6341), .S1(n6207), .Y(n5833) );
  MX4X1 U6492 ( .A(\ram[12][13] ), .B(\ram[13][13] ), .C(\ram[14][13] ), .D(
        \ram[15][13] ), .S0(n6342), .S1(n6208), .Y(n5843) );
  MX4X1 U6493 ( .A(\ram[252][14] ), .B(\ram[253][14] ), .C(\ram[254][14] ), 
        .D(\ram[255][14] ), .S0(n6342), .S1(n6208), .Y(n5849) );
  MX4X1 U6494 ( .A(\ram[220][14] ), .B(\ram[221][14] ), .C(\ram[222][14] ), 
        .D(\ram[223][14] ), .S0(n6343), .S1(n6209), .Y(n5859) );
  MX4X1 U6495 ( .A(\ram[236][14] ), .B(\ram[237][14] ), .C(\ram[238][14] ), 
        .D(\ram[239][14] ), .S0(n6342), .S1(n6208), .Y(n5854) );
  MX4X1 U6496 ( .A(\ram[204][14] ), .B(\ram[205][14] ), .C(\ram[206][14] ), 
        .D(\ram[207][14] ), .S0(n6343), .S1(n6209), .Y(n5864) );
  MX4X1 U6497 ( .A(\ram[124][14] ), .B(\ram[125][14] ), .C(\ram[126][14] ), 
        .D(\ram[127][14] ), .S0(n6345), .S1(n6211), .Y(n5891) );
  MX4X1 U6498 ( .A(\ram[92][14] ), .B(\ram[93][14] ), .C(\ram[94][14] ), .D(
        \ram[95][14] ), .S0(n6345), .S1(n6211), .Y(n5901) );
  MX4X1 U6499 ( .A(\ram[108][14] ), .B(\ram[109][14] ), .C(\ram[110][14] ), 
        .D(\ram[111][14] ), .S0(n6345), .S1(n6211), .Y(n5896) );
  MX4X1 U6500 ( .A(\ram[76][14] ), .B(\ram[77][14] ), .C(\ram[78][14] ), .D(
        \ram[79][14] ), .S0(n6346), .S1(n6212), .Y(n5906) );
  MX4X1 U6501 ( .A(\ram[188][14] ), .B(\ram[189][14] ), .C(\ram[190][14] ), 
        .D(\ram[191][14] ), .S0(n6343), .S1(n6209), .Y(n5870) );
  MX4X1 U6502 ( .A(\ram[156][14] ), .B(\ram[157][14] ), .C(\ram[158][14] ), 
        .D(\ram[159][14] ), .S0(n6344), .S1(n6210), .Y(n5880) );
  MX4X1 U6503 ( .A(\ram[172][14] ), .B(\ram[173][14] ), .C(\ram[174][14] ), 
        .D(\ram[175][14] ), .S0(n6344), .S1(n6210), .Y(n5875) );
  MX4X1 U6504 ( .A(\ram[140][14] ), .B(\ram[141][14] ), .C(\ram[142][14] ), 
        .D(\ram[143][14] ), .S0(n6344), .S1(n6210), .Y(n5885) );
  MX4X1 U6505 ( .A(\ram[60][14] ), .B(\ram[61][14] ), .C(\ram[62][14] ), .D(
        \ram[63][14] ), .S0(n6346), .S1(n6212), .Y(n5912) );
  MX4X1 U6506 ( .A(\ram[44][14] ), .B(\ram[45][14] ), .C(\ram[46][14] ), .D(
        \ram[47][14] ), .S0(n6346), .S1(n6212), .Y(n5917) );
  MX4X1 U6507 ( .A(\ram[28][14] ), .B(\ram[29][14] ), .C(\ram[30][14] ), .D(
        \ram[31][14] ), .S0(n6347), .S1(n6140), .Y(n5922) );
  MX4X1 U6508 ( .A(\ram[12][14] ), .B(\ram[13][14] ), .C(\ram[14][14] ), .D(
        \ram[15][14] ), .S0(n6347), .S1(n6155), .Y(n5927) );
  MX4X1 U6509 ( .A(\ram[252][15] ), .B(\ram[253][15] ), .C(\ram[254][15] ), 
        .D(\ram[255][15] ), .S0(n6347), .S1(n6092), .Y(n5933) );
  MX4X1 U6510 ( .A(\ram[220][15] ), .B(\ram[221][15] ), .C(\ram[222][15] ), 
        .D(\ram[223][15] ), .S0(n6348), .S1(n6213), .Y(n5943) );
  MX4X1 U6511 ( .A(\ram[236][15] ), .B(\ram[237][15] ), .C(\ram[238][15] ), 
        .D(\ram[239][15] ), .S0(n6348), .S1(n6213), .Y(n5938) );
  MX4X1 U6512 ( .A(\ram[204][15] ), .B(\ram[205][15] ), .C(\ram[206][15] ), 
        .D(\ram[207][15] ), .S0(n6348), .S1(n6213), .Y(n5948) );
  MX4X1 U6513 ( .A(\ram[124][15] ), .B(\ram[125][15] ), .C(\ram[126][15] ), 
        .D(\ram[127][15] ), .S0(n6350), .S1(n6213), .Y(n5975) );
  MX4X1 U6514 ( .A(\ram[92][15] ), .B(\ram[93][15] ), .C(\ram[94][15] ), .D(
        \ram[95][15] ), .S0(n6351), .S1(n6091), .Y(n5985) );
  MX4X1 U6515 ( .A(\ram[108][15] ), .B(\ram[109][15] ), .C(\ram[110][15] ), 
        .D(\ram[111][15] ), .S0(n6350), .S1(n6139), .Y(n5980) );
  MX4X1 U6516 ( .A(\ram[76][15] ), .B(\ram[77][15] ), .C(\ram[78][15] ), .D(
        \ram[79][15] ), .S0(n6351), .S1(n6192), .Y(n5990) );
  MX4X1 U6517 ( .A(\ram[188][15] ), .B(\ram[189][15] ), .C(\ram[190][15] ), 
        .D(\ram[191][15] ), .S0(n6349), .S1(n6214), .Y(n5954) );
  MX4X1 U6518 ( .A(\ram[156][15] ), .B(\ram[157][15] ), .C(\ram[158][15] ), 
        .D(\ram[159][15] ), .S0(n6349), .S1(n6214), .Y(n5964) );
  MX4X1 U6519 ( .A(\ram[172][15] ), .B(\ram[173][15] ), .C(\ram[174][15] ), 
        .D(\ram[175][15] ), .S0(n6349), .S1(n6214), .Y(n5959) );
  MX4X1 U6520 ( .A(\ram[140][15] ), .B(\ram[141][15] ), .C(\ram[142][15] ), 
        .D(\ram[143][15] ), .S0(n6350), .S1(n6214), .Y(n5969) );
  MX4X1 U6521 ( .A(\ram[60][15] ), .B(\ram[61][15] ), .C(\ram[62][15] ), .D(
        \ram[63][15] ), .S0(n6351), .S1(n6190), .Y(n5996) );
  MX4X1 U6522 ( .A(\ram[28][15] ), .B(\ram[29][15] ), .C(\ram[30][15] ), .D(
        \ram[31][15] ), .S0(n6352), .S1(n6191), .Y(n6006) );
  MX4X1 U6523 ( .A(\ram[44][15] ), .B(\ram[45][15] ), .C(\ram[46][15] ), .D(
        \ram[47][15] ), .S0(n6352), .S1(n6139), .Y(n6001) );
  MX4X1 U6524 ( .A(\ram[12][15] ), .B(\ram[13][15] ), .C(\ram[14][15] ), .D(
        \ram[15][15] ), .S0(n6352), .S1(n6189), .Y(n6011) );
  MX4X1 U6525 ( .A(n4718), .B(n4716), .C(n4717), .D(n4715), .S0(n6037), .S1(
        n6061), .Y(n4719) );
  MX4X1 U6526 ( .A(\ram[112][0] ), .B(\ram[113][0] ), .C(\ram[114][0] ), .D(
        \ram[115][0] ), .S0(n6270), .S1(n6136), .Y(n4718) );
  MX4X1 U6527 ( .A(\ram[120][0] ), .B(\ram[121][0] ), .C(\ram[122][0] ), .D(
        \ram[123][0] ), .S0(n6270), .S1(n6136), .Y(n4716) );
  MX4X1 U6528 ( .A(\ram[116][0] ), .B(\ram[117][0] ), .C(\ram[118][0] ), .D(
        \ram[119][0] ), .S0(n6270), .S1(n6136), .Y(n4717) );
  MX4X1 U6529 ( .A(n4697), .B(n4695), .C(n4696), .D(n4694), .S0(n6041), .S1(
        n6057), .Y(n4698) );
  MX4X1 U6530 ( .A(\ram[176][0] ), .B(\ram[177][0] ), .C(\ram[178][0] ), .D(
        \ram[179][0] ), .S0(n6269), .S1(n6135), .Y(n4697) );
  MX4X1 U6531 ( .A(\ram[184][0] ), .B(\ram[185][0] ), .C(\ram[186][0] ), .D(
        \ram[187][0] ), .S0(n6269), .S1(n6135), .Y(n4695) );
  MX4X1 U6532 ( .A(\ram[180][0] ), .B(\ram[181][0] ), .C(\ram[182][0] ), .D(
        \ram[183][0] ), .S0(n6269), .S1(n6135), .Y(n4696) );
  MX4X1 U6533 ( .A(n4739), .B(n4737), .C(n4738), .D(n4736), .S0(n6033), .S1(
        n6056), .Y(n4740) );
  MX4X1 U6534 ( .A(\ram[48][0] ), .B(\ram[49][0] ), .C(\ram[50][0] ), .D(
        \ram[51][0] ), .S0(n6271), .S1(n6137), .Y(n4739) );
  MX4X1 U6535 ( .A(\ram[56][0] ), .B(\ram[57][0] ), .C(\ram[58][0] ), .D(
        \ram[59][0] ), .S0(n6271), .S1(n6137), .Y(n4737) );
  MX4X1 U6536 ( .A(\ram[52][0] ), .B(\ram[53][0] ), .C(\ram[54][0] ), .D(
        \ram[55][0] ), .S0(n6271), .S1(n6137), .Y(n4738) );
  MX4X1 U6537 ( .A(n4760), .B(n4758), .C(n4759), .D(n4757), .S0(n6033), .S1(
        n6056), .Y(n4761) );
  MX4X1 U6538 ( .A(\ram[240][1] ), .B(\ram[241][1] ), .C(\ram[242][1] ), .D(
        \ram[243][1] ), .S0(n6273), .S1(n6139), .Y(n4760) );
  MX4X1 U6539 ( .A(\ram[248][1] ), .B(\ram[249][1] ), .C(\ram[250][1] ), .D(
        \ram[251][1] ), .S0(n6273), .S1(n6139), .Y(n4758) );
  MX4X1 U6540 ( .A(\ram[244][1] ), .B(\ram[245][1] ), .C(\ram[246][1] ), .D(
        \ram[247][1] ), .S0(n6273), .S1(n6139), .Y(n4759) );
  MX4X1 U6541 ( .A(n4802), .B(n4800), .C(n4801), .D(n4799), .S0(n6033), .S1(
        n6056), .Y(n4803) );
  MX4X1 U6542 ( .A(\ram[112][1] ), .B(\ram[113][1] ), .C(\ram[114][1] ), .D(
        \ram[115][1] ), .S0(n6275), .S1(n6141), .Y(n4802) );
  MX4X1 U6543 ( .A(\ram[120][1] ), .B(\ram[121][1] ), .C(\ram[122][1] ), .D(
        \ram[123][1] ), .S0(n6275), .S1(n6141), .Y(n4800) );
  MX4X1 U6544 ( .A(\ram[116][1] ), .B(\ram[117][1] ), .C(\ram[118][1] ), .D(
        \ram[119][1] ), .S0(n6275), .S1(n6141), .Y(n4801) );
  MX4X1 U6545 ( .A(n4781), .B(n4779), .C(n4780), .D(n4778), .S0(n6033), .S1(
        n6056), .Y(n4782) );
  MX4X1 U6546 ( .A(\ram[176][1] ), .B(\ram[177][1] ), .C(\ram[178][1] ), .D(
        \ram[179][1] ), .S0(n6274), .S1(n6140), .Y(n4781) );
  MX4X1 U6547 ( .A(\ram[184][1] ), .B(\ram[185][1] ), .C(\ram[186][1] ), .D(
        \ram[187][1] ), .S0(n6274), .S1(n6140), .Y(n4779) );
  MX4X1 U6548 ( .A(\ram[180][1] ), .B(\ram[181][1] ), .C(\ram[182][1] ), .D(
        \ram[183][1] ), .S0(n6274), .S1(n6140), .Y(n4780) );
  MX4X1 U6549 ( .A(n4823), .B(n4821), .C(n4822), .D(n4820), .S0(n6046), .S1(
        n6057), .Y(n4824) );
  MX4X1 U6550 ( .A(\ram[48][1] ), .B(\ram[49][1] ), .C(\ram[50][1] ), .D(
        \ram[51][1] ), .S0(n6277), .S1(n6143), .Y(n4823) );
  MX4X1 U6551 ( .A(\ram[56][1] ), .B(\ram[57][1] ), .C(\ram[58][1] ), .D(
        \ram[59][1] ), .S0(n6277), .S1(n6143), .Y(n4821) );
  MX4X1 U6552 ( .A(\ram[52][1] ), .B(\ram[53][1] ), .C(\ram[54][1] ), .D(
        \ram[55][1] ), .S0(n6277), .S1(n6143), .Y(n4822) );
  MX4X1 U6553 ( .A(n4844), .B(n4842), .C(n4843), .D(n4841), .S0(n6036), .S1(
        n6057), .Y(n4845) );
  MX4X1 U6554 ( .A(\ram[240][2] ), .B(\ram[241][2] ), .C(\ram[242][2] ), .D(
        \ram[243][2] ), .S0(n6278), .S1(n6144), .Y(n4844) );
  MX4X1 U6555 ( .A(\ram[248][2] ), .B(\ram[249][2] ), .C(\ram[250][2] ), .D(
        \ram[251][2] ), .S0(n6278), .S1(n6144), .Y(n4842) );
  MX4X1 U6556 ( .A(\ram[244][2] ), .B(\ram[245][2] ), .C(\ram[246][2] ), .D(
        \ram[247][2] ), .S0(n6278), .S1(n6144), .Y(n4843) );
  MX4X1 U6557 ( .A(n4886), .B(n4884), .C(n4885), .D(n4883), .S0(n6044), .S1(
        n6058), .Y(n4887) );
  MX4X1 U6558 ( .A(\ram[112][2] ), .B(\ram[113][2] ), .C(\ram[114][2] ), .D(
        \ram[115][2] ), .S0(n6281), .S1(n6147), .Y(n4886) );
  MX4X1 U6559 ( .A(\ram[120][2] ), .B(\ram[121][2] ), .C(\ram[122][2] ), .D(
        \ram[123][2] ), .S0(n6281), .S1(n6147), .Y(n4884) );
  MX4X1 U6560 ( .A(\ram[116][2] ), .B(\ram[117][2] ), .C(\ram[118][2] ), .D(
        \ram[119][2] ), .S0(n6281), .S1(n6147), .Y(n4885) );
  MX4X1 U6561 ( .A(n4865), .B(n4863), .C(n4864), .D(n4862), .S0(n6040), .S1(
        n6057), .Y(n4866) );
  MX4X1 U6562 ( .A(\ram[176][2] ), .B(\ram[177][2] ), .C(\ram[178][2] ), .D(
        \ram[179][2] ), .S0(n6279), .S1(n6145), .Y(n4865) );
  MX4X1 U6563 ( .A(\ram[184][2] ), .B(\ram[185][2] ), .C(\ram[186][2] ), .D(
        \ram[187][2] ), .S0(n6279), .S1(n6145), .Y(n4863) );
  MX4X1 U6564 ( .A(\ram[180][2] ), .B(\ram[181][2] ), .C(\ram[182][2] ), .D(
        \ram[183][2] ), .S0(n6279), .S1(n6145), .Y(n4864) );
  MX4X1 U6565 ( .A(n4907), .B(n4905), .C(n4906), .D(n4904), .S0(n6037), .S1(
        n6058), .Y(n4908) );
  MX4X1 U6566 ( .A(\ram[48][2] ), .B(\ram[49][2] ), .C(\ram[50][2] ), .D(
        \ram[51][2] ), .S0(n6282), .S1(n6148), .Y(n4907) );
  MX4X1 U6567 ( .A(\ram[56][2] ), .B(\ram[57][2] ), .C(\ram[58][2] ), .D(
        \ram[59][2] ), .S0(n6282), .S1(n6148), .Y(n4905) );
  MX4X1 U6568 ( .A(\ram[52][2] ), .B(\ram[53][2] ), .C(\ram[54][2] ), .D(
        \ram[55][2] ), .S0(n6282), .S1(n6148), .Y(n4906) );
  MX4X1 U6569 ( .A(n4928), .B(n4926), .C(n4927), .D(n4925), .S0(n6036), .S1(
        n6058), .Y(n4929) );
  MX4X1 U6570 ( .A(\ram[240][3] ), .B(\ram[241][3] ), .C(\ram[242][3] ), .D(
        \ram[243][3] ), .S0(n6283), .S1(n6149), .Y(n4928) );
  MX4X1 U6571 ( .A(\ram[248][3] ), .B(\ram[249][3] ), .C(\ram[250][3] ), .D(
        \ram[251][3] ), .S0(n6283), .S1(n6149), .Y(n4926) );
  MX4X1 U6572 ( .A(\ram[244][3] ), .B(\ram[245][3] ), .C(\ram[246][3] ), .D(
        \ram[247][3] ), .S0(n6283), .S1(n6149), .Y(n4927) );
  MX4X1 U6573 ( .A(n4991), .B(n4989), .C(n4990), .D(n4988), .S0(n6037), .S1(
        n6059), .Y(n4992) );
  MX4X1 U6574 ( .A(\ram[48][3] ), .B(\ram[49][3] ), .C(\ram[50][3] ), .D(
        \ram[51][3] ), .S0(n6287), .S1(n6153), .Y(n4991) );
  MX4X1 U6575 ( .A(\ram[56][3] ), .B(\ram[57][3] ), .C(\ram[58][3] ), .D(
        \ram[59][3] ), .S0(n6287), .S1(n6153), .Y(n4989) );
  MX4X1 U6576 ( .A(\ram[52][3] ), .B(\ram[53][3] ), .C(\ram[54][3] ), .D(
        \ram[55][3] ), .S0(n6287), .S1(n6153), .Y(n4990) );
  MX4X1 U6577 ( .A(n4949), .B(n4947), .C(n4948), .D(n4946), .S0(n6040), .S1(
        n6059), .Y(n4950) );
  MX4X1 U6578 ( .A(\ram[176][3] ), .B(\ram[177][3] ), .C(\ram[178][3] ), .D(
        \ram[179][3] ), .S0(n6285), .S1(n6151), .Y(n4949) );
  MX4X1 U6579 ( .A(\ram[184][3] ), .B(\ram[185][3] ), .C(\ram[186][3] ), .D(
        \ram[187][3] ), .S0(n6285), .S1(n6151), .Y(n4947) );
  MX4X1 U6580 ( .A(\ram[180][3] ), .B(\ram[181][3] ), .C(\ram[182][3] ), .D(
        \ram[183][3] ), .S0(n6285), .S1(n6151), .Y(n4948) );
  MX4X1 U6581 ( .A(n5012), .B(n5010), .C(n5011), .D(n5009), .S0(n6034), .S1(
        n6060), .Y(n5013) );
  MX4X1 U6582 ( .A(\ram[240][4] ), .B(\ram[241][4] ), .C(\ram[242][4] ), .D(
        \ram[243][4] ), .S0(n6289), .S1(n6155), .Y(n5012) );
  MX4X1 U6583 ( .A(\ram[248][4] ), .B(\ram[249][4] ), .C(\ram[250][4] ), .D(
        \ram[251][4] ), .S0(n6289), .S1(n6155), .Y(n5010) );
  MX4X1 U6584 ( .A(\ram[244][4] ), .B(\ram[245][4] ), .C(\ram[246][4] ), .D(
        \ram[247][4] ), .S0(n6289), .S1(n6155), .Y(n5011) );
  MX4X1 U6585 ( .A(n5054), .B(n5052), .C(n5053), .D(n5051), .S0(n6034), .S1(
        n6060), .Y(n5055) );
  MX4X1 U6586 ( .A(\ram[112][4] ), .B(\ram[113][4] ), .C(\ram[114][4] ), .D(
        \ram[115][4] ), .S0(n6291), .S1(n6157), .Y(n5054) );
  MX4X1 U6587 ( .A(\ram[120][4] ), .B(\ram[121][4] ), .C(\ram[122][4] ), .D(
        \ram[123][4] ), .S0(n6291), .S1(n6157), .Y(n5052) );
  MX4X1 U6588 ( .A(\ram[116][4] ), .B(\ram[117][4] ), .C(\ram[118][4] ), .D(
        \ram[119][4] ), .S0(n6291), .S1(n6157), .Y(n5053) );
  MX4X1 U6589 ( .A(n5033), .B(n5031), .C(n5032), .D(n5030), .S0(n6034), .S1(
        n6060), .Y(n5034) );
  MX4X1 U6590 ( .A(\ram[176][4] ), .B(\ram[177][4] ), .C(\ram[178][4] ), .D(
        \ram[179][4] ), .S0(n6290), .S1(n6156), .Y(n5033) );
  MX4X1 U6591 ( .A(\ram[184][4] ), .B(\ram[185][4] ), .C(\ram[186][4] ), .D(
        \ram[187][4] ), .S0(n6290), .S1(n6156), .Y(n5031) );
  MX4X1 U6592 ( .A(\ram[180][4] ), .B(\ram[181][4] ), .C(\ram[182][4] ), .D(
        \ram[183][4] ), .S0(n6290), .S1(n6156), .Y(n5032) );
  MX4X1 U6593 ( .A(n5075), .B(n5073), .C(n5074), .D(n5072), .S0(n6038), .S1(
        n6061), .Y(n5076) );
  MX4X1 U6594 ( .A(\ram[48][4] ), .B(\ram[49][4] ), .C(\ram[50][4] ), .D(
        \ram[51][4] ), .S0(n6293), .S1(n6159), .Y(n5075) );
  MX4X1 U6595 ( .A(\ram[56][4] ), .B(\ram[57][4] ), .C(\ram[58][4] ), .D(
        \ram[59][4] ), .S0(n6293), .S1(n6159), .Y(n5073) );
  MX4X1 U6596 ( .A(\ram[52][4] ), .B(\ram[53][4] ), .C(\ram[54][4] ), .D(
        \ram[55][4] ), .S0(n6293), .S1(n6159), .Y(n5074) );
  MX4X1 U6597 ( .A(n5096), .B(n5094), .C(n5095), .D(n5093), .S0(n6044), .S1(
        n6061), .Y(n5097) );
  MX4X1 U6598 ( .A(\ram[240][5] ), .B(\ram[241][5] ), .C(\ram[242][5] ), .D(
        \ram[243][5] ), .S0(n6294), .S1(n6160), .Y(n5096) );
  MX4X1 U6599 ( .A(\ram[248][5] ), .B(\ram[249][5] ), .C(\ram[250][5] ), .D(
        \ram[251][5] ), .S0(n6294), .S1(n6160), .Y(n5094) );
  MX4X1 U6600 ( .A(\ram[244][5] ), .B(\ram[245][5] ), .C(\ram[246][5] ), .D(
        \ram[247][5] ), .S0(n6294), .S1(n6160), .Y(n5095) );
  MX4X1 U6601 ( .A(n5138), .B(n5136), .C(n5137), .D(n5135), .S0(n6035), .S1(
        n6062), .Y(n5139) );
  MX4X1 U6602 ( .A(\ram[112][5] ), .B(\ram[113][5] ), .C(\ram[114][5] ), .D(
        \ram[115][5] ), .S0(n6297), .S1(n6163), .Y(n5138) );
  MX4X1 U6603 ( .A(\ram[120][5] ), .B(\ram[121][5] ), .C(\ram[122][5] ), .D(
        \ram[123][5] ), .S0(n6297), .S1(n6163), .Y(n5136) );
  MX4X1 U6604 ( .A(\ram[116][5] ), .B(\ram[117][5] ), .C(\ram[118][5] ), .D(
        \ram[119][5] ), .S0(n6297), .S1(n6163), .Y(n5137) );
  MX4X1 U6605 ( .A(n5117), .B(n5115), .C(n5116), .D(n5114), .S0(n6041), .S1(
        n6061), .Y(n5118) );
  MX4X1 U6606 ( .A(\ram[176][5] ), .B(\ram[177][5] ), .C(\ram[178][5] ), .D(
        \ram[179][5] ), .S0(n6295), .S1(n6161), .Y(n5117) );
  MX4X1 U6607 ( .A(\ram[184][5] ), .B(\ram[185][5] ), .C(\ram[186][5] ), .D(
        \ram[187][5] ), .S0(n6295), .S1(n6161), .Y(n5115) );
  MX4X1 U6608 ( .A(\ram[180][5] ), .B(\ram[181][5] ), .C(\ram[182][5] ), .D(
        \ram[183][5] ), .S0(n6295), .S1(n6161), .Y(n5116) );
  MX4X1 U6609 ( .A(n5159), .B(n5157), .C(n5158), .D(n5156), .S0(n6035), .S1(
        n6062), .Y(n5160) );
  MX4X1 U6610 ( .A(\ram[48][5] ), .B(\ram[49][5] ), .C(\ram[50][5] ), .D(
        \ram[51][5] ), .S0(n6298), .S1(n6164), .Y(n5159) );
  MX4X1 U6611 ( .A(\ram[56][5] ), .B(\ram[57][5] ), .C(\ram[58][5] ), .D(
        \ram[59][5] ), .S0(n6298), .S1(n6164), .Y(n5157) );
  MX4X1 U6612 ( .A(\ram[52][5] ), .B(\ram[53][5] ), .C(\ram[54][5] ), .D(
        \ram[55][5] ), .S0(n6298), .S1(n6164), .Y(n5158) );
  MX4X1 U6613 ( .A(n5180), .B(n5178), .C(n5179), .D(n5177), .S0(n6035), .S1(
        n6062), .Y(n5181) );
  MX4X1 U6614 ( .A(\ram[240][6] ), .B(\ram[241][6] ), .C(\ram[242][6] ), .D(
        \ram[243][6] ), .S0(n6299), .S1(n6165), .Y(n5180) );
  MX4X1 U6615 ( .A(\ram[248][6] ), .B(\ram[249][6] ), .C(\ram[250][6] ), .D(
        \ram[251][6] ), .S0(n6299), .S1(n6165), .Y(n5178) );
  MX4X1 U6616 ( .A(\ram[244][6] ), .B(\ram[245][6] ), .C(\ram[246][6] ), .D(
        \ram[247][6] ), .S0(n6299), .S1(n6165), .Y(n5179) );
  MX4X1 U6617 ( .A(n5222), .B(n5220), .C(n5221), .D(n5219), .S0(n6046), .S1(
        n6063), .Y(n5223) );
  MX4X1 U6618 ( .A(\ram[112][6] ), .B(\ram[113][6] ), .C(\ram[114][6] ), .D(
        \ram[115][6] ), .S0(n6302), .S1(n6168), .Y(n5222) );
  MX4X1 U6619 ( .A(\ram[120][6] ), .B(\ram[121][6] ), .C(\ram[122][6] ), .D(
        \ram[123][6] ), .S0(n6302), .S1(n6168), .Y(n5220) );
  MX4X1 U6620 ( .A(\ram[116][6] ), .B(\ram[117][6] ), .C(\ram[118][6] ), .D(
        \ram[119][6] ), .S0(n6302), .S1(n6168), .Y(n5221) );
  MX4X1 U6621 ( .A(n5201), .B(n5199), .C(n5200), .D(n5198), .S0(n6042), .S1(
        n6063), .Y(n5202) );
  MX4X1 U6622 ( .A(\ram[176][6] ), .B(\ram[177][6] ), .C(\ram[178][6] ), .D(
        \ram[179][6] ), .S0(n6301), .S1(n6167), .Y(n5201) );
  MX4X1 U6623 ( .A(\ram[184][6] ), .B(\ram[185][6] ), .C(\ram[186][6] ), .D(
        \ram[187][6] ), .S0(n6301), .S1(n6167), .Y(n5199) );
  MX4X1 U6624 ( .A(\ram[180][6] ), .B(\ram[181][6] ), .C(\ram[182][6] ), .D(
        \ram[183][6] ), .S0(n6301), .S1(n6167), .Y(n5200) );
  MX4X1 U6625 ( .A(n5243), .B(n5241), .C(n5242), .D(n5240), .S0(n6037), .S1(
        n6063), .Y(n5244) );
  MX4X1 U6626 ( .A(\ram[48][6] ), .B(\ram[49][6] ), .C(\ram[50][6] ), .D(
        \ram[51][6] ), .S0(n6303), .S1(n6169), .Y(n5243) );
  MX4X1 U6627 ( .A(\ram[56][6] ), .B(\ram[57][6] ), .C(\ram[58][6] ), .D(
        \ram[59][6] ), .S0(n6303), .S1(n6169), .Y(n5241) );
  MX4X1 U6628 ( .A(\ram[52][6] ), .B(\ram[53][6] ), .C(\ram[54][6] ), .D(
        \ram[55][6] ), .S0(n6303), .S1(n6169), .Y(n5242) );
  MX4X1 U6629 ( .A(n5264), .B(n5262), .C(n5263), .D(n5261), .S0(n6036), .S1(
        n6064), .Y(n5265) );
  MX4X1 U6630 ( .A(\ram[240][7] ), .B(\ram[241][7] ), .C(\ram[242][7] ), .D(
        \ram[243][7] ), .S0(n6305), .S1(n6171), .Y(n5264) );
  MX4X1 U6631 ( .A(\ram[248][7] ), .B(\ram[249][7] ), .C(\ram[250][7] ), .D(
        \ram[251][7] ), .S0(n6305), .S1(n6171), .Y(n5262) );
  MX4X1 U6632 ( .A(\ram[244][7] ), .B(\ram[245][7] ), .C(\ram[246][7] ), .D(
        \ram[247][7] ), .S0(n6305), .S1(n6171), .Y(n5263) );
  MX4X1 U6633 ( .A(n5306), .B(n5304), .C(n5305), .D(n5303), .S0(n6036), .S1(
        n6064), .Y(n5307) );
  MX4X1 U6634 ( .A(\ram[112][7] ), .B(\ram[113][7] ), .C(\ram[114][7] ), .D(
        \ram[115][7] ), .S0(n6307), .S1(n6173), .Y(n5306) );
  MX4X1 U6635 ( .A(\ram[120][7] ), .B(\ram[121][7] ), .C(\ram[122][7] ), .D(
        \ram[123][7] ), .S0(n6307), .S1(n6173), .Y(n5304) );
  MX4X1 U6636 ( .A(\ram[116][7] ), .B(\ram[117][7] ), .C(\ram[118][7] ), .D(
        \ram[119][7] ), .S0(n6307), .S1(n6173), .Y(n5305) );
  MX4X1 U6637 ( .A(n5285), .B(n5283), .C(n5284), .D(n5282), .S0(n6036), .S1(
        n6064), .Y(n5286) );
  MX4X1 U6638 ( .A(\ram[176][7] ), .B(\ram[177][7] ), .C(\ram[178][7] ), .D(
        \ram[179][7] ), .S0(n6306), .S1(n6172), .Y(n5285) );
  MX4X1 U6639 ( .A(\ram[184][7] ), .B(\ram[185][7] ), .C(\ram[186][7] ), .D(
        \ram[187][7] ), .S0(n6306), .S1(n6172), .Y(n5283) );
  MX4X1 U6640 ( .A(\ram[180][7] ), .B(\ram[181][7] ), .C(\ram[182][7] ), .D(
        \ram[183][7] ), .S0(n6306), .S1(n6172), .Y(n5284) );
  MX4X1 U6641 ( .A(n5327), .B(n5325), .C(n5326), .D(n5324), .S0(n6037), .S1(
        n6065), .Y(n5328) );
  MX4X1 U6642 ( .A(\ram[48][7] ), .B(\ram[49][7] ), .C(\ram[50][7] ), .D(
        \ram[51][7] ), .S0(n6309), .S1(n6175), .Y(n5327) );
  MX4X1 U6643 ( .A(\ram[56][7] ), .B(\ram[57][7] ), .C(\ram[58][7] ), .D(
        \ram[59][7] ), .S0(n6309), .S1(n6175), .Y(n5325) );
  MX4X1 U6644 ( .A(\ram[52][7] ), .B(\ram[53][7] ), .C(\ram[54][7] ), .D(
        \ram[55][7] ), .S0(n6309), .S1(n6175), .Y(n5326) );
  MX4X1 U6645 ( .A(n5348), .B(n5346), .C(n5347), .D(n5345), .S0(n6037), .S1(
        n6065), .Y(n5349) );
  MX4X1 U6646 ( .A(\ram[240][8] ), .B(\ram[241][8] ), .C(\ram[242][8] ), .D(
        \ram[243][8] ), .S0(n6310), .S1(n6176), .Y(n5348) );
  MX4X1 U6647 ( .A(\ram[248][8] ), .B(\ram[249][8] ), .C(\ram[250][8] ), .D(
        \ram[251][8] ), .S0(n6310), .S1(n6176), .Y(n5346) );
  MX4X1 U6648 ( .A(\ram[244][8] ), .B(\ram[245][8] ), .C(\ram[246][8] ), .D(
        \ram[247][8] ), .S0(n6310), .S1(n6176), .Y(n5347) );
  MX4X1 U6649 ( .A(n5390), .B(n5388), .C(n5389), .D(n5387), .S0(n6038), .S1(
        n6066), .Y(n5391) );
  MX4X1 U6650 ( .A(\ram[112][8] ), .B(\ram[113][8] ), .C(\ram[114][8] ), .D(
        \ram[115][8] ), .S0(n6313), .S1(n6179), .Y(n5390) );
  MX4X1 U6651 ( .A(\ram[120][8] ), .B(\ram[121][8] ), .C(\ram[122][8] ), .D(
        \ram[123][8] ), .S0(n6313), .S1(n6179), .Y(n5388) );
  MX4X1 U6652 ( .A(\ram[116][8] ), .B(\ram[117][8] ), .C(\ram[118][8] ), .D(
        \ram[119][8] ), .S0(n6313), .S1(n6179), .Y(n5389) );
  MX4X1 U6653 ( .A(n5369), .B(n5367), .C(n5368), .D(n5366), .S0(n6037), .S1(
        n6065), .Y(n5370) );
  MX4X1 U6654 ( .A(\ram[176][8] ), .B(\ram[177][8] ), .C(\ram[178][8] ), .D(
        \ram[179][8] ), .S0(n6311), .S1(n6177), .Y(n5369) );
  MX4X1 U6655 ( .A(\ram[184][8] ), .B(\ram[185][8] ), .C(\ram[186][8] ), .D(
        \ram[187][8] ), .S0(n6311), .S1(n6177), .Y(n5367) );
  MX4X1 U6656 ( .A(\ram[180][8] ), .B(\ram[181][8] ), .C(\ram[182][8] ), .D(
        \ram[183][8] ), .S0(n6311), .S1(n6177), .Y(n5368) );
  MX4X1 U6657 ( .A(n5411), .B(n5409), .C(n5410), .D(n5408), .S0(n6038), .S1(
        n6066), .Y(n5412) );
  MX4X1 U6658 ( .A(\ram[48][8] ), .B(\ram[49][8] ), .C(\ram[50][8] ), .D(
        \ram[51][8] ), .S0(n6314), .S1(n6180), .Y(n5411) );
  MX4X1 U6659 ( .A(\ram[56][8] ), .B(\ram[57][8] ), .C(\ram[58][8] ), .D(
        \ram[59][8] ), .S0(n6314), .S1(n6180), .Y(n5409) );
  MX4X1 U6660 ( .A(\ram[52][8] ), .B(\ram[53][8] ), .C(\ram[54][8] ), .D(
        \ram[55][8] ), .S0(n6314), .S1(n6180), .Y(n5410) );
  MX4X1 U6661 ( .A(n5432), .B(n5430), .C(n5431), .D(n5429), .S0(n6038), .S1(
        n6066), .Y(n5433) );
  MX4X1 U6662 ( .A(\ram[240][9] ), .B(\ram[241][9] ), .C(\ram[242][9] ), .D(
        \ram[243][9] ), .S0(n6315), .S1(n6181), .Y(n5432) );
  MX4X1 U6663 ( .A(\ram[248][9] ), .B(\ram[249][9] ), .C(\ram[250][9] ), .D(
        \ram[251][9] ), .S0(n6315), .S1(n6181), .Y(n5430) );
  MX4X1 U6664 ( .A(\ram[244][9] ), .B(\ram[245][9] ), .C(\ram[246][9] ), .D(
        \ram[247][9] ), .S0(n6315), .S1(n6181), .Y(n5431) );
  MX4X1 U6665 ( .A(n5474), .B(n5472), .C(n5473), .D(n5471), .S0(n6039), .S1(
        n6067), .Y(n5475) );
  MX4X1 U6666 ( .A(\ram[112][9] ), .B(\ram[113][9] ), .C(\ram[114][9] ), .D(
        \ram[115][9] ), .S0(n6318), .S1(n6184), .Y(n5474) );
  MX4X1 U6667 ( .A(\ram[120][9] ), .B(\ram[121][9] ), .C(\ram[122][9] ), .D(
        \ram[123][9] ), .S0(n6318), .S1(n6184), .Y(n5472) );
  MX4X1 U6668 ( .A(\ram[116][9] ), .B(\ram[117][9] ), .C(\ram[118][9] ), .D(
        \ram[119][9] ), .S0(n6318), .S1(n6184), .Y(n5473) );
  MX4X1 U6669 ( .A(n5453), .B(n5451), .C(n5452), .D(n5450), .S0(n6039), .S1(
        n6067), .Y(n5454) );
  MX4X1 U6670 ( .A(\ram[176][9] ), .B(\ram[177][9] ), .C(\ram[178][9] ), .D(
        \ram[179][9] ), .S0(n6317), .S1(n6183), .Y(n5453) );
  MX4X1 U6671 ( .A(\ram[184][9] ), .B(\ram[185][9] ), .C(\ram[186][9] ), .D(
        \ram[187][9] ), .S0(n6317), .S1(n6183), .Y(n5451) );
  MX4X1 U6672 ( .A(\ram[180][9] ), .B(\ram[181][9] ), .C(\ram[182][9] ), .D(
        \ram[183][9] ), .S0(n6317), .S1(n6183), .Y(n5452) );
  MX4X1 U6673 ( .A(n5495), .B(n5493), .C(n5494), .D(n5492), .S0(n6039), .S1(
        n6067), .Y(n5496) );
  MX4X1 U6674 ( .A(\ram[48][9] ), .B(\ram[49][9] ), .C(\ram[50][9] ), .D(
        \ram[51][9] ), .S0(n6319), .S1(n6185), .Y(n5495) );
  MX4X1 U6675 ( .A(\ram[56][9] ), .B(\ram[57][9] ), .C(\ram[58][9] ), .D(
        \ram[59][9] ), .S0(n6319), .S1(n6185), .Y(n5493) );
  MX4X1 U6676 ( .A(\ram[52][9] ), .B(\ram[53][9] ), .C(\ram[54][9] ), .D(
        \ram[55][9] ), .S0(n6319), .S1(n6185), .Y(n5494) );
  MX4X1 U6677 ( .A(n5516), .B(n5514), .C(n5515), .D(n5513), .S0(n6040), .S1(
        n6068), .Y(n5517) );
  MX4X1 U6678 ( .A(\ram[240][10] ), .B(\ram[241][10] ), .C(\ram[242][10] ), 
        .D(\ram[243][10] ), .S0(n6321), .S1(n6187), .Y(n5516) );
  MX4X1 U6679 ( .A(\ram[248][10] ), .B(\ram[249][10] ), .C(\ram[250][10] ), 
        .D(\ram[251][10] ), .S0(n6321), .S1(n6187), .Y(n5514) );
  MX4X1 U6680 ( .A(\ram[244][10] ), .B(\ram[245][10] ), .C(\ram[246][10] ), 
        .D(\ram[247][10] ), .S0(n6321), .S1(n6187), .Y(n5515) );
  MX4X1 U6681 ( .A(n5537), .B(n5535), .C(n5536), .D(n5534), .S0(n6040), .S1(
        n6068), .Y(n5538) );
  MX4X1 U6682 ( .A(\ram[176][10] ), .B(\ram[177][10] ), .C(\ram[178][10] ), 
        .D(\ram[179][10] ), .S0(n6322), .S1(n6188), .Y(n5537) );
  MX4X1 U6683 ( .A(\ram[184][10] ), .B(\ram[185][10] ), .C(\ram[186][10] ), 
        .D(\ram[187][10] ), .S0(n6322), .S1(n6188), .Y(n5535) );
  MX4X1 U6684 ( .A(\ram[180][10] ), .B(\ram[181][10] ), .C(\ram[182][10] ), 
        .D(\ram[183][10] ), .S0(n6322), .S1(n6188), .Y(n5536) );
  MX4X1 U6685 ( .A(n5558), .B(n5556), .C(n5557), .D(n5555), .S0(n6040), .S1(
        n6068), .Y(n5559) );
  MX4X1 U6686 ( .A(\ram[112][10] ), .B(\ram[113][10] ), .C(\ram[114][10] ), 
        .D(\ram[115][10] ), .S0(n6323), .S1(n6189), .Y(n5558) );
  MX4X1 U6687 ( .A(\ram[120][10] ), .B(\ram[121][10] ), .C(\ram[122][10] ), 
        .D(\ram[123][10] ), .S0(n6323), .S1(n6189), .Y(n5556) );
  MX4X1 U6688 ( .A(\ram[116][10] ), .B(\ram[117][10] ), .C(\ram[118][10] ), 
        .D(\ram[119][10] ), .S0(n6323), .S1(n6189), .Y(n5557) );
  MX4X1 U6689 ( .A(n5579), .B(n5577), .C(n5578), .D(n5576), .S0(n6041), .S1(
        n6069), .Y(n5580) );
  MX4X1 U6690 ( .A(\ram[48][10] ), .B(\ram[49][10] ), .C(\ram[50][10] ), .D(
        \ram[51][10] ), .S0(n6325), .S1(n6191), .Y(n5579) );
  MX4X1 U6691 ( .A(\ram[56][10] ), .B(\ram[57][10] ), .C(\ram[58][10] ), .D(
        \ram[59][10] ), .S0(n6325), .S1(n6191), .Y(n5577) );
  MX4X1 U6692 ( .A(\ram[52][10] ), .B(\ram[53][10] ), .C(\ram[54][10] ), .D(
        \ram[55][10] ), .S0(n6325), .S1(n6191), .Y(n5578) );
  MX4X1 U6693 ( .A(n5600), .B(n5598), .C(n5599), .D(n5597), .S0(n6041), .S1(
        n6069), .Y(n5601) );
  MX4X1 U6694 ( .A(\ram[240][11] ), .B(\ram[241][11] ), .C(\ram[242][11] ), 
        .D(\ram[243][11] ), .S0(n6326), .S1(n6192), .Y(n5600) );
  MX4X1 U6695 ( .A(\ram[248][11] ), .B(\ram[249][11] ), .C(\ram[250][11] ), 
        .D(\ram[251][11] ), .S0(n6326), .S1(n6192), .Y(n5598) );
  MX4X1 U6696 ( .A(\ram[244][11] ), .B(\ram[245][11] ), .C(\ram[246][11] ), 
        .D(\ram[247][11] ), .S0(n6326), .S1(n6192), .Y(n5599) );
  MX4X1 U6697 ( .A(n5642), .B(n5640), .C(n5641), .D(n5639), .S0(n6042), .S1(
        n6070), .Y(n5643) );
  MX4X1 U6698 ( .A(\ram[112][11] ), .B(\ram[113][11] ), .C(\ram[114][11] ), 
        .D(\ram[115][11] ), .S0(n6329), .S1(n6195), .Y(n5642) );
  MX4X1 U6699 ( .A(\ram[120][11] ), .B(\ram[121][11] ), .C(\ram[122][11] ), 
        .D(\ram[123][11] ), .S0(n6329), .S1(n6195), .Y(n5640) );
  MX4X1 U6700 ( .A(\ram[116][11] ), .B(\ram[117][11] ), .C(\ram[118][11] ), 
        .D(\ram[119][11] ), .S0(n6329), .S1(n6195), .Y(n5641) );
  MX4X1 U6701 ( .A(n5621), .B(n5619), .C(n5620), .D(n5618), .S0(n6041), .S1(
        n6069), .Y(n5622) );
  MX4X1 U6702 ( .A(\ram[176][11] ), .B(\ram[177][11] ), .C(\ram[178][11] ), 
        .D(\ram[179][11] ), .S0(n6327), .S1(n6193), .Y(n5621) );
  MX4X1 U6703 ( .A(\ram[184][11] ), .B(\ram[185][11] ), .C(\ram[186][11] ), 
        .D(\ram[187][11] ), .S0(n6327), .S1(n6193), .Y(n5619) );
  MX4X1 U6704 ( .A(\ram[180][11] ), .B(\ram[181][11] ), .C(\ram[182][11] ), 
        .D(\ram[183][11] ), .S0(n6327), .S1(n6193), .Y(n5620) );
  MX4X1 U6705 ( .A(n5663), .B(n5661), .C(n5662), .D(n5660), .S0(n6042), .S1(
        n6070), .Y(n5664) );
  MX4X1 U6706 ( .A(\ram[48][11] ), .B(\ram[49][11] ), .C(\ram[50][11] ), .D(
        \ram[51][11] ), .S0(n6330), .S1(n6196), .Y(n5663) );
  MX4X1 U6707 ( .A(\ram[56][11] ), .B(\ram[57][11] ), .C(\ram[58][11] ), .D(
        \ram[59][11] ), .S0(n6330), .S1(n6196), .Y(n5661) );
  MX4X1 U6708 ( .A(\ram[52][11] ), .B(\ram[53][11] ), .C(\ram[54][11] ), .D(
        \ram[55][11] ), .S0(n6330), .S1(n6196), .Y(n5662) );
  MX4X1 U6709 ( .A(n5684), .B(n5682), .C(n5683), .D(n5681), .S0(n6042), .S1(
        n6070), .Y(n5685) );
  MX4X1 U6710 ( .A(\ram[240][12] ), .B(\ram[241][12] ), .C(\ram[242][12] ), 
        .D(\ram[243][12] ), .S0(n6331), .S1(n6197), .Y(n5684) );
  MX4X1 U6711 ( .A(\ram[248][12] ), .B(\ram[249][12] ), .C(\ram[250][12] ), 
        .D(\ram[251][12] ), .S0(n6331), .S1(n6197), .Y(n5682) );
  MX4X1 U6712 ( .A(\ram[244][12] ), .B(\ram[245][12] ), .C(\ram[246][12] ), 
        .D(\ram[247][12] ), .S0(n6331), .S1(n6197), .Y(n5683) );
  MX4X1 U6713 ( .A(n5726), .B(n5724), .C(n5725), .D(n5723), .S0(n6043), .S1(
        n6071), .Y(n5727) );
  MX4X1 U6714 ( .A(\ram[112][12] ), .B(\ram[113][12] ), .C(\ram[114][12] ), 
        .D(\ram[115][12] ), .S0(n6334), .S1(n6200), .Y(n5726) );
  MX4X1 U6715 ( .A(\ram[120][12] ), .B(\ram[121][12] ), .C(\ram[122][12] ), 
        .D(\ram[123][12] ), .S0(n6334), .S1(n6200), .Y(n5724) );
  MX4X1 U6716 ( .A(\ram[116][12] ), .B(\ram[117][12] ), .C(\ram[118][12] ), 
        .D(\ram[119][12] ), .S0(n6334), .S1(n6200), .Y(n5725) );
  MX4X1 U6717 ( .A(n5705), .B(n5703), .C(n5704), .D(n5702), .S0(n6043), .S1(
        n6071), .Y(n5706) );
  MX4X1 U6718 ( .A(\ram[176][12] ), .B(\ram[177][12] ), .C(\ram[178][12] ), 
        .D(\ram[179][12] ), .S0(n6333), .S1(n6199), .Y(n5705) );
  MX4X1 U6719 ( .A(\ram[184][12] ), .B(\ram[185][12] ), .C(\ram[186][12] ), 
        .D(\ram[187][12] ), .S0(n6333), .S1(n6199), .Y(n5703) );
  MX4X1 U6720 ( .A(\ram[180][12] ), .B(\ram[181][12] ), .C(\ram[182][12] ), 
        .D(\ram[183][12] ), .S0(n6333), .S1(n6199), .Y(n5704) );
  MX4X1 U6721 ( .A(n5747), .B(n5745), .C(n5746), .D(n5744), .S0(n6043), .S1(
        n6071), .Y(n5748) );
  MX4X1 U6722 ( .A(\ram[48][12] ), .B(\ram[49][12] ), .C(\ram[50][12] ), .D(
        \ram[51][12] ), .S0(n6335), .S1(n6201), .Y(n5747) );
  MX4X1 U6723 ( .A(\ram[56][12] ), .B(\ram[57][12] ), .C(\ram[58][12] ), .D(
        \ram[59][12] ), .S0(n6335), .S1(n6201), .Y(n5745) );
  MX4X1 U6724 ( .A(\ram[52][12] ), .B(\ram[53][12] ), .C(\ram[54][12] ), .D(
        \ram[55][12] ), .S0(n6335), .S1(n6201), .Y(n5746) );
  MX4X1 U6725 ( .A(n5768), .B(n5766), .C(n5767), .D(n5765), .S0(n6044), .S1(
        n6072), .Y(n5769) );
  MX4X1 U6726 ( .A(\ram[240][13] ), .B(\ram[241][13] ), .C(\ram[242][13] ), 
        .D(\ram[243][13] ), .S0(n6337), .S1(n6203), .Y(n5768) );
  MX4X1 U6727 ( .A(\ram[248][13] ), .B(\ram[249][13] ), .C(\ram[250][13] ), 
        .D(\ram[251][13] ), .S0(n6337), .S1(n6203), .Y(n5766) );
  MX4X1 U6728 ( .A(\ram[244][13] ), .B(\ram[245][13] ), .C(\ram[246][13] ), 
        .D(\ram[247][13] ), .S0(n6337), .S1(n6203), .Y(n5767) );
  MX4X1 U6729 ( .A(n5810), .B(n5808), .C(n5809), .D(n5807), .S0(n6044), .S1(
        n6072), .Y(n5811) );
  MX4X1 U6730 ( .A(\ram[112][13] ), .B(\ram[113][13] ), .C(\ram[114][13] ), 
        .D(\ram[115][13] ), .S0(n6339), .S1(n6205), .Y(n5810) );
  MX4X1 U6731 ( .A(\ram[120][13] ), .B(\ram[121][13] ), .C(\ram[122][13] ), 
        .D(\ram[123][13] ), .S0(n6339), .S1(n6205), .Y(n5808) );
  MX4X1 U6732 ( .A(\ram[116][13] ), .B(\ram[117][13] ), .C(\ram[118][13] ), 
        .D(\ram[119][13] ), .S0(n6339), .S1(n6205), .Y(n5809) );
  MX4X1 U6733 ( .A(n5789), .B(n5787), .C(n5788), .D(n5786), .S0(n6044), .S1(
        n6072), .Y(n5790) );
  MX4X1 U6734 ( .A(\ram[176][13] ), .B(\ram[177][13] ), .C(\ram[178][13] ), 
        .D(\ram[179][13] ), .S0(n6338), .S1(n6204), .Y(n5789) );
  MX4X1 U6735 ( .A(\ram[184][13] ), .B(\ram[185][13] ), .C(\ram[186][13] ), 
        .D(\ram[187][13] ), .S0(n6338), .S1(n6204), .Y(n5787) );
  MX4X1 U6736 ( .A(\ram[180][13] ), .B(\ram[181][13] ), .C(\ram[182][13] ), 
        .D(\ram[183][13] ), .S0(n6338), .S1(n6204), .Y(n5788) );
  MX4X1 U6737 ( .A(n5831), .B(n5829), .C(n5830), .D(n5828), .S0(n6045), .S1(
        n6073), .Y(n5832) );
  MX4X1 U6738 ( .A(\ram[48][13] ), .B(\ram[49][13] ), .C(\ram[50][13] ), .D(
        \ram[51][13] ), .S0(n6341), .S1(n6207), .Y(n5831) );
  MX4X1 U6739 ( .A(\ram[56][13] ), .B(\ram[57][13] ), .C(\ram[58][13] ), .D(
        \ram[59][13] ), .S0(n6341), .S1(n6207), .Y(n5829) );
  MX4X1 U6740 ( .A(\ram[52][13] ), .B(\ram[53][13] ), .C(\ram[54][13] ), .D(
        \ram[55][13] ), .S0(n6341), .S1(n6207), .Y(n5830) );
  MX4X1 U6741 ( .A(n5852), .B(n5850), .C(n5851), .D(n5849), .S0(n6045), .S1(
        n6073), .Y(n5853) );
  MX4X1 U6742 ( .A(\ram[240][14] ), .B(\ram[241][14] ), .C(\ram[242][14] ), 
        .D(\ram[243][14] ), .S0(n6342), .S1(n6208), .Y(n5852) );
  MX4X1 U6743 ( .A(\ram[248][14] ), .B(\ram[249][14] ), .C(\ram[250][14] ), 
        .D(\ram[251][14] ), .S0(n6342), .S1(n6208), .Y(n5850) );
  MX4X1 U6744 ( .A(\ram[244][14] ), .B(\ram[245][14] ), .C(\ram[246][14] ), 
        .D(\ram[247][14] ), .S0(n6342), .S1(n6208), .Y(n5851) );
  MX4X1 U6745 ( .A(n5894), .B(n5892), .C(n5893), .D(n5891), .S0(n6046), .S1(
        n6060), .Y(n5895) );
  MX4X1 U6746 ( .A(\ram[112][14] ), .B(\ram[113][14] ), .C(\ram[114][14] ), 
        .D(\ram[115][14] ), .S0(n6345), .S1(n6211), .Y(n5894) );
  MX4X1 U6747 ( .A(\ram[120][14] ), .B(\ram[121][14] ), .C(\ram[122][14] ), 
        .D(\ram[123][14] ), .S0(n6345), .S1(n6211), .Y(n5892) );
  MX4X1 U6748 ( .A(\ram[116][14] ), .B(\ram[117][14] ), .C(\ram[118][14] ), 
        .D(\ram[119][14] ), .S0(n6345), .S1(n6211), .Y(n5893) );
  MX4X1 U6749 ( .A(n5873), .B(n5871), .C(n5872), .D(n5870), .S0(n6045), .S1(
        n6073), .Y(n5874) );
  MX4X1 U6750 ( .A(\ram[176][14] ), .B(\ram[177][14] ), .C(\ram[178][14] ), 
        .D(\ram[179][14] ), .S0(n6343), .S1(n6209), .Y(n5873) );
  MX4X1 U6751 ( .A(\ram[184][14] ), .B(\ram[185][14] ), .C(\ram[186][14] ), 
        .D(\ram[187][14] ), .S0(n6343), .S1(n6209), .Y(n5871) );
  MX4X1 U6752 ( .A(\ram[180][14] ), .B(\ram[181][14] ), .C(\ram[182][14] ), 
        .D(\ram[183][14] ), .S0(n6343), .S1(n6209), .Y(n5872) );
  MX4X1 U6753 ( .A(n5915), .B(n5913), .C(n5914), .D(n5912), .S0(n6046), .S1(
        n6073), .Y(n5916) );
  MX4X1 U6754 ( .A(\ram[48][14] ), .B(\ram[49][14] ), .C(\ram[50][14] ), .D(
        \ram[51][14] ), .S0(n6346), .S1(n6212), .Y(n5915) );
  MX4X1 U6755 ( .A(\ram[56][14] ), .B(\ram[57][14] ), .C(\ram[58][14] ), .D(
        \ram[59][14] ), .S0(n6346), .S1(n6212), .Y(n5913) );
  MX4X1 U6756 ( .A(\ram[52][14] ), .B(\ram[53][14] ), .C(\ram[54][14] ), .D(
        \ram[55][14] ), .S0(n6346), .S1(n6212), .Y(n5914) );
  MX4X1 U6757 ( .A(n5936), .B(n5934), .C(n5935), .D(n5933), .S0(n6046), .S1(
        n6073), .Y(n5937) );
  MX4X1 U6758 ( .A(\ram[240][15] ), .B(\ram[241][15] ), .C(\ram[242][15] ), 
        .D(\ram[243][15] ), .S0(n6347), .S1(n6214), .Y(n5936) );
  MX4X1 U6759 ( .A(\ram[248][15] ), .B(\ram[249][15] ), .C(\ram[250][15] ), 
        .D(\ram[251][15] ), .S0(n6347), .S1(n6189), .Y(n5934) );
  MX4X1 U6760 ( .A(\ram[244][15] ), .B(\ram[245][15] ), .C(\ram[246][15] ), 
        .D(\ram[247][15] ), .S0(n6347), .S1(n6093), .Y(n5935) );
  MX4X1 U6761 ( .A(n5978), .B(n5976), .C(n5977), .D(n5975), .S0(n6047), .S1(
        n6063), .Y(n5979) );
  MX4X1 U6762 ( .A(\ram[112][15] ), .B(\ram[113][15] ), .C(\ram[114][15] ), 
        .D(\ram[115][15] ), .S0(n6350), .S1(n6214), .Y(n5978) );
  MX4X1 U6763 ( .A(\ram[120][15] ), .B(\ram[121][15] ), .C(\ram[122][15] ), 
        .D(\ram[123][15] ), .S0(n6350), .S1(n6213), .Y(n5976) );
  MX4X1 U6764 ( .A(\ram[116][15] ), .B(\ram[117][15] ), .C(\ram[118][15] ), 
        .D(\ram[119][15] ), .S0(n6350), .S1(n6139), .Y(n5977) );
  MX4X1 U6765 ( .A(n5957), .B(n5955), .C(n5956), .D(n5954), .S0(n6047), .S1(
        n6063), .Y(n5958) );
  MX4X1 U6766 ( .A(\ram[176][15] ), .B(\ram[177][15] ), .C(\ram[178][15] ), 
        .D(\ram[179][15] ), .S0(n6349), .S1(n6214), .Y(n5957) );
  MX4X1 U6767 ( .A(\ram[184][15] ), .B(\ram[185][15] ), .C(\ram[186][15] ), 
        .D(\ram[187][15] ), .S0(n6349), .S1(n6214), .Y(n5955) );
  MX4X1 U6768 ( .A(\ram[180][15] ), .B(\ram[181][15] ), .C(\ram[182][15] ), 
        .D(\ram[183][15] ), .S0(n6349), .S1(n6214), .Y(n5956) );
  MX4X1 U6769 ( .A(n5999), .B(n5997), .C(n5998), .D(n5996), .S0(n6047), .S1(
        n6060), .Y(n6000) );
  MX4X1 U6770 ( .A(\ram[48][15] ), .B(\ram[49][15] ), .C(\ram[50][15] ), .D(
        \ram[51][15] ), .S0(n6351), .S1(n6090), .Y(n5999) );
  MX4X1 U6771 ( .A(\ram[56][15] ), .B(\ram[57][15] ), .C(\ram[58][15] ), .D(
        \ram[59][15] ), .S0(n6351), .S1(n6193), .Y(n5997) );
  MX4X1 U6772 ( .A(\ram[52][15] ), .B(\ram[53][15] ), .C(\ram[54][15] ), .D(
        \ram[55][15] ), .S0(n6351), .S1(n6194), .Y(n5998) );
  MX4X1 U6773 ( .A(\ram[88][0] ), .B(\ram[89][0] ), .C(\ram[90][0] ), .D(
        \ram[91][0] ), .S0(n6271), .S1(n6137), .Y(n4726) );
  MX4X1 U6774 ( .A(\ram[104][0] ), .B(\ram[105][0] ), .C(\ram[106][0] ), .D(
        \ram[107][0] ), .S0(n6270), .S1(n6136), .Y(n4721) );
  MX4X1 U6775 ( .A(\ram[72][0] ), .B(\ram[73][0] ), .C(\ram[74][0] ), .D(
        \ram[75][0] ), .S0(n6271), .S1(n6137), .Y(n4731) );
  MX4X1 U6776 ( .A(\ram[216][1] ), .B(\ram[217][1] ), .C(\ram[218][1] ), .D(
        \ram[219][1] ), .S0(n6273), .S1(n6139), .Y(n4768) );
  MX4X1 U6777 ( .A(\ram[232][1] ), .B(\ram[233][1] ), .C(\ram[234][1] ), .D(
        \ram[235][1] ), .S0(n6273), .S1(n6139), .Y(n4763) );
  MX4X1 U6778 ( .A(\ram[200][1] ), .B(\ram[201][1] ), .C(\ram[202][1] ), .D(
        \ram[203][1] ), .S0(n6274), .S1(n6140), .Y(n4773) );
  MX4X1 U6779 ( .A(\ram[216][2] ), .B(\ram[217][2] ), .C(\ram[218][2] ), .D(
        \ram[219][2] ), .S0(n6279), .S1(n6145), .Y(n4852) );
  MX4X1 U6780 ( .A(\ram[232][2] ), .B(\ram[233][2] ), .C(\ram[234][2] ), .D(
        \ram[235][2] ), .S0(n6278), .S1(n6144), .Y(n4847) );
  MX4X1 U6781 ( .A(\ram[200][2] ), .B(\ram[201][2] ), .C(\ram[202][2] ), .D(
        \ram[203][2] ), .S0(n6279), .S1(n6145), .Y(n4857) );
  MX4X1 U6782 ( .A(\ram[120][3] ), .B(\ram[121][3] ), .C(\ram[122][3] ), .D(
        \ram[123][3] ), .S0(n6286), .S1(n6152), .Y(n4968) );
  MX4X1 U6783 ( .A(\ram[72][3] ), .B(\ram[73][3] ), .C(\ram[74][3] ), .D(
        \ram[75][3] ), .S0(n6287), .S1(n6153), .Y(n4983) );
  MX4X1 U6784 ( .A(\ram[104][3] ), .B(\ram[105][3] ), .C(\ram[106][3] ), .D(
        \ram[107][3] ), .S0(n6286), .S1(n6152), .Y(n4973) );
  MX4X1 U6785 ( .A(\ram[216][4] ), .B(\ram[217][4] ), .C(\ram[218][4] ), .D(
        \ram[219][4] ), .S0(n6289), .S1(n6155), .Y(n5020) );
  MX4X1 U6786 ( .A(\ram[232][4] ), .B(\ram[233][4] ), .C(\ram[234][4] ), .D(
        \ram[235][4] ), .S0(n6289), .S1(n6155), .Y(n5015) );
  MX4X1 U6787 ( .A(\ram[200][4] ), .B(\ram[201][4] ), .C(\ram[202][4] ), .D(
        \ram[203][4] ), .S0(n6290), .S1(n6156), .Y(n5025) );
  MX4X1 U6788 ( .A(\ram[216][5] ), .B(\ram[217][5] ), .C(\ram[218][5] ), .D(
        \ram[219][5] ), .S0(n6295), .S1(n6161), .Y(n5104) );
  MX4X1 U6789 ( .A(\ram[232][5] ), .B(\ram[233][5] ), .C(\ram[234][5] ), .D(
        \ram[235][5] ), .S0(n6294), .S1(n6160), .Y(n5099) );
  MX4X1 U6790 ( .A(\ram[200][5] ), .B(\ram[201][5] ), .C(\ram[202][5] ), .D(
        \ram[203][5] ), .S0(n6295), .S1(n6161), .Y(n5109) );
  MX4X1 U6791 ( .A(\ram[216][6] ), .B(\ram[217][6] ), .C(\ram[218][6] ), .D(
        \ram[219][6] ), .S0(n6300), .S1(n6166), .Y(n5188) );
  MX4X1 U6792 ( .A(\ram[232][6] ), .B(\ram[233][6] ), .C(\ram[234][6] ), .D(
        \ram[235][6] ), .S0(n6300), .S1(n6166), .Y(n5183) );
  MX4X1 U6793 ( .A(\ram[200][6] ), .B(\ram[201][6] ), .C(\ram[202][6] ), .D(
        \ram[203][6] ), .S0(n6300), .S1(n6166), .Y(n5193) );
  MX4X1 U6794 ( .A(\ram[216][7] ), .B(\ram[217][7] ), .C(\ram[218][7] ), .D(
        \ram[219][7] ), .S0(n6305), .S1(n6171), .Y(n5272) );
  MX4X1 U6795 ( .A(\ram[232][7] ), .B(\ram[233][7] ), .C(\ram[234][7] ), .D(
        \ram[235][7] ), .S0(n6305), .S1(n6171), .Y(n5267) );
  MX4X1 U6796 ( .A(\ram[200][7] ), .B(\ram[201][7] ), .C(\ram[202][7] ), .D(
        \ram[203][7] ), .S0(n6306), .S1(n6172), .Y(n5277) );
  MX4X1 U6797 ( .A(\ram[216][8] ), .B(\ram[217][8] ), .C(\ram[218][8] ), .D(
        \ram[219][8] ), .S0(n6311), .S1(n6177), .Y(n5356) );
  MX4X1 U6798 ( .A(\ram[232][8] ), .B(\ram[233][8] ), .C(\ram[234][8] ), .D(
        \ram[235][8] ), .S0(n6310), .S1(n6176), .Y(n5351) );
  MX4X1 U6799 ( .A(\ram[200][8] ), .B(\ram[201][8] ), .C(\ram[202][8] ), .D(
        \ram[203][8] ), .S0(n6311), .S1(n6177), .Y(n5361) );
  MX4X1 U6800 ( .A(\ram[216][9] ), .B(\ram[217][9] ), .C(\ram[218][9] ), .D(
        \ram[219][9] ), .S0(n6316), .S1(n6182), .Y(n5440) );
  MX4X1 U6801 ( .A(\ram[232][9] ), .B(\ram[233][9] ), .C(\ram[234][9] ), .D(
        \ram[235][9] ), .S0(n6316), .S1(n6182), .Y(n5435) );
  MX4X1 U6802 ( .A(\ram[200][9] ), .B(\ram[201][9] ), .C(\ram[202][9] ), .D(
        \ram[203][9] ), .S0(n6316), .S1(n6182), .Y(n5445) );
  MX4X1 U6803 ( .A(\ram[216][10] ), .B(\ram[217][10] ), .C(\ram[218][10] ), 
        .D(\ram[219][10] ), .S0(n6321), .S1(n6187), .Y(n5524) );
  MX4X1 U6804 ( .A(\ram[232][10] ), .B(\ram[233][10] ), .C(\ram[234][10] ), 
        .D(\ram[235][10] ), .S0(n6321), .S1(n6187), .Y(n5519) );
  MX4X1 U6805 ( .A(\ram[200][10] ), .B(\ram[201][10] ), .C(\ram[202][10] ), 
        .D(\ram[203][10] ), .S0(n6322), .S1(n6188), .Y(n5529) );
  MX4X1 U6806 ( .A(\ram[216][11] ), .B(\ram[217][11] ), .C(\ram[218][11] ), 
        .D(\ram[219][11] ), .S0(n6327), .S1(n6193), .Y(n5608) );
  MX4X1 U6807 ( .A(\ram[232][11] ), .B(\ram[233][11] ), .C(\ram[234][11] ), 
        .D(\ram[235][11] ), .S0(n6326), .S1(n6192), .Y(n5603) );
  MX4X1 U6808 ( .A(\ram[200][11] ), .B(\ram[201][11] ), .C(\ram[202][11] ), 
        .D(\ram[203][11] ), .S0(n6327), .S1(n6193), .Y(n5613) );
  MX4X1 U6809 ( .A(\ram[216][12] ), .B(\ram[217][12] ), .C(\ram[218][12] ), 
        .D(\ram[219][12] ), .S0(n6332), .S1(n6198), .Y(n5692) );
  MX4X1 U6810 ( .A(\ram[232][12] ), .B(\ram[233][12] ), .C(\ram[234][12] ), 
        .D(\ram[235][12] ), .S0(n6332), .S1(n6198), .Y(n5687) );
  MX4X1 U6811 ( .A(\ram[200][12] ), .B(\ram[201][12] ), .C(\ram[202][12] ), 
        .D(\ram[203][12] ), .S0(n6332), .S1(n6198), .Y(n5697) );
  MX4X1 U6812 ( .A(\ram[216][13] ), .B(\ram[217][13] ), .C(\ram[218][13] ), 
        .D(\ram[219][13] ), .S0(n6337), .S1(n6203), .Y(n5776) );
  MX4X1 U6813 ( .A(\ram[232][13] ), .B(\ram[233][13] ), .C(\ram[234][13] ), 
        .D(\ram[235][13] ), .S0(n6337), .S1(n6203), .Y(n5771) );
  MX4X1 U6814 ( .A(\ram[200][13] ), .B(\ram[201][13] ), .C(\ram[202][13] ), 
        .D(\ram[203][13] ), .S0(n6338), .S1(n6204), .Y(n5781) );
  MX4X1 U6815 ( .A(\ram[216][14] ), .B(\ram[217][14] ), .C(\ram[218][14] ), 
        .D(\ram[219][14] ), .S0(n6343), .S1(n6209), .Y(n5860) );
  MX4X1 U6816 ( .A(\ram[232][14] ), .B(\ram[233][14] ), .C(\ram[234][14] ), 
        .D(\ram[235][14] ), .S0(n6342), .S1(n6208), .Y(n5855) );
  MX4X1 U6817 ( .A(\ram[200][14] ), .B(\ram[201][14] ), .C(\ram[202][14] ), 
        .D(\ram[203][14] ), .S0(n6343), .S1(n6209), .Y(n5865) );
  MX4X1 U6818 ( .A(\ram[216][15] ), .B(\ram[217][15] ), .C(\ram[218][15] ), 
        .D(\ram[219][15] ), .S0(n6348), .S1(n6213), .Y(n5944) );
  MX4X1 U6819 ( .A(\ram[232][15] ), .B(\ram[233][15] ), .C(\ram[234][15] ), 
        .D(\ram[235][15] ), .S0(n6348), .S1(n6213), .Y(n5939) );
  MX4X1 U6820 ( .A(\ram[200][15] ), .B(\ram[201][15] ), .C(\ram[202][15] ), 
        .D(\ram[203][15] ), .S0(n6348), .S1(n6213), .Y(n5949) );
  MX4X1 U6821 ( .A(n4702), .B(n4700), .C(n4701), .D(n4699), .S0(n6035), .S1(
        n6073), .Y(n4703) );
  MX4X1 U6822 ( .A(\ram[160][0] ), .B(\ram[161][0] ), .C(\ram[162][0] ), .D(
        \ram[163][0] ), .S0(n6269), .S1(n6135), .Y(n4702) );
  MX4X1 U6823 ( .A(\ram[168][0] ), .B(\ram[169][0] ), .C(\ram[170][0] ), .D(
        \ram[171][0] ), .S0(n6269), .S1(n6135), .Y(n4700) );
  MX4X1 U6824 ( .A(\ram[164][0] ), .B(\ram[165][0] ), .C(\ram[166][0] ), .D(
        \ram[167][0] ), .S0(n6269), .S1(n6135), .Y(n4701) );
  MX4X1 U6825 ( .A(n4744), .B(n4742), .C(n4743), .D(n4741), .S0(n6043), .S1(
        n6059), .Y(n4745) );
  MX4X1 U6826 ( .A(\ram[32][0] ), .B(\ram[33][0] ), .C(\ram[34][0] ), .D(
        \ram[35][0] ), .S0(n6272), .S1(n6138), .Y(n4744) );
  MX4X1 U6827 ( .A(\ram[40][0] ), .B(\ram[41][0] ), .C(\ram[42][0] ), .D(
        \ram[43][0] ), .S0(n6272), .S1(n6138), .Y(n4742) );
  MX4X1 U6828 ( .A(\ram[36][0] ), .B(\ram[37][0] ), .C(\ram[38][0] ), .D(
        \ram[39][0] ), .S0(n6272), .S1(n6138), .Y(n4743) );
  MX4X1 U6829 ( .A(n4807), .B(n4805), .C(n4806), .D(n4804), .S0(n6033), .S1(
        n6056), .Y(n4808) );
  MX4X1 U6830 ( .A(\ram[96][1] ), .B(\ram[97][1] ), .C(\ram[98][1] ), .D(
        \ram[99][1] ), .S0(n6276), .S1(n6142), .Y(n4807) );
  MX4X1 U6831 ( .A(\ram[104][1] ), .B(\ram[105][1] ), .C(\ram[106][1] ), .D(
        \ram[107][1] ), .S0(n6276), .S1(n6142), .Y(n4805) );
  MX4X1 U6832 ( .A(\ram[100][1] ), .B(\ram[101][1] ), .C(\ram[102][1] ), .D(
        \ram[103][1] ), .S0(n6276), .S1(n6142), .Y(n4806) );
  MX4X1 U6833 ( .A(n4786), .B(n4784), .C(n4785), .D(n4783), .S0(n6033), .S1(
        n6056), .Y(n4787) );
  MX4X1 U6834 ( .A(\ram[160][1] ), .B(\ram[161][1] ), .C(\ram[162][1] ), .D(
        \ram[163][1] ), .S0(n6274), .S1(n6140), .Y(n4786) );
  MX4X1 U6835 ( .A(\ram[168][1] ), .B(\ram[169][1] ), .C(\ram[170][1] ), .D(
        \ram[171][1] ), .S0(n6274), .S1(n6140), .Y(n4784) );
  MX4X1 U6836 ( .A(\ram[164][1] ), .B(\ram[165][1] ), .C(\ram[166][1] ), .D(
        \ram[167][1] ), .S0(n6274), .S1(n6140), .Y(n4785) );
  MX4X1 U6837 ( .A(n4828), .B(n4826), .C(n4827), .D(n4825), .S0(n6042), .S1(
        n6057), .Y(n4829) );
  MX4X1 U6838 ( .A(\ram[32][1] ), .B(\ram[33][1] ), .C(\ram[34][1] ), .D(
        \ram[35][1] ), .S0(n6277), .S1(n6143), .Y(n4828) );
  MX4X1 U6839 ( .A(\ram[40][1] ), .B(\ram[41][1] ), .C(\ram[42][1] ), .D(
        \ram[43][1] ), .S0(n6277), .S1(n6143), .Y(n4826) );
  MX4X1 U6840 ( .A(\ram[36][1] ), .B(\ram[37][1] ), .C(\ram[38][1] ), .D(
        \ram[39][1] ), .S0(n6277), .S1(n6143), .Y(n4827) );
  MX4X1 U6841 ( .A(n4891), .B(n4889), .C(n4890), .D(n4888), .S0(n6047), .S1(
        n6058), .Y(n4892) );
  MX4X1 U6842 ( .A(\ram[96][2] ), .B(\ram[97][2] ), .C(\ram[98][2] ), .D(
        \ram[99][2] ), .S0(n6281), .S1(n6147), .Y(n4891) );
  MX4X1 U6843 ( .A(\ram[104][2] ), .B(\ram[105][2] ), .C(\ram[106][2] ), .D(
        \ram[107][2] ), .S0(n6281), .S1(n6147), .Y(n4889) );
  MX4X1 U6844 ( .A(\ram[100][2] ), .B(\ram[101][2] ), .C(\ram[102][2] ), .D(
        \ram[103][2] ), .S0(n6281), .S1(n6147), .Y(n4890) );
  MX4X1 U6845 ( .A(n4870), .B(n4868), .C(n4869), .D(n4867), .S0(n6046), .S1(
        n6057), .Y(n4871) );
  MX4X1 U6846 ( .A(\ram[160][2] ), .B(\ram[161][2] ), .C(\ram[162][2] ), .D(
        \ram[163][2] ), .S0(n6280), .S1(n6146), .Y(n4870) );
  MX4X1 U6847 ( .A(\ram[168][2] ), .B(\ram[169][2] ), .C(\ram[170][2] ), .D(
        \ram[171][2] ), .S0(n6280), .S1(n6146), .Y(n4868) );
  MX4X1 U6848 ( .A(\ram[164][2] ), .B(\ram[165][2] ), .C(\ram[166][2] ), .D(
        \ram[167][2] ), .S0(n6280), .S1(n6146), .Y(n4869) );
  MX4X1 U6849 ( .A(n4912), .B(n4910), .C(n4911), .D(n4909), .S0(n6038), .S1(
        n6058), .Y(n4913) );
  MX4X1 U6850 ( .A(\ram[32][2] ), .B(\ram[33][2] ), .C(\ram[34][2] ), .D(
        \ram[35][2] ), .S0(n6282), .S1(n6148), .Y(n4912) );
  MX4X1 U6851 ( .A(\ram[40][2] ), .B(\ram[41][2] ), .C(\ram[42][2] ), .D(
        \ram[43][2] ), .S0(n6282), .S1(n6148), .Y(n4910) );
  MX4X1 U6852 ( .A(\ram[36][2] ), .B(\ram[37][2] ), .C(\ram[38][2] ), .D(
        \ram[39][2] ), .S0(n6282), .S1(n6148), .Y(n4911) );
  MX4X1 U6853 ( .A(n4933), .B(n4931), .C(n4932), .D(n4930), .S0(n6046), .S1(
        n6058), .Y(n4934) );
  MX4X1 U6854 ( .A(\ram[224][3] ), .B(\ram[225][3] ), .C(\ram[226][3] ), .D(
        \ram[227][3] ), .S0(n6284), .S1(n6150), .Y(n4933) );
  MX4X1 U6855 ( .A(\ram[232][3] ), .B(\ram[233][3] ), .C(\ram[234][3] ), .D(
        \ram[235][3] ), .S0(n6284), .S1(n6150), .Y(n4931) );
  MX4X1 U6856 ( .A(\ram[228][3] ), .B(\ram[229][3] ), .C(\ram[230][3] ), .D(
        \ram[231][3] ), .S0(n6284), .S1(n6150), .Y(n4932) );
  MX4X1 U6857 ( .A(n4996), .B(n4994), .C(n4995), .D(n4993), .S0(n6026), .S1(
        n6059), .Y(n4997) );
  MX4X1 U6858 ( .A(\ram[32][3] ), .B(\ram[33][3] ), .C(\ram[34][3] ), .D(
        \ram[35][3] ), .S0(n6288), .S1(n6154), .Y(n4996) );
  MX4X1 U6859 ( .A(\ram[40][3] ), .B(\ram[41][3] ), .C(\ram[42][3] ), .D(
        \ram[43][3] ), .S0(n6288), .S1(n6154), .Y(n4994) );
  MX4X1 U6860 ( .A(\ram[36][3] ), .B(\ram[37][3] ), .C(\ram[38][3] ), .D(
        \ram[39][3] ), .S0(n6288), .S1(n6154), .Y(n4995) );
  MX4X1 U6861 ( .A(n4954), .B(n4952), .C(n4953), .D(n4951), .S0(n6046), .S1(
        n6059), .Y(n4955) );
  MX4X1 U6862 ( .A(\ram[160][3] ), .B(\ram[161][3] ), .C(\ram[162][3] ), .D(
        \ram[163][3] ), .S0(n6285), .S1(n6151), .Y(n4954) );
  MX4X1 U6863 ( .A(\ram[168][3] ), .B(\ram[169][3] ), .C(\ram[170][3] ), .D(
        \ram[171][3] ), .S0(n6285), .S1(n6151), .Y(n4952) );
  MX4X1 U6864 ( .A(\ram[164][3] ), .B(\ram[165][3] ), .C(\ram[166][3] ), .D(
        \ram[167][3] ), .S0(n6285), .S1(n6151), .Y(n4953) );
  MX4X1 U6865 ( .A(n5059), .B(n5057), .C(n5058), .D(n5056), .S0(n6034), .S1(
        n6060), .Y(n5060) );
  MX4X1 U6866 ( .A(\ram[96][4] ), .B(\ram[97][4] ), .C(\ram[98][4] ), .D(
        \ram[99][4] ), .S0(n6292), .S1(n6158), .Y(n5059) );
  MX4X1 U6867 ( .A(\ram[104][4] ), .B(\ram[105][4] ), .C(\ram[106][4] ), .D(
        \ram[107][4] ), .S0(n6292), .S1(n6158), .Y(n5057) );
  MX4X1 U6868 ( .A(\ram[100][4] ), .B(\ram[101][4] ), .C(\ram[102][4] ), .D(
        \ram[103][4] ), .S0(n6292), .S1(n6158), .Y(n5058) );
  MX4X1 U6869 ( .A(n5038), .B(n5036), .C(n5037), .D(n5035), .S0(n6034), .S1(
        n6060), .Y(n5039) );
  MX4X1 U6870 ( .A(\ram[160][4] ), .B(\ram[161][4] ), .C(\ram[162][4] ), .D(
        \ram[163][4] ), .S0(n6290), .S1(n6156), .Y(n5038) );
  MX4X1 U6871 ( .A(\ram[168][4] ), .B(\ram[169][4] ), .C(\ram[170][4] ), .D(
        \ram[171][4] ), .S0(n6290), .S1(n6156), .Y(n5036) );
  MX4X1 U6872 ( .A(\ram[164][4] ), .B(\ram[165][4] ), .C(\ram[166][4] ), .D(
        \ram[167][4] ), .S0(n6290), .S1(n6156), .Y(n5037) );
  MX4X1 U6873 ( .A(n5080), .B(n5078), .C(n5079), .D(n5077), .S0(n6044), .S1(
        n6061), .Y(n5081) );
  MX4X1 U6874 ( .A(\ram[32][4] ), .B(\ram[33][4] ), .C(\ram[34][4] ), .D(
        \ram[35][4] ), .S0(n6293), .S1(n6159), .Y(n5080) );
  MX4X1 U6875 ( .A(\ram[40][4] ), .B(\ram[41][4] ), .C(\ram[42][4] ), .D(
        \ram[43][4] ), .S0(n6293), .S1(n6159), .Y(n5078) );
  MX4X1 U6876 ( .A(\ram[36][4] ), .B(\ram[37][4] ), .C(\ram[38][4] ), .D(
        \ram[39][4] ), .S0(n6293), .S1(n6159), .Y(n5079) );
  MX4X1 U6877 ( .A(n5143), .B(n5141), .C(n5142), .D(n5140), .S0(n6035), .S1(
        n6062), .Y(n5144) );
  MX4X1 U6878 ( .A(\ram[96][5] ), .B(\ram[97][5] ), .C(\ram[98][5] ), .D(
        \ram[99][5] ), .S0(n6297), .S1(n6163), .Y(n5143) );
  MX4X1 U6879 ( .A(\ram[104][5] ), .B(\ram[105][5] ), .C(\ram[106][5] ), .D(
        \ram[107][5] ), .S0(n6297), .S1(n6163), .Y(n5141) );
  MX4X1 U6880 ( .A(\ram[100][5] ), .B(\ram[101][5] ), .C(\ram[102][5] ), .D(
        \ram[103][5] ), .S0(n6297), .S1(n6163), .Y(n5142) );
  MX4X1 U6881 ( .A(n5122), .B(n5120), .C(n5121), .D(n5119), .S0(n6035), .S1(
        n6061), .Y(n5123) );
  MX4X1 U6882 ( .A(\ram[160][5] ), .B(\ram[161][5] ), .C(\ram[162][5] ), .D(
        \ram[163][5] ), .S0(n6296), .S1(n6162), .Y(n5122) );
  MX4X1 U6883 ( .A(\ram[168][5] ), .B(\ram[169][5] ), .C(\ram[170][5] ), .D(
        \ram[171][5] ), .S0(n6296), .S1(n6162), .Y(n5120) );
  MX4X1 U6884 ( .A(\ram[164][5] ), .B(\ram[165][5] ), .C(\ram[166][5] ), .D(
        \ram[167][5] ), .S0(n6296), .S1(n6162), .Y(n5121) );
  MX4X1 U6885 ( .A(n5164), .B(n5162), .C(n5163), .D(n5161), .S0(n6035), .S1(
        n6062), .Y(n5165) );
  MX4X1 U6886 ( .A(\ram[32][5] ), .B(\ram[33][5] ), .C(\ram[34][5] ), .D(
        \ram[35][5] ), .S0(n6298), .S1(n6164), .Y(n5164) );
  MX4X1 U6887 ( .A(\ram[40][5] ), .B(\ram[41][5] ), .C(\ram[42][5] ), .D(
        \ram[43][5] ), .S0(n6298), .S1(n6164), .Y(n5162) );
  MX4X1 U6888 ( .A(\ram[36][5] ), .B(\ram[37][5] ), .C(\ram[38][5] ), .D(
        \ram[39][5] ), .S0(n6298), .S1(n6164), .Y(n5163) );
  MX4X1 U6889 ( .A(n5227), .B(n5225), .C(n5226), .D(n5224), .S0(n6035), .S1(
        n6063), .Y(n5228) );
  MX4X1 U6890 ( .A(\ram[96][6] ), .B(\ram[97][6] ), .C(\ram[98][6] ), .D(
        \ram[99][6] ), .S0(n6302), .S1(n6168), .Y(n5227) );
  MX4X1 U6891 ( .A(\ram[104][6] ), .B(\ram[105][6] ), .C(\ram[106][6] ), .D(
        \ram[107][6] ), .S0(n6302), .S1(n6168), .Y(n5225) );
  MX4X1 U6892 ( .A(\ram[100][6] ), .B(\ram[101][6] ), .C(\ram[102][6] ), .D(
        \ram[103][6] ), .S0(n6302), .S1(n6168), .Y(n5226) );
  MX4X1 U6893 ( .A(n5206), .B(n5204), .C(n5205), .D(n5203), .S0(n6040), .S1(
        n6063), .Y(n5207) );
  MX4X1 U6894 ( .A(\ram[160][6] ), .B(\ram[161][6] ), .C(\ram[162][6] ), .D(
        \ram[163][6] ), .S0(n6301), .S1(n6167), .Y(n5206) );
  MX4X1 U6895 ( .A(\ram[168][6] ), .B(\ram[169][6] ), .C(\ram[170][6] ), .D(
        \ram[171][6] ), .S0(n6301), .S1(n6167), .Y(n5204) );
  MX4X1 U6896 ( .A(\ram[164][6] ), .B(\ram[165][6] ), .C(\ram[166][6] ), .D(
        \ram[167][6] ), .S0(n6301), .S1(n6167), .Y(n5205) );
  MX4X1 U6897 ( .A(n5248), .B(n5246), .C(n5247), .D(n5245), .S0(n6034), .S1(
        n6063), .Y(n5249) );
  MX4X1 U6898 ( .A(\ram[32][6] ), .B(\ram[33][6] ), .C(\ram[34][6] ), .D(
        \ram[35][6] ), .S0(n6304), .S1(n6170), .Y(n5248) );
  MX4X1 U6899 ( .A(\ram[40][6] ), .B(\ram[41][6] ), .C(\ram[42][6] ), .D(
        \ram[43][6] ), .S0(n6304), .S1(n6170), .Y(n5246) );
  MX4X1 U6900 ( .A(\ram[36][6] ), .B(\ram[37][6] ), .C(\ram[38][6] ), .D(
        \ram[39][6] ), .S0(n6304), .S1(n6170), .Y(n5247) );
  MX4X1 U6901 ( .A(n5311), .B(n5309), .C(n5310), .D(n5308), .S0(n6036), .S1(
        n6064), .Y(n5312) );
  MX4X1 U6902 ( .A(\ram[96][7] ), .B(\ram[97][7] ), .C(\ram[98][7] ), .D(
        \ram[99][7] ), .S0(n6308), .S1(n6174), .Y(n5311) );
  MX4X1 U6903 ( .A(\ram[104][7] ), .B(\ram[105][7] ), .C(\ram[106][7] ), .D(
        \ram[107][7] ), .S0(n6308), .S1(n6174), .Y(n5309) );
  MX4X1 U6904 ( .A(\ram[100][7] ), .B(\ram[101][7] ), .C(\ram[102][7] ), .D(
        \ram[103][7] ), .S0(n6308), .S1(n6174), .Y(n5310) );
  MX4X1 U6905 ( .A(n5290), .B(n5288), .C(n5289), .D(n5287), .S0(n6036), .S1(
        n6064), .Y(n5291) );
  MX4X1 U6906 ( .A(\ram[160][7] ), .B(\ram[161][7] ), .C(\ram[162][7] ), .D(
        \ram[163][7] ), .S0(n6306), .S1(n6172), .Y(n5290) );
  MX4X1 U6907 ( .A(\ram[168][7] ), .B(\ram[169][7] ), .C(\ram[170][7] ), .D(
        \ram[171][7] ), .S0(n6306), .S1(n6172), .Y(n5288) );
  MX4X1 U6908 ( .A(\ram[164][7] ), .B(\ram[165][7] ), .C(\ram[166][7] ), .D(
        \ram[167][7] ), .S0(n6306), .S1(n6172), .Y(n5289) );
  MX4X1 U6909 ( .A(n5332), .B(n5330), .C(n5331), .D(n5329), .S0(n6037), .S1(
        n6065), .Y(n5333) );
  MX4X1 U6910 ( .A(\ram[32][7] ), .B(\ram[33][7] ), .C(\ram[34][7] ), .D(
        \ram[35][7] ), .S0(n6309), .S1(n6175), .Y(n5332) );
  MX4X1 U6911 ( .A(\ram[40][7] ), .B(\ram[41][7] ), .C(\ram[42][7] ), .D(
        \ram[43][7] ), .S0(n6309), .S1(n6175), .Y(n5330) );
  MX4X1 U6912 ( .A(\ram[36][7] ), .B(\ram[37][7] ), .C(\ram[38][7] ), .D(
        \ram[39][7] ), .S0(n6309), .S1(n6175), .Y(n5331) );
  MX4X1 U6913 ( .A(n5395), .B(n5393), .C(n5394), .D(n5392), .S0(n6038), .S1(
        n6066), .Y(n5396) );
  MX4X1 U6914 ( .A(\ram[96][8] ), .B(\ram[97][8] ), .C(\ram[98][8] ), .D(
        \ram[99][8] ), .S0(n6313), .S1(n6179), .Y(n5395) );
  MX4X1 U6915 ( .A(\ram[104][8] ), .B(\ram[105][8] ), .C(\ram[106][8] ), .D(
        \ram[107][8] ), .S0(n6313), .S1(n6179), .Y(n5393) );
  MX4X1 U6916 ( .A(\ram[100][8] ), .B(\ram[101][8] ), .C(\ram[102][8] ), .D(
        \ram[103][8] ), .S0(n6313), .S1(n6179), .Y(n5394) );
  MX4X1 U6917 ( .A(n5374), .B(n5372), .C(n5373), .D(n5371), .S0(n6037), .S1(
        n6065), .Y(n5375) );
  MX4X1 U6918 ( .A(\ram[160][8] ), .B(\ram[161][8] ), .C(\ram[162][8] ), .D(
        \ram[163][8] ), .S0(n6312), .S1(n6178), .Y(n5374) );
  MX4X1 U6919 ( .A(\ram[168][8] ), .B(\ram[169][8] ), .C(\ram[170][8] ), .D(
        \ram[171][8] ), .S0(n6312), .S1(n6178), .Y(n5372) );
  MX4X1 U6920 ( .A(\ram[164][8] ), .B(\ram[165][8] ), .C(\ram[166][8] ), .D(
        \ram[167][8] ), .S0(n6312), .S1(n6178), .Y(n5373) );
  MX4X1 U6921 ( .A(n5416), .B(n5414), .C(n5415), .D(n5413), .S0(n6038), .S1(
        n6066), .Y(n5417) );
  MX4X1 U6922 ( .A(\ram[32][8] ), .B(\ram[33][8] ), .C(\ram[34][8] ), .D(
        \ram[35][8] ), .S0(n6314), .S1(n6180), .Y(n5416) );
  MX4X1 U6923 ( .A(\ram[40][8] ), .B(\ram[41][8] ), .C(\ram[42][8] ), .D(
        \ram[43][8] ), .S0(n6314), .S1(n6180), .Y(n5414) );
  MX4X1 U6924 ( .A(\ram[36][8] ), .B(\ram[37][8] ), .C(\ram[38][8] ), .D(
        \ram[39][8] ), .S0(n6314), .S1(n6180), .Y(n5415) );
  MX4X1 U6925 ( .A(n5479), .B(n5477), .C(n5478), .D(n5476), .S0(n6039), .S1(
        n6067), .Y(n5480) );
  MX4X1 U6926 ( .A(\ram[96][9] ), .B(\ram[97][9] ), .C(\ram[98][9] ), .D(
        \ram[99][9] ), .S0(n6318), .S1(n6184), .Y(n5479) );
  MX4X1 U6927 ( .A(\ram[104][9] ), .B(\ram[105][9] ), .C(\ram[106][9] ), .D(
        \ram[107][9] ), .S0(n6318), .S1(n6184), .Y(n5477) );
  MX4X1 U6928 ( .A(\ram[100][9] ), .B(\ram[101][9] ), .C(\ram[102][9] ), .D(
        \ram[103][9] ), .S0(n6318), .S1(n6184), .Y(n5478) );
  MX4X1 U6929 ( .A(n5458), .B(n5456), .C(n5457), .D(n5455), .S0(n6039), .S1(
        n6067), .Y(n5459) );
  MX4X1 U6930 ( .A(\ram[160][9] ), .B(\ram[161][9] ), .C(\ram[162][9] ), .D(
        \ram[163][9] ), .S0(n6317), .S1(n6183), .Y(n5458) );
  MX4X1 U6931 ( .A(\ram[168][9] ), .B(\ram[169][9] ), .C(\ram[170][9] ), .D(
        \ram[171][9] ), .S0(n6317), .S1(n6183), .Y(n5456) );
  MX4X1 U6932 ( .A(\ram[164][9] ), .B(\ram[165][9] ), .C(\ram[166][9] ), .D(
        \ram[167][9] ), .S0(n6317), .S1(n6183), .Y(n5457) );
  MX4X1 U6933 ( .A(n5500), .B(n5498), .C(n5499), .D(n5497), .S0(n6039), .S1(
        n6067), .Y(n5501) );
  MX4X1 U6934 ( .A(\ram[32][9] ), .B(\ram[33][9] ), .C(\ram[34][9] ), .D(
        \ram[35][9] ), .S0(n6320), .S1(n6186), .Y(n5500) );
  MX4X1 U6935 ( .A(\ram[40][9] ), .B(\ram[41][9] ), .C(\ram[42][9] ), .D(
        \ram[43][9] ), .S0(n6320), .S1(n6186), .Y(n5498) );
  MX4X1 U6936 ( .A(\ram[36][9] ), .B(\ram[37][9] ), .C(\ram[38][9] ), .D(
        \ram[39][9] ), .S0(n6320), .S1(n6186), .Y(n5499) );
  MX4X1 U6937 ( .A(n5542), .B(n5540), .C(n5541), .D(n5539), .S0(n6040), .S1(
        n6068), .Y(n5543) );
  MX4X1 U6938 ( .A(\ram[160][10] ), .B(\ram[161][10] ), .C(\ram[162][10] ), 
        .D(\ram[163][10] ), .S0(n6322), .S1(n6188), .Y(n5542) );
  MX4X1 U6939 ( .A(\ram[168][10] ), .B(\ram[169][10] ), .C(\ram[170][10] ), 
        .D(\ram[171][10] ), .S0(n6322), .S1(n6188), .Y(n5540) );
  MX4X1 U6940 ( .A(\ram[164][10] ), .B(\ram[165][10] ), .C(\ram[166][10] ), 
        .D(\ram[167][10] ), .S0(n6322), .S1(n6188), .Y(n5541) );
  MX4X1 U6941 ( .A(n5563), .B(n5561), .C(n5562), .D(n5560), .S0(n6040), .S1(
        n6068), .Y(n5564) );
  MX4X1 U6942 ( .A(\ram[96][10] ), .B(\ram[97][10] ), .C(\ram[98][10] ), .D(
        \ram[99][10] ), .S0(n6324), .S1(n6190), .Y(n5563) );
  MX4X1 U6943 ( .A(\ram[104][10] ), .B(\ram[105][10] ), .C(\ram[106][10] ), 
        .D(\ram[107][10] ), .S0(n6324), .S1(n6190), .Y(n5561) );
  MX4X1 U6944 ( .A(\ram[100][10] ), .B(\ram[101][10] ), .C(\ram[102][10] ), 
        .D(\ram[103][10] ), .S0(n6324), .S1(n6190), .Y(n5562) );
  MX4X1 U6945 ( .A(n5584), .B(n5582), .C(n5583), .D(n5581), .S0(n6041), .S1(
        n6069), .Y(n5585) );
  MX4X1 U6946 ( .A(\ram[32][10] ), .B(\ram[33][10] ), .C(\ram[34][10] ), .D(
        \ram[35][10] ), .S0(n6325), .S1(n6191), .Y(n5584) );
  MX4X1 U6947 ( .A(\ram[40][10] ), .B(\ram[41][10] ), .C(\ram[42][10] ), .D(
        \ram[43][10] ), .S0(n6325), .S1(n6191), .Y(n5582) );
  MX4X1 U6948 ( .A(\ram[36][10] ), .B(\ram[37][10] ), .C(\ram[38][10] ), .D(
        \ram[39][10] ), .S0(n6325), .S1(n6191), .Y(n5583) );
  MX4X1 U6949 ( .A(n5647), .B(n5645), .C(n5646), .D(n5644), .S0(n6042), .S1(
        n6070), .Y(n5648) );
  MX4X1 U6950 ( .A(\ram[96][11] ), .B(\ram[97][11] ), .C(\ram[98][11] ), .D(
        \ram[99][11] ), .S0(n6329), .S1(n6195), .Y(n5647) );
  MX4X1 U6951 ( .A(\ram[104][11] ), .B(\ram[105][11] ), .C(\ram[106][11] ), 
        .D(\ram[107][11] ), .S0(n6329), .S1(n6195), .Y(n5645) );
  MX4X1 U6952 ( .A(\ram[100][11] ), .B(\ram[101][11] ), .C(\ram[102][11] ), 
        .D(\ram[103][11] ), .S0(n6329), .S1(n6195), .Y(n5646) );
  MX4X1 U6953 ( .A(n5626), .B(n5624), .C(n5625), .D(n5623), .S0(n6041), .S1(
        n6069), .Y(n5627) );
  MX4X1 U6954 ( .A(\ram[160][11] ), .B(\ram[161][11] ), .C(\ram[162][11] ), 
        .D(\ram[163][11] ), .S0(n6328), .S1(n6194), .Y(n5626) );
  MX4X1 U6955 ( .A(\ram[168][11] ), .B(\ram[169][11] ), .C(\ram[170][11] ), 
        .D(\ram[171][11] ), .S0(n6328), .S1(n6194), .Y(n5624) );
  MX4X1 U6956 ( .A(\ram[164][11] ), .B(\ram[165][11] ), .C(\ram[166][11] ), 
        .D(\ram[167][11] ), .S0(n6328), .S1(n6194), .Y(n5625) );
  MX4X1 U6957 ( .A(n5668), .B(n5666), .C(n5667), .D(n5665), .S0(n6042), .S1(
        n6070), .Y(n5669) );
  MX4X1 U6958 ( .A(\ram[32][11] ), .B(\ram[33][11] ), .C(\ram[34][11] ), .D(
        \ram[35][11] ), .S0(n6330), .S1(n6196), .Y(n5668) );
  MX4X1 U6959 ( .A(\ram[40][11] ), .B(\ram[41][11] ), .C(\ram[42][11] ), .D(
        \ram[43][11] ), .S0(n6330), .S1(n6196), .Y(n5666) );
  MX4X1 U6960 ( .A(\ram[36][11] ), .B(\ram[37][11] ), .C(\ram[38][11] ), .D(
        \ram[39][11] ), .S0(n6330), .S1(n6196), .Y(n5667) );
  MX4X1 U6961 ( .A(n5731), .B(n5729), .C(n5730), .D(n5728), .S0(n6043), .S1(
        n6071), .Y(n5732) );
  MX4X1 U6962 ( .A(\ram[96][12] ), .B(\ram[97][12] ), .C(\ram[98][12] ), .D(
        \ram[99][12] ), .S0(n6334), .S1(n6200), .Y(n5731) );
  MX4X1 U6963 ( .A(\ram[104][12] ), .B(\ram[105][12] ), .C(\ram[106][12] ), 
        .D(\ram[107][12] ), .S0(n6334), .S1(n6200), .Y(n5729) );
  MX4X1 U6964 ( .A(\ram[100][12] ), .B(\ram[101][12] ), .C(\ram[102][12] ), 
        .D(\ram[103][12] ), .S0(n6334), .S1(n6200), .Y(n5730) );
  MX4X1 U6965 ( .A(n5710), .B(n5708), .C(n5709), .D(n5707), .S0(n6043), .S1(
        n6071), .Y(n5711) );
  MX4X1 U6966 ( .A(\ram[160][12] ), .B(\ram[161][12] ), .C(\ram[162][12] ), 
        .D(\ram[163][12] ), .S0(n6333), .S1(n6199), .Y(n5710) );
  MX4X1 U6967 ( .A(\ram[168][12] ), .B(\ram[169][12] ), .C(\ram[170][12] ), 
        .D(\ram[171][12] ), .S0(n6333), .S1(n6199), .Y(n5708) );
  MX4X1 U6968 ( .A(\ram[164][12] ), .B(\ram[165][12] ), .C(\ram[166][12] ), 
        .D(\ram[167][12] ), .S0(n6333), .S1(n6199), .Y(n5709) );
  MX4X1 U6969 ( .A(n5752), .B(n5750), .C(n5751), .D(n5749), .S0(n6043), .S1(
        n6071), .Y(n5753) );
  MX4X1 U6970 ( .A(\ram[32][12] ), .B(\ram[33][12] ), .C(\ram[34][12] ), .D(
        \ram[35][12] ), .S0(n6336), .S1(n6202), .Y(n5752) );
  MX4X1 U6971 ( .A(\ram[40][12] ), .B(\ram[41][12] ), .C(\ram[42][12] ), .D(
        \ram[43][12] ), .S0(n6336), .S1(n6202), .Y(n5750) );
  MX4X1 U6972 ( .A(\ram[36][12] ), .B(\ram[37][12] ), .C(\ram[38][12] ), .D(
        \ram[39][12] ), .S0(n6336), .S1(n6202), .Y(n5751) );
  MX4X1 U6973 ( .A(n5815), .B(n5813), .C(n5814), .D(n5812), .S0(n6044), .S1(
        n6072), .Y(n5816) );
  MX4X1 U6974 ( .A(\ram[96][13] ), .B(\ram[97][13] ), .C(\ram[98][13] ), .D(
        \ram[99][13] ), .S0(n6340), .S1(n6206), .Y(n5815) );
  MX4X1 U6975 ( .A(\ram[104][13] ), .B(\ram[105][13] ), .C(\ram[106][13] ), 
        .D(\ram[107][13] ), .S0(n6340), .S1(n6206), .Y(n5813) );
  MX4X1 U6976 ( .A(\ram[100][13] ), .B(\ram[101][13] ), .C(\ram[102][13] ), 
        .D(\ram[103][13] ), .S0(n6340), .S1(n6206), .Y(n5814) );
  MX4X1 U6977 ( .A(n5794), .B(n5792), .C(n5793), .D(n5791), .S0(n6044), .S1(
        n6072), .Y(n5795) );
  MX4X1 U6978 ( .A(\ram[160][13] ), .B(\ram[161][13] ), .C(\ram[162][13] ), 
        .D(\ram[163][13] ), .S0(n6338), .S1(n6204), .Y(n5794) );
  MX4X1 U6979 ( .A(\ram[168][13] ), .B(\ram[169][13] ), .C(\ram[170][13] ), 
        .D(\ram[171][13] ), .S0(n6338), .S1(n6204), .Y(n5792) );
  MX4X1 U6980 ( .A(\ram[164][13] ), .B(\ram[165][13] ), .C(\ram[166][13] ), 
        .D(\ram[167][13] ), .S0(n6338), .S1(n6204), .Y(n5793) );
  MX4X1 U6981 ( .A(n5836), .B(n5834), .C(n5835), .D(n5833), .S0(n6045), .S1(
        n6073), .Y(n5837) );
  MX4X1 U6982 ( .A(\ram[32][13] ), .B(\ram[33][13] ), .C(\ram[34][13] ), .D(
        \ram[35][13] ), .S0(n6341), .S1(n6207), .Y(n5836) );
  MX4X1 U6983 ( .A(\ram[40][13] ), .B(\ram[41][13] ), .C(\ram[42][13] ), .D(
        \ram[43][13] ), .S0(n6341), .S1(n6207), .Y(n5834) );
  MX4X1 U6984 ( .A(\ram[36][13] ), .B(\ram[37][13] ), .C(\ram[38][13] ), .D(
        \ram[39][13] ), .S0(n6341), .S1(n6207), .Y(n5835) );
  MX4X1 U6985 ( .A(n5899), .B(n5897), .C(n5898), .D(n5896), .S0(n6046), .S1(
        n6063), .Y(n5900) );
  MX4X1 U6986 ( .A(\ram[96][14] ), .B(\ram[97][14] ), .C(\ram[98][14] ), .D(
        \ram[99][14] ), .S0(n6345), .S1(n6211), .Y(n5899) );
  MX4X1 U6987 ( .A(\ram[104][14] ), .B(\ram[105][14] ), .C(\ram[106][14] ), 
        .D(\ram[107][14] ), .S0(n6345), .S1(n6211), .Y(n5897) );
  MX4X1 U6988 ( .A(\ram[100][14] ), .B(\ram[101][14] ), .C(\ram[102][14] ), 
        .D(\ram[103][14] ), .S0(n6345), .S1(n6211), .Y(n5898) );
  MX4X1 U6989 ( .A(n5878), .B(n5876), .C(n5877), .D(n5875), .S0(n6045), .S1(
        n6073), .Y(n5879) );
  MX4X1 U6990 ( .A(\ram[160][14] ), .B(\ram[161][14] ), .C(\ram[162][14] ), 
        .D(\ram[163][14] ), .S0(n6344), .S1(n6210), .Y(n5878) );
  MX4X1 U6991 ( .A(\ram[168][14] ), .B(\ram[169][14] ), .C(\ram[170][14] ), 
        .D(\ram[171][14] ), .S0(n6344), .S1(n6210), .Y(n5876) );
  MX4X1 U6992 ( .A(\ram[164][14] ), .B(\ram[165][14] ), .C(\ram[166][14] ), 
        .D(\ram[167][14] ), .S0(n6344), .S1(n6210), .Y(n5877) );
  MX4X1 U6993 ( .A(n5920), .B(n5918), .C(n5919), .D(n5917), .S0(n6046), .S1(
        n6061), .Y(n5921) );
  MX4X1 U6994 ( .A(\ram[32][14] ), .B(\ram[33][14] ), .C(\ram[34][14] ), .D(
        \ram[35][14] ), .S0(n6346), .S1(n6212), .Y(n5920) );
  MX4X1 U6995 ( .A(\ram[40][14] ), .B(\ram[41][14] ), .C(\ram[42][14] ), .D(
        \ram[43][14] ), .S0(n6346), .S1(n6212), .Y(n5918) );
  MX4X1 U6996 ( .A(\ram[36][14] ), .B(\ram[37][14] ), .C(\ram[38][14] ), .D(
        \ram[39][14] ), .S0(n6346), .S1(n6212), .Y(n5919) );
  MX4X1 U6997 ( .A(n5983), .B(n5981), .C(n5982), .D(n5980), .S0(n6047), .S1(
        n6061), .Y(n5984) );
  MX4X1 U6998 ( .A(\ram[96][15] ), .B(\ram[97][15] ), .C(\ram[98][15] ), .D(
        \ram[99][15] ), .S0(n6350), .S1(n6213), .Y(n5983) );
  MX4X1 U6999 ( .A(\ram[104][15] ), .B(\ram[105][15] ), .C(\ram[106][15] ), 
        .D(\ram[107][15] ), .S0(n6350), .S1(n6139), .Y(n5981) );
  MX4X1 U7000 ( .A(\ram[100][15] ), .B(\ram[101][15] ), .C(\ram[102][15] ), 
        .D(\ram[103][15] ), .S0(n6350), .S1(n6140), .Y(n5982) );
  MX4X1 U7001 ( .A(n5962), .B(n5960), .C(n5961), .D(n5959), .S0(n6047), .S1(
        n6063), .Y(n5963) );
  MX4X1 U7002 ( .A(\ram[160][15] ), .B(\ram[161][15] ), .C(\ram[162][15] ), 
        .D(\ram[163][15] ), .S0(n6349), .S1(n6214), .Y(n5962) );
  MX4X1 U7003 ( .A(\ram[168][15] ), .B(\ram[169][15] ), .C(\ram[170][15] ), 
        .D(\ram[171][15] ), .S0(n6349), .S1(n6214), .Y(n5960) );
  MX4X1 U7004 ( .A(\ram[164][15] ), .B(\ram[165][15] ), .C(\ram[166][15] ), 
        .D(\ram[167][15] ), .S0(n6349), .S1(n6214), .Y(n5961) );
  MX4X1 U7005 ( .A(n6004), .B(n6002), .C(n6003), .D(n6001), .S0(n6047), .S1(
        n6060), .Y(n6005) );
  MX4X1 U7006 ( .A(\ram[32][15] ), .B(\ram[33][15] ), .C(\ram[34][15] ), .D(
        \ram[35][15] ), .S0(n6352), .S1(n6214), .Y(n6004) );
  MX4X1 U7007 ( .A(\ram[40][15] ), .B(\ram[41][15] ), .C(\ram[42][15] ), .D(
        \ram[43][15] ), .S0(n6352), .S1(n6139), .Y(n6002) );
  MX4X1 U7008 ( .A(\ram[36][15] ), .B(\ram[37][15] ), .C(\ram[38][15] ), .D(
        \ram[39][15] ), .S0(n6352), .S1(n6139), .Y(n6003) );
  MX4X1 U7009 ( .A(n4686), .B(n4684), .C(n4685), .D(n4683), .S0(n6038), .S1(
        n6060), .Y(n4687) );
  MX4X1 U7010 ( .A(\ram[208][0] ), .B(\ram[209][0] ), .C(\ram[210][0] ), .D(
        \ram[211][0] ), .S0(n6268), .S1(n6134), .Y(n4686) );
  MX4X1 U7011 ( .A(\ram[216][0] ), .B(\ram[217][0] ), .C(\ram[218][0] ), .D(
        \ram[219][0] ), .S0(n6268), .S1(n6134), .Y(n4684) );
  MX4X1 U7012 ( .A(\ram[212][0] ), .B(\ram[213][0] ), .C(\ram[214][0] ), .D(
        \ram[215][0] ), .S0(n6268), .S1(n6134), .Y(n4685) );
  MX4X1 U7013 ( .A(n4691), .B(n4689), .C(n4690), .D(n4688), .S0(n6041), .S1(
        n6068), .Y(n4692) );
  MX4X1 U7014 ( .A(\ram[192][0] ), .B(\ram[193][0] ), .C(\ram[194][0] ), .D(
        \ram[195][0] ), .S0(n6268), .S1(n6134), .Y(n4691) );
  MX4X1 U7015 ( .A(\ram[200][0] ), .B(\ram[201][0] ), .C(\ram[202][0] ), .D(
        \ram[203][0] ), .S0(n6268), .S1(n6134), .Y(n4689) );
  MX4X1 U7016 ( .A(\ram[196][0] ), .B(\ram[197][0] ), .C(\ram[198][0] ), .D(
        \ram[199][0] ), .S0(n6268), .S1(n6134), .Y(n4690) );
  MX4X1 U7017 ( .A(n4681), .B(n4679), .C(n4680), .D(n4678), .S0(n6040), .S1(
        n6062), .Y(n4682) );
  MX4X1 U7018 ( .A(\ram[224][0] ), .B(\ram[225][0] ), .C(\ram[226][0] ), .D(
        \ram[227][0] ), .S0(n6268), .S1(n6134), .Y(n4681) );
  MX4X1 U7019 ( .A(\ram[232][0] ), .B(\ram[233][0] ), .C(\ram[234][0] ), .D(
        \ram[235][0] ), .S0(n6268), .S1(n6134), .Y(n4679) );
  MX4X1 U7020 ( .A(\ram[228][0] ), .B(\ram[229][0] ), .C(\ram[230][0] ), .D(
        \ram[231][0] ), .S0(n6268), .S1(n6134), .Y(n4680) );
  MX4X1 U7021 ( .A(\ram[252][0] ), .B(\ram[253][0] ), .C(\ram[254][0] ), .D(
        \ram[255][0] ), .S0(n6267), .S1(n6133), .Y(n571) );
  MX4X1 U7022 ( .A(n578), .B(n573), .C(n576), .D(n571), .S0(n6036), .S1(n6058), 
        .Y(n580) );
  MX4X1 U7023 ( .A(\ram[240][0] ), .B(\ram[241][0] ), .C(\ram[242][0] ), .D(
        \ram[243][0] ), .S0(n6267), .S1(n6133), .Y(n578) );
  MX4X1 U7024 ( .A(\ram[248][0] ), .B(\ram[249][0] ), .C(\ram[250][0] ), .D(
        \ram[251][0] ), .S0(n6267), .S1(n6133), .Y(n573) );
  MX4X1 U7025 ( .A(\ram[244][0] ), .B(\ram[245][0] ), .C(\ram[246][0] ), .D(
        \ram[247][0] ), .S0(n6267), .S1(n6133), .Y(n576) );
  NOR2X1 U7026 ( .A(N24), .B(N25), .Y(n71) );
  NOR2X1 U7027 ( .A(n7017), .B(N25), .Y(n208) );
  AND2X2 U7028 ( .A(N25), .B(n7017), .Y(n341) );
  AND2X2 U7029 ( .A(N25), .B(N24), .Y(n474) );
  NAND2X1 U7030 ( .A(mem_write_data[0]), .B(n6991), .Y(n7) );
  NAND2X1 U7031 ( .A(mem_write_data[1]), .B(n6991), .Y(n9) );
  NAND2X1 U7032 ( .A(mem_write_data[2]), .B(n6991), .Y(n10) );
  NAND2X1 U7033 ( .A(mem_write_data[3]), .B(n6991), .Y(n11) );
  INVX1 U7034 ( .A(N24), .Y(n7017) );
endmodule


module MEM_stage ( clk, rst, pipeline_reg_in, pipeline_reg_out, mem_op_dest );
  input [37:0] pipeline_reg_in;
  output [36:0] pipeline_reg_out;
  output [2:0] mem_op_dest;
  input clk, rst;
  wire   pipeline_reg_in_0, \pipeline_reg_in[3] , \pipeline_reg_in[2] ,
         \pipeline_reg_in[1] , n38, n39, n40, n41, n42, n43, n44;
  wire   [15:0] mem_read_data;
  assign pipeline_reg_in_0 = pipeline_reg_in[0];
  assign mem_op_dest[2] = \pipeline_reg_in[3] ;
  assign \pipeline_reg_in[3]  = pipeline_reg_in[3];
  assign mem_op_dest[1] = \pipeline_reg_in[2] ;
  assign \pipeline_reg_in[2]  = pipeline_reg_in[2];
  assign mem_op_dest[0] = \pipeline_reg_in[1] ;
  assign \pipeline_reg_in[1]  = pipeline_reg_in[1];

  data_mem dmem ( .clk(clk), .mem_access_addr({pipeline_reg_in[37:25], n42, 
        pipeline_reg_in[23], n40}), .mem_write_data(pipeline_reg_in[20:5]), 
        .mem_write_en(n38), .mem_read_data(mem_read_data) );
  DFFTRX2 \pipeline_reg_out_reg[4]  ( .D(pipeline_reg_in[4]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[4]) );
  DFFTRXL \pipeline_reg_out_reg[0]  ( .D(pipeline_reg_in_0), .RN(n44), .CK(clk), .Q(pipeline_reg_out[0]) );
  DFFTRXL \pipeline_reg_out_reg[36]  ( .D(pipeline_reg_in[37]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[36]) );
  DFFTRXL \pipeline_reg_out_reg[35]  ( .D(pipeline_reg_in[36]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[35]) );
  DFFTRXL \pipeline_reg_out_reg[34]  ( .D(pipeline_reg_in[35]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[34]) );
  DFFTRXL \pipeline_reg_out_reg[33]  ( .D(pipeline_reg_in[34]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[33]) );
  DFFTRXL \pipeline_reg_out_reg[32]  ( .D(pipeline_reg_in[33]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[32]) );
  DFFTRXL \pipeline_reg_out_reg[31]  ( .D(pipeline_reg_in[32]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[31]) );
  DFFTRXL \pipeline_reg_out_reg[30]  ( .D(pipeline_reg_in[31]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[30]) );
  DFFTRXL \pipeline_reg_out_reg[29]  ( .D(pipeline_reg_in[30]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[29]) );
  DFFTRXL \pipeline_reg_out_reg[28]  ( .D(pipeline_reg_in[29]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[28]) );
  DFFTRXL \pipeline_reg_out_reg[27]  ( .D(pipeline_reg_in[28]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[27]) );
  DFFTRXL \pipeline_reg_out_reg[26]  ( .D(pipeline_reg_in[27]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[26]) );
  DFFTRXL \pipeline_reg_out_reg[25]  ( .D(pipeline_reg_in[26]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[25]) );
  DFFTRXL \pipeline_reg_out_reg[24]  ( .D(pipeline_reg_in[25]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[24]) );
  DFFTRXL \pipeline_reg_out_reg[23]  ( .D(n42), .RN(n44), .CK(clk), .Q(
        pipeline_reg_out[23]) );
  DFFTRXL \pipeline_reg_out_reg[22]  ( .D(pipeline_reg_in[23]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[22]) );
  DFFTRXL \pipeline_reg_out_reg[21]  ( .D(n40), .RN(n44), .CK(clk), .Q(
        pipeline_reg_out[21]) );
  DFFTRXL \pipeline_reg_out_reg[20]  ( .D(mem_read_data[15]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[20]) );
  DFFTRXL \pipeline_reg_out_reg[5]  ( .D(mem_read_data[0]), .RN(n44), .CK(clk), 
        .Q(pipeline_reg_out[5]) );
  DFFTRXL \pipeline_reg_out_reg[7]  ( .D(mem_read_data[2]), .RN(n44), .CK(clk), 
        .Q(pipeline_reg_out[7]) );
  DFFTRXL \pipeline_reg_out_reg[6]  ( .D(mem_read_data[1]), .RN(n44), .CK(clk), 
        .Q(pipeline_reg_out[6]) );
  DFFTRXL \pipeline_reg_out_reg[19]  ( .D(mem_read_data[14]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[19]) );
  DFFTRXL \pipeline_reg_out_reg[18]  ( .D(mem_read_data[13]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[18]) );
  DFFTRXL \pipeline_reg_out_reg[17]  ( .D(mem_read_data[12]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[17]) );
  DFFTRXL \pipeline_reg_out_reg[16]  ( .D(mem_read_data[11]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[16]) );
  DFFTRXL \pipeline_reg_out_reg[8]  ( .D(mem_read_data[3]), .RN(n44), .CK(clk), 
        .Q(pipeline_reg_out[8]) );
  DFFTRXL \pipeline_reg_out_reg[15]  ( .D(mem_read_data[10]), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[15]) );
  DFFTRXL \pipeline_reg_out_reg[14]  ( .D(mem_read_data[9]), .RN(n44), .CK(clk), .Q(pipeline_reg_out[14]) );
  DFFTRXL \pipeline_reg_out_reg[13]  ( .D(mem_read_data[8]), .RN(n44), .CK(clk), .Q(pipeline_reg_out[13]) );
  DFFTRXL \pipeline_reg_out_reg[12]  ( .D(mem_read_data[7]), .RN(n44), .CK(clk), .Q(pipeline_reg_out[12]) );
  DFFTRXL \pipeline_reg_out_reg[11]  ( .D(mem_read_data[6]), .RN(n44), .CK(clk), .Q(pipeline_reg_out[11]) );
  DFFTRXL \pipeline_reg_out_reg[10]  ( .D(mem_read_data[5]), .RN(n44), .CK(clk), .Q(pipeline_reg_out[10]) );
  DFFTRXL \pipeline_reg_out_reg[9]  ( .D(mem_read_data[4]), .RN(n44), .CK(clk), 
        .Q(pipeline_reg_out[9]) );
  DFFTRX1 \pipeline_reg_out_reg[3]  ( .D(\pipeline_reg_in[3] ), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[3]) );
  DFFTRX1 \pipeline_reg_out_reg[1]  ( .D(\pipeline_reg_in[1] ), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[1]) );
  DFFTRX1 \pipeline_reg_out_reg[2]  ( .D(\pipeline_reg_in[2] ), .RN(n44), .CK(
        clk), .Q(pipeline_reg_out[2]) );
  INVX8 U3 ( .A(rst), .Y(n44) );
  INVX1 U4 ( .A(n39), .Y(n38) );
  INVX1 U5 ( .A(pipeline_reg_in[21]), .Y(n39) );
  INVX1 U6 ( .A(n41), .Y(n40) );
  INVX1 U7 ( .A(pipeline_reg_in[22]), .Y(n41) );
  INVX1 U8 ( .A(n43), .Y(n42) );
  INVX1 U9 ( .A(pipeline_reg_in[24]), .Y(n43) );
endmodule


module WB_stage ( pipeline_reg_in, reg_write_en, reg_write_dest, 
        reg_write_data, wb_op_dest );
  input [36:0] pipeline_reg_in;
  output [2:0] reg_write_dest;
  output [15:0] reg_write_data;
  output [2:0] wb_op_dest;
  output reg_write_en;
  wire   pipeline_reg_in_0, \pipeline_reg_in[3] , \pipeline_reg_in[2] ,
         \pipeline_reg_in[1] , n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n1, n2, n35;
  assign reg_write_en = pipeline_reg_in[4];
  assign pipeline_reg_in_0 = pipeline_reg_in[0];
  assign wb_op_dest[2] = \pipeline_reg_in[3] ;
  assign reg_write_dest[2] = \pipeline_reg_in[3] ;
  assign \pipeline_reg_in[3]  = pipeline_reg_in[3];
  assign wb_op_dest[1] = \pipeline_reg_in[2] ;
  assign reg_write_dest[1] = \pipeline_reg_in[2] ;
  assign \pipeline_reg_in[2]  = pipeline_reg_in[2];
  assign wb_op_dest[0] = \pipeline_reg_in[1] ;
  assign reg_write_dest[0] = \pipeline_reg_in[1] ;
  assign \pipeline_reg_in[1]  = pipeline_reg_in[1];

  BUFX3 U1 ( .A(pipeline_reg_in_0), .Y(n2) );
  BUFX3 U2 ( .A(n35), .Y(n1) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n34), .Y(reg_write_data[0]) );
  AOI22X1 U5 ( .A0(pipeline_reg_in[21]), .A1(n1), .B0(pipeline_reg_in[5]), 
        .B1(n2), .Y(n34) );
  INVX1 U6 ( .A(n27), .Y(reg_write_data[1]) );
  AOI22X1 U7 ( .A0(pipeline_reg_in[22]), .A1(n1), .B0(pipeline_reg_in[6]), 
        .B1(n2), .Y(n27) );
  INVX1 U8 ( .A(n26), .Y(reg_write_data[2]) );
  AOI22X1 U9 ( .A0(pipeline_reg_in[23]), .A1(n1), .B0(pipeline_reg_in[7]), 
        .B1(n2), .Y(n26) );
  INVX1 U10 ( .A(n25), .Y(reg_write_data[3]) );
  AOI22X1 U11 ( .A0(pipeline_reg_in[24]), .A1(n1), .B0(pipeline_reg_in[8]), 
        .B1(n2), .Y(n25) );
  INVX1 U12 ( .A(n24), .Y(reg_write_data[4]) );
  AOI22X1 U13 ( .A0(pipeline_reg_in[25]), .A1(n1), .B0(pipeline_reg_in[9]), 
        .B1(n2), .Y(n24) );
  INVX1 U14 ( .A(n23), .Y(reg_write_data[5]) );
  AOI22X1 U15 ( .A0(pipeline_reg_in[10]), .A1(n2), .B0(pipeline_reg_in[26]), 
        .B1(n1), .Y(n23) );
  INVX1 U16 ( .A(n22), .Y(reg_write_data[6]) );
  AOI22X1 U17 ( .A0(pipeline_reg_in[11]), .A1(n2), .B0(pipeline_reg_in[27]), 
        .B1(n1), .Y(n22) );
  INVX1 U18 ( .A(n21), .Y(reg_write_data[7]) );
  AOI22X1 U19 ( .A0(pipeline_reg_in[12]), .A1(n2), .B0(pipeline_reg_in[28]), 
        .B1(n1), .Y(n21) );
  INVX1 U20 ( .A(n20), .Y(reg_write_data[8]) );
  AOI22X1 U21 ( .A0(pipeline_reg_in[13]), .A1(n2), .B0(pipeline_reg_in[29]), 
        .B1(n1), .Y(n20) );
  INVX1 U22 ( .A(n19), .Y(reg_write_data[9]) );
  AOI22X1 U23 ( .A0(n2), .A1(pipeline_reg_in[14]), .B0(pipeline_reg_in[30]), 
        .B1(n1), .Y(n19) );
  INVX1 U24 ( .A(n33), .Y(reg_write_data[10]) );
  AOI22X1 U25 ( .A0(pipeline_reg_in[15]), .A1(n2), .B0(pipeline_reg_in[31]), 
        .B1(n1), .Y(n33) );
  INVX1 U26 ( .A(n32), .Y(reg_write_data[11]) );
  AOI22X1 U27 ( .A0(pipeline_reg_in[16]), .A1(n2), .B0(pipeline_reg_in[32]), 
        .B1(n1), .Y(n32) );
  INVX1 U28 ( .A(n31), .Y(reg_write_data[12]) );
  AOI22X1 U29 ( .A0(pipeline_reg_in[17]), .A1(n2), .B0(pipeline_reg_in[33]), 
        .B1(n1), .Y(n31) );
  INVX1 U30 ( .A(n30), .Y(reg_write_data[13]) );
  AOI22X1 U31 ( .A0(pipeline_reg_in[18]), .A1(n2), .B0(pipeline_reg_in[34]), 
        .B1(n1), .Y(n30) );
  INVX1 U32 ( .A(n29), .Y(reg_write_data[14]) );
  AOI22X1 U33 ( .A0(pipeline_reg_in[19]), .A1(n2), .B0(pipeline_reg_in[35]), 
        .B1(n1), .Y(n29) );
  INVX1 U34 ( .A(n28), .Y(reg_write_data[15]) );
  AOI22X1 U35 ( .A0(pipeline_reg_in[20]), .A1(n2), .B0(pipeline_reg_in[36]), 
        .B1(n1), .Y(n28) );
endmodule


module register_file ( clk, rst, reg_write_en, reg_write_dest, reg_write_data, 
        reg_read_addr_1, reg_read_data_1, reg_read_addr_2, reg_read_data_2 );
  input [2:0] reg_write_dest;
  input [15:0] reg_write_data;
  input [2:0] reg_read_addr_1;
  output [15:0] reg_read_data_1;
  input [2:0] reg_read_addr_2;
  output [15:0] reg_read_data_2;
  input clk, rst, reg_write_en;
  wire   N18, N19, N20, N21, N22, N23, \reg_array[7][15] , \reg_array[7][14] ,
         \reg_array[7][13] , \reg_array[7][12] , \reg_array[7][11] ,
         \reg_array[7][10] , \reg_array[7][9] , \reg_array[7][8] ,
         \reg_array[7][7] , \reg_array[7][6] , \reg_array[7][5] ,
         \reg_array[7][4] , \reg_array[7][3] , \reg_array[7][2] ,
         \reg_array[7][1] , \reg_array[7][0] , \reg_array[6][15] ,
         \reg_array[6][14] , \reg_array[6][13] , \reg_array[6][12] ,
         \reg_array[6][11] , \reg_array[6][10] , \reg_array[6][9] ,
         \reg_array[6][8] , \reg_array[6][7] , \reg_array[6][6] ,
         \reg_array[6][5] , \reg_array[6][4] , \reg_array[6][3] ,
         \reg_array[6][2] , \reg_array[6][1] , \reg_array[6][0] ,
         \reg_array[5][15] , \reg_array[5][14] , \reg_array[5][13] ,
         \reg_array[5][12] , \reg_array[5][11] , \reg_array[5][10] ,
         \reg_array[5][9] , \reg_array[5][8] , \reg_array[5][7] ,
         \reg_array[5][6] , \reg_array[5][5] , \reg_array[5][4] ,
         \reg_array[5][3] , \reg_array[5][2] , \reg_array[5][1] ,
         \reg_array[5][0] , \reg_array[4][15] , \reg_array[4][14] ,
         \reg_array[4][13] , \reg_array[4][12] , \reg_array[4][11] ,
         \reg_array[4][10] , \reg_array[4][9] , \reg_array[4][8] ,
         \reg_array[4][7] , \reg_array[4][6] , \reg_array[4][5] ,
         \reg_array[4][4] , \reg_array[4][3] , \reg_array[4][2] ,
         \reg_array[4][1] , \reg_array[4][0] , \reg_array[3][15] ,
         \reg_array[3][14] , \reg_array[3][13] , \reg_array[3][12] ,
         \reg_array[3][11] , \reg_array[3][10] , \reg_array[3][9] ,
         \reg_array[3][8] , \reg_array[3][7] , \reg_array[3][6] ,
         \reg_array[3][5] , \reg_array[3][4] , \reg_array[3][3] ,
         \reg_array[3][2] , \reg_array[3][1] , \reg_array[3][0] ,
         \reg_array[2][15] , \reg_array[2][14] , \reg_array[2][13] ,
         \reg_array[2][12] , \reg_array[2][11] , \reg_array[2][10] ,
         \reg_array[2][9] , \reg_array[2][8] , \reg_array[2][7] ,
         \reg_array[2][6] , \reg_array[2][5] , \reg_array[2][4] ,
         \reg_array[2][3] , \reg_array[2][2] , \reg_array[2][1] ,
         \reg_array[2][0] , \reg_array[1][15] , \reg_array[1][14] ,
         \reg_array[1][13] , \reg_array[1][12] , \reg_array[1][11] ,
         \reg_array[1][10] , \reg_array[1][9] , \reg_array[1][8] ,
         \reg_array[1][7] , \reg_array[1][6] , \reg_array[1][5] ,
         \reg_array[1][4] , \reg_array[1][3] , \reg_array[1][2] ,
         \reg_array[1][1] , \reg_array[1][0] , \reg_array[0][15] ,
         \reg_array[0][14] , \reg_array[0][13] , \reg_array[0][12] ,
         \reg_array[0][11] , \reg_array[0][10] , \reg_array[0][9] ,
         \reg_array[0][8] , \reg_array[0][7] , \reg_array[0][6] ,
         \reg_array[0][5] , \reg_array[0][4] , \reg_array[0][3] ,
         \reg_array[0][2] , \reg_array[0][1] , \reg_array[0][0] , N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, n24, n27, n28, n29,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26,
         n30, n31, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263;
  assign N18 = reg_read_addr_1[0];
  assign N19 = reg_read_addr_1[1];
  assign N20 = reg_read_addr_1[2];
  assign N21 = reg_read_addr_2[0];
  assign N22 = reg_read_addr_2[1];
  assign N23 = reg_read_addr_2[2];

  DFFRHQX1 \reg_array_reg[5][15]  ( .D(n127), .CK(clk), .RN(n220), .Q(
        \reg_array[5][15] ) );
  DFFRHQX1 \reg_array_reg[5][14]  ( .D(n126), .CK(clk), .RN(n222), .Q(
        \reg_array[5][14] ) );
  DFFRHQX1 \reg_array_reg[5][13]  ( .D(n125), .CK(clk), .RN(n220), .Q(
        \reg_array[5][13] ) );
  DFFRHQX1 \reg_array_reg[5][12]  ( .D(n124), .CK(clk), .RN(n218), .Q(
        \reg_array[5][12] ) );
  DFFRHQX1 \reg_array_reg[5][11]  ( .D(n123), .CK(clk), .RN(n218), .Q(
        \reg_array[5][11] ) );
  DFFRHQX1 \reg_array_reg[5][10]  ( .D(n122), .CK(clk), .RN(n222), .Q(
        \reg_array[5][10] ) );
  DFFRHQX1 \reg_array_reg[5][9]  ( .D(n121), .CK(clk), .RN(n220), .Q(
        \reg_array[5][9] ) );
  DFFRHQX1 \reg_array_reg[5][8]  ( .D(n120), .CK(clk), .RN(n218), .Q(
        \reg_array[5][8] ) );
  DFFRHQX1 \reg_array_reg[5][7]  ( .D(n119), .CK(clk), .RN(n217), .Q(
        \reg_array[5][7] ) );
  DFFRHQX1 \reg_array_reg[5][6]  ( .D(n118), .CK(clk), .RN(n222), .Q(
        \reg_array[5][6] ) );
  DFFRHQX1 \reg_array_reg[5][5]  ( .D(n117), .CK(clk), .RN(n220), .Q(
        \reg_array[5][5] ) );
  DFFRHQX1 \reg_array_reg[5][4]  ( .D(n116), .CK(clk), .RN(n216), .Q(
        \reg_array[5][4] ) );
  DFFRHQX1 \reg_array_reg[5][3]  ( .D(n115), .CK(clk), .RN(n221), .Q(
        \reg_array[5][3] ) );
  DFFRHQX1 \reg_array_reg[5][2]  ( .D(n114), .CK(clk), .RN(n221), .Q(
        \reg_array[5][2] ) );
  DFFRHQX1 \reg_array_reg[5][1]  ( .D(n113), .CK(clk), .RN(n221), .Q(
        \reg_array[5][1] ) );
  DFFRHQX1 \reg_array_reg[5][0]  ( .D(n112), .CK(clk), .RN(n221), .Q(
        \reg_array[5][0] ) );
  DFFRHQX1 \reg_array_reg[1][15]  ( .D(n63), .CK(clk), .RN(n218), .Q(
        \reg_array[1][15] ) );
  DFFRHQX1 \reg_array_reg[1][14]  ( .D(n62), .CK(clk), .RN(n218), .Q(
        \reg_array[1][14] ) );
  DFFRHQX1 \reg_array_reg[1][13]  ( .D(n61), .CK(clk), .RN(n218), .Q(
        \reg_array[1][13] ) );
  DFFRHQX1 \reg_array_reg[1][12]  ( .D(n60), .CK(clk), .RN(n218), .Q(
        \reg_array[1][12] ) );
  DFFRHQX1 \reg_array_reg[1][11]  ( .D(n59), .CK(clk), .RN(n218), .Q(
        \reg_array[1][11] ) );
  DFFRHQX1 \reg_array_reg[1][10]  ( .D(n58), .CK(clk), .RN(n218), .Q(
        \reg_array[1][10] ) );
  DFFRHQX1 \reg_array_reg[1][9]  ( .D(n57), .CK(clk), .RN(n218), .Q(
        \reg_array[1][9] ) );
  DFFRHQX1 \reg_array_reg[1][8]  ( .D(n56), .CK(clk), .RN(n218), .Q(
        \reg_array[1][8] ) );
  DFFRHQX1 \reg_array_reg[1][7]  ( .D(n55), .CK(clk), .RN(n217), .Q(
        \reg_array[1][7] ) );
  DFFRHQX1 \reg_array_reg[1][6]  ( .D(n54), .CK(clk), .RN(n217), .Q(
        \reg_array[1][6] ) );
  DFFRHQX1 \reg_array_reg[1][5]  ( .D(n53), .CK(clk), .RN(n217), .Q(
        \reg_array[1][5] ) );
  DFFRHQX1 \reg_array_reg[1][4]  ( .D(n52), .CK(clk), .RN(n217), .Q(
        \reg_array[1][4] ) );
  DFFRHQX1 \reg_array_reg[1][3]  ( .D(n51), .CK(clk), .RN(n217), .Q(
        \reg_array[1][3] ) );
  DFFRHQX1 \reg_array_reg[1][2]  ( .D(n50), .CK(clk), .RN(n217), .Q(
        \reg_array[1][2] ) );
  DFFRHQX1 \reg_array_reg[1][1]  ( .D(n49), .CK(clk), .RN(n217), .Q(
        \reg_array[1][1] ) );
  DFFRHQX1 \reg_array_reg[1][0]  ( .D(n48), .CK(clk), .RN(n217), .Q(
        \reg_array[1][0] ) );
  DFFRHQX1 \reg_array_reg[7][15]  ( .D(n159), .CK(clk), .RN(n219), .Q(
        \reg_array[7][15] ) );
  DFFRHQX1 \reg_array_reg[7][14]  ( .D(n158), .CK(clk), .RN(n218), .Q(
        \reg_array[7][14] ) );
  DFFRHQX1 \reg_array_reg[7][13]  ( .D(n157), .CK(clk), .RN(n217), .Q(
        \reg_array[7][13] ) );
  DFFRHQX1 \reg_array_reg[7][12]  ( .D(n156), .CK(clk), .RN(n221), .Q(
        \reg_array[7][12] ) );
  DFFRHQX1 \reg_array_reg[7][11]  ( .D(n155), .CK(clk), .RN(n216), .Q(
        \reg_array[7][11] ) );
  DFFRHQX1 \reg_array_reg[7][10]  ( .D(n154), .CK(clk), .RN(n216), .Q(
        \reg_array[7][10] ) );
  DFFRHQX1 \reg_array_reg[7][9]  ( .D(n153), .CK(clk), .RN(n216), .Q(
        \reg_array[7][9] ) );
  DFFRHQX1 \reg_array_reg[7][8]  ( .D(n152), .CK(clk), .RN(n216), .Q(
        \reg_array[7][8] ) );
  DFFRHQX1 \reg_array_reg[7][7]  ( .D(n151), .CK(clk), .RN(n222), .Q(
        \reg_array[7][7] ) );
  DFFRHQX1 \reg_array_reg[7][6]  ( .D(n150), .CK(clk), .RN(n220), .Q(
        \reg_array[7][6] ) );
  DFFRHQX1 \reg_array_reg[7][5]  ( .D(n149), .CK(clk), .RN(n218), .Q(
        \reg_array[7][5] ) );
  DFFRHQX1 \reg_array_reg[7][4]  ( .D(n148), .CK(clk), .RN(n219), .Q(
        \reg_array[7][4] ) );
  DFFRHQX1 \reg_array_reg[7][3]  ( .D(n147), .CK(clk), .RN(n219), .Q(
        \reg_array[7][3] ) );
  DFFRHQX1 \reg_array_reg[7][2]  ( .D(n146), .CK(clk), .RN(n217), .Q(
        \reg_array[7][2] ) );
  DFFRHQX1 \reg_array_reg[7][1]  ( .D(n145), .CK(clk), .RN(n221), .Q(
        \reg_array[7][1] ) );
  DFFRHQX1 \reg_array_reg[7][0]  ( .D(n144), .CK(clk), .RN(n219), .Q(
        \reg_array[7][0] ) );
  DFFRHQX1 \reg_array_reg[3][15]  ( .D(n95), .CK(clk), .RN(n222), .Q(
        \reg_array[3][15] ) );
  DFFRHQX1 \reg_array_reg[3][14]  ( .D(n94), .CK(clk), .RN(n220), .Q(
        \reg_array[3][14] ) );
  DFFRHQX1 \reg_array_reg[3][13]  ( .D(n93), .CK(clk), .RN(n218), .Q(
        \reg_array[3][13] ) );
  DFFRHQX1 \reg_array_reg[3][12]  ( .D(n92), .CK(clk), .RN(n217), .Q(
        \reg_array[3][12] ) );
  DFFRHQX1 \reg_array_reg[3][11]  ( .D(n91), .CK(clk), .RN(n220), .Q(
        \reg_array[3][11] ) );
  DFFRHQX1 \reg_array_reg[3][10]  ( .D(n90), .CK(clk), .RN(n220), .Q(
        \reg_array[3][10] ) );
  DFFRHQX1 \reg_array_reg[3][9]  ( .D(n89), .CK(clk), .RN(n220), .Q(
        \reg_array[3][9] ) );
  DFFRHQX1 \reg_array_reg[3][8]  ( .D(n88), .CK(clk), .RN(n220), .Q(
        \reg_array[3][8] ) );
  DFFRHQX1 \reg_array_reg[3][7]  ( .D(n87), .CK(clk), .RN(n220), .Q(
        \reg_array[3][7] ) );
  DFFRHQX1 \reg_array_reg[3][6]  ( .D(n86), .CK(clk), .RN(n220), .Q(
        \reg_array[3][6] ) );
  DFFRHQX1 \reg_array_reg[3][5]  ( .D(n85), .CK(clk), .RN(n220), .Q(
        \reg_array[3][5] ) );
  DFFRHQX1 \reg_array_reg[3][4]  ( .D(n84), .CK(clk), .RN(n220), .Q(
        \reg_array[3][4] ) );
  DFFRHQX1 \reg_array_reg[3][3]  ( .D(n83), .CK(clk), .RN(n220), .Q(
        \reg_array[3][3] ) );
  DFFRHQX1 \reg_array_reg[3][2]  ( .D(n82), .CK(clk), .RN(n220), .Q(
        \reg_array[3][2] ) );
  DFFRHQX1 \reg_array_reg[3][1]  ( .D(n81), .CK(clk), .RN(n220), .Q(
        \reg_array[3][1] ) );
  DFFRHQX1 \reg_array_reg[3][0]  ( .D(n80), .CK(clk), .RN(n220), .Q(
        \reg_array[3][0] ) );
  DFFRHQX1 \reg_array_reg[4][15]  ( .D(n111), .CK(clk), .RN(n221), .Q(
        \reg_array[4][15] ) );
  DFFRHQX1 \reg_array_reg[4][14]  ( .D(n110), .CK(clk), .RN(n221), .Q(
        \reg_array[4][14] ) );
  DFFRHQX1 \reg_array_reg[4][13]  ( .D(n109), .CK(clk), .RN(n221), .Q(
        \reg_array[4][13] ) );
  DFFRHQX1 \reg_array_reg[4][12]  ( .D(n108), .CK(clk), .RN(n221), .Q(
        \reg_array[4][12] ) );
  DFFRHQX1 \reg_array_reg[4][11]  ( .D(n107), .CK(clk), .RN(n221), .Q(
        \reg_array[4][11] ) );
  DFFRHQX1 \reg_array_reg[4][10]  ( .D(n106), .CK(clk), .RN(n221), .Q(
        \reg_array[4][10] ) );
  DFFRHQX1 \reg_array_reg[4][9]  ( .D(n105), .CK(clk), .RN(n221), .Q(
        \reg_array[4][9] ) );
  DFFRHQX1 \reg_array_reg[4][8]  ( .D(n104), .CK(clk), .RN(n221), .Q(
        \reg_array[4][8] ) );
  DFFRHQX1 \reg_array_reg[4][7]  ( .D(n103), .CK(clk), .RN(n221), .Q(
        \reg_array[4][7] ) );
  DFFRHQX1 \reg_array_reg[4][6]  ( .D(n102), .CK(clk), .RN(n221), .Q(
        \reg_array[4][6] ) );
  DFFRHQX1 \reg_array_reg[4][5]  ( .D(n101), .CK(clk), .RN(n217), .Q(
        \reg_array[4][5] ) );
  DFFRHQX1 \reg_array_reg[4][4]  ( .D(n100), .CK(clk), .RN(n221), .Q(
        \reg_array[4][4] ) );
  DFFRHQX1 \reg_array_reg[4][3]  ( .D(n99), .CK(clk), .RN(n216), .Q(
        \reg_array[4][3] ) );
  DFFRHQX1 \reg_array_reg[4][2]  ( .D(n98), .CK(clk), .RN(n219), .Q(
        \reg_array[4][2] ) );
  DFFRHQX1 \reg_array_reg[4][1]  ( .D(n97), .CK(clk), .RN(n219), .Q(
        \reg_array[4][1] ) );
  DFFRHQX1 \reg_array_reg[4][0]  ( .D(n96), .CK(clk), .RN(n219), .Q(
        \reg_array[4][0] ) );
  DFFRHQX1 \reg_array_reg[0][15]  ( .D(n47), .CK(clk), .RN(n217), .Q(
        \reg_array[0][15] ) );
  DFFRHQX1 \reg_array_reg[0][14]  ( .D(n46), .CK(clk), .RN(n217), .Q(
        \reg_array[0][14] ) );
  DFFRHQX1 \reg_array_reg[0][13]  ( .D(n45), .CK(clk), .RN(n217), .Q(
        \reg_array[0][13] ) );
  DFFRHQX1 \reg_array_reg[0][12]  ( .D(n44), .CK(clk), .RN(n217), .Q(
        \reg_array[0][12] ) );
  DFFRHQX1 \reg_array_reg[0][11]  ( .D(n43), .CK(clk), .RN(n221), .Q(
        \reg_array[0][11] ) );
  DFFRHQX1 \reg_array_reg[0][10]  ( .D(n42), .CK(clk), .RN(n222), .Q(
        \reg_array[0][10] ) );
  DFFRHQX1 \reg_array_reg[0][9]  ( .D(n41), .CK(clk), .RN(n220), .Q(
        \reg_array[0][9] ) );
  DFFRHQX1 \reg_array_reg[0][8]  ( .D(n40), .CK(clk), .RN(n218), .Q(
        \reg_array[0][8] ) );
  DFFRHQX1 \reg_array_reg[0][7]  ( .D(n39), .CK(clk), .RN(n217), .Q(
        \reg_array[0][7] ) );
  DFFRHQX1 \reg_array_reg[0][6]  ( .D(n38), .CK(clk), .RN(n221), .Q(
        \reg_array[0][6] ) );
  DFFRHQX1 \reg_array_reg[0][5]  ( .D(n37), .CK(clk), .RN(n222), .Q(
        \reg_array[0][5] ) );
  DFFRHQX1 \reg_array_reg[0][4]  ( .D(n36), .CK(clk), .RN(n220), .Q(
        \reg_array[0][4] ) );
  DFFRHQX1 \reg_array_reg[0][3]  ( .D(n35), .CK(clk), .RN(n218), .Q(
        \reg_array[0][3] ) );
  DFFRHQX1 \reg_array_reg[0][2]  ( .D(n34), .CK(clk), .RN(n217), .Q(
        \reg_array[0][2] ) );
  DFFRHQX1 \reg_array_reg[0][1]  ( .D(n33), .CK(clk), .RN(n221), .Q(
        \reg_array[0][1] ) );
  DFFRHQX1 \reg_array_reg[0][0]  ( .D(n32), .CK(clk), .RN(n222), .Q(
        \reg_array[0][0] ) );
  DFFRHQX1 \reg_array_reg[6][15]  ( .D(n143), .CK(clk), .RN(n219), .Q(
        \reg_array[6][15] ) );
  DFFRHQX1 \reg_array_reg[6][14]  ( .D(n142), .CK(clk), .RN(n217), .Q(
        \reg_array[6][14] ) );
  DFFRHQX1 \reg_array_reg[6][13]  ( .D(n141), .CK(clk), .RN(n221), .Q(
        \reg_array[6][13] ) );
  DFFRHQX1 \reg_array_reg[6][12]  ( .D(n140), .CK(clk), .RN(n219), .Q(
        \reg_array[6][12] ) );
  DFFRHQX1 \reg_array_reg[6][11]  ( .D(n139), .CK(clk), .RN(n222), .Q(
        \reg_array[6][11] ) );
  DFFRHQX1 \reg_array_reg[6][10]  ( .D(n138), .CK(clk), .RN(n222), .Q(
        \reg_array[6][10] ) );
  DFFRHQX1 \reg_array_reg[6][9]  ( .D(n137), .CK(clk), .RN(n222), .Q(
        \reg_array[6][9] ) );
  DFFRHQX1 \reg_array_reg[6][8]  ( .D(n136), .CK(clk), .RN(n222), .Q(
        \reg_array[6][8] ) );
  DFFRHQX1 \reg_array_reg[6][7]  ( .D(n135), .CK(clk), .RN(n222), .Q(
        \reg_array[6][7] ) );
  DFFRHQX1 \reg_array_reg[6][6]  ( .D(n134), .CK(clk), .RN(n222), .Q(
        \reg_array[6][6] ) );
  DFFRHQX1 \reg_array_reg[6][5]  ( .D(n133), .CK(clk), .RN(n222), .Q(
        \reg_array[6][5] ) );
  DFFRHQX1 \reg_array_reg[6][4]  ( .D(n132), .CK(clk), .RN(n222), .Q(
        \reg_array[6][4] ) );
  DFFRHQX1 \reg_array_reg[6][3]  ( .D(n131), .CK(clk), .RN(n222), .Q(
        \reg_array[6][3] ) );
  DFFRHQX1 \reg_array_reg[6][2]  ( .D(n130), .CK(clk), .RN(n222), .Q(
        \reg_array[6][2] ) );
  DFFRHQX1 \reg_array_reg[6][1]  ( .D(n129), .CK(clk), .RN(n222), .Q(
        \reg_array[6][1] ) );
  DFFRHQX1 \reg_array_reg[6][0]  ( .D(n128), .CK(clk), .RN(n222), .Q(
        \reg_array[6][0] ) );
  DFFRHQX1 \reg_array_reg[2][15]  ( .D(n79), .CK(clk), .RN(n219), .Q(
        \reg_array[2][15] ) );
  DFFRHQX1 \reg_array_reg[2][14]  ( .D(n78), .CK(clk), .RN(n219), .Q(
        \reg_array[2][14] ) );
  DFFRHQX1 \reg_array_reg[2][13]  ( .D(n77), .CK(clk), .RN(n219), .Q(
        \reg_array[2][13] ) );
  DFFRHQX1 \reg_array_reg[2][12]  ( .D(n76), .CK(clk), .RN(n219), .Q(
        \reg_array[2][12] ) );
  DFFRHQX1 \reg_array_reg[2][11]  ( .D(n75), .CK(clk), .RN(n219), .Q(
        \reg_array[2][11] ) );
  DFFRHQX1 \reg_array_reg[2][10]  ( .D(n74), .CK(clk), .RN(n219), .Q(
        \reg_array[2][10] ) );
  DFFRHQX1 \reg_array_reg[2][9]  ( .D(n73), .CK(clk), .RN(n219), .Q(
        \reg_array[2][9] ) );
  DFFRHQX1 \reg_array_reg[2][8]  ( .D(n72), .CK(clk), .RN(n219), .Q(
        \reg_array[2][8] ) );
  DFFRHQX1 \reg_array_reg[2][7]  ( .D(n71), .CK(clk), .RN(n219), .Q(
        \reg_array[2][7] ) );
  DFFRHQX1 \reg_array_reg[2][6]  ( .D(n70), .CK(clk), .RN(n219), .Q(
        \reg_array[2][6] ) );
  DFFRHQX1 \reg_array_reg[2][5]  ( .D(n69), .CK(clk), .RN(n219), .Q(
        \reg_array[2][5] ) );
  DFFRHQX1 \reg_array_reg[2][4]  ( .D(n68), .CK(clk), .RN(n219), .Q(
        \reg_array[2][4] ) );
  DFFRHQX1 \reg_array_reg[2][3]  ( .D(n67), .CK(clk), .RN(n218), .Q(
        \reg_array[2][3] ) );
  DFFRHQX1 \reg_array_reg[2][2]  ( .D(n66), .CK(clk), .RN(n218), .Q(
        \reg_array[2][2] ) );
  DFFRHQX1 \reg_array_reg[2][1]  ( .D(n65), .CK(clk), .RN(n218), .Q(
        \reg_array[2][1] ) );
  DFFRHQX1 \reg_array_reg[2][0]  ( .D(n64), .CK(clk), .RN(n218), .Q(
        \reg_array[2][0] ) );
  AND4X2 U2 ( .A(reg_write_dest[2]), .B(reg_write_dest[1]), .C(reg_write_en), 
        .D(n263), .Y(n1) );
  AND4X2 U3 ( .A(reg_write_dest[0]), .B(reg_write_en), .C(n262), .D(n261), .Y(
        n2) );
  AND4X2 U4 ( .A(reg_write_dest[1]), .B(reg_write_en), .C(n263), .D(n261), .Y(
        n3) );
  AND4X1 U5 ( .A(reg_write_dest[2]), .B(reg_write_dest[1]), .C(
        reg_write_dest[0]), .D(reg_write_en), .Y(n4) );
  OR3X4 U6 ( .A(N22), .B(N23), .C(N21), .Y(n5) );
  OR3X4 U7 ( .A(N19), .B(N20), .C(n175), .Y(n6) );
  NAND4X1 U8 ( .A(reg_write_dest[1]), .B(reg_write_dest[0]), .C(reg_write_en), 
        .D(n261), .Y(n27) );
  AND2X1 U9 ( .A(N166), .B(n6), .Y(reg_read_data_1[2]) );
  AND2X1 U10 ( .A(N167), .B(n6), .Y(reg_read_data_1[1]) );
  AND2X1 U11 ( .A(N165), .B(n6), .Y(reg_read_data_1[3]) );
  AND2X1 U12 ( .A(N153), .B(n6), .Y(reg_read_data_1[15]) );
  AND2X1 U13 ( .A(N164), .B(n6), .Y(reg_read_data_1[4]) );
  AND2X1 U14 ( .A(N162), .B(n6), .Y(reg_read_data_1[6]) );
  CLKINVX3 U15 ( .A(n214), .Y(n213) );
  CLKINVX3 U16 ( .A(n214), .Y(n212) );
  CLKINVX3 U17 ( .A(n209), .Y(n211) );
  CLKINVX3 U18 ( .A(n209), .Y(n210) );
  INVX1 U19 ( .A(N22), .Y(n209) );
  CLKINVX3 U20 ( .A(n244), .Y(n175) );
  CLKINVX3 U21 ( .A(n244), .Y(n174) );
  CLKINVX3 U22 ( .A(n171), .Y(n172) );
  INVX1 U23 ( .A(N21), .Y(n214) );
  CLKINVX3 U24 ( .A(n171), .Y(n173) );
  CLKINVX3 U25 ( .A(n223), .Y(n217) );
  CLKINVX3 U26 ( .A(n223), .Y(n218) );
  CLKINVX3 U27 ( .A(rst), .Y(n219) );
  CLKINVX3 U28 ( .A(n223), .Y(n220) );
  CLKINVX3 U29 ( .A(n223), .Y(n221) );
  CLKINVX3 U30 ( .A(n223), .Y(n222) );
  INVX1 U31 ( .A(N19), .Y(n171) );
  BUFX3 U32 ( .A(N23), .Y(n215) );
  CLKINVX3 U33 ( .A(n243), .Y(n241) );
  CLKINVX3 U34 ( .A(n2), .Y(n240) );
  CLKINVX3 U35 ( .A(n3), .Y(n238) );
  CLKINVX3 U36 ( .A(n236), .Y(n234) );
  CLKINVX3 U37 ( .A(n233), .Y(n231) );
  CLKINVX3 U38 ( .A(n230), .Y(n228) );
  CLKINVX3 U39 ( .A(n1), .Y(n227) );
  CLKINVX3 U40 ( .A(n4), .Y(n225) );
  INVX1 U41 ( .A(n243), .Y(n242) );
  INVX1 U42 ( .A(n236), .Y(n235) );
  INVX1 U43 ( .A(n233), .Y(n232) );
  INVX1 U44 ( .A(n230), .Y(n229) );
  INVX1 U45 ( .A(n216), .Y(n223) );
  CLKINVX3 U46 ( .A(n1), .Y(n226) );
  CLKINVX3 U47 ( .A(n4), .Y(n224) );
  INVX1 U48 ( .A(n24), .Y(n243) );
  INVX1 U49 ( .A(n28), .Y(n233) );
  INVX1 U50 ( .A(n27), .Y(n236) );
  INVX1 U51 ( .A(n29), .Y(n230) );
  CLKINVX3 U52 ( .A(n2), .Y(n239) );
  CLKINVX3 U53 ( .A(n3), .Y(n237) );
  INVX1 U54 ( .A(rst), .Y(n216) );
  AND2X1 U55 ( .A(N154), .B(n6), .Y(reg_read_data_1[14]) );
  MX2X1 U56 ( .A(n168), .B(n167), .S0(n176), .Y(N154) );
  MX4X1 U57 ( .A(\reg_array[0][14] ), .B(\reg_array[1][14] ), .C(
        \reg_array[2][14] ), .D(\reg_array[3][14] ), .S0(n174), .S1(n172), .Y(
        n168) );
  MX4X1 U58 ( .A(\reg_array[4][14] ), .B(\reg_array[5][14] ), .C(
        \reg_array[6][14] ), .D(\reg_array[7][14] ), .S0(n174), .S1(n172), .Y(
        n167) );
  AND2X2 U59 ( .A(N180), .B(n5), .Y(reg_read_data_2[4]) );
  MX2X1 U60 ( .A(n186), .B(n185), .S0(n215), .Y(N180) );
  MX4X1 U61 ( .A(\reg_array[0][4] ), .B(\reg_array[1][4] ), .C(
        \reg_array[2][4] ), .D(\reg_array[3][4] ), .S0(n213), .S1(n211), .Y(
        n186) );
  MX4X1 U62 ( .A(\reg_array[4][4] ), .B(\reg_array[5][4] ), .C(
        \reg_array[6][4] ), .D(\reg_array[7][4] ), .S0(n213), .S1(n211), .Y(
        n185) );
  AND2X1 U63 ( .A(N168), .B(n6), .Y(reg_read_data_1[0]) );
  MX2X1 U64 ( .A(n8), .B(n7), .S0(n176), .Y(N168) );
  MX4X1 U65 ( .A(\reg_array[0][0] ), .B(\reg_array[1][0] ), .C(
        \reg_array[2][0] ), .D(\reg_array[3][0] ), .S0(n174), .S1(n172), .Y(n8) );
  MX4X1 U66 ( .A(\reg_array[4][0] ), .B(\reg_array[5][0] ), .C(
        \reg_array[6][0] ), .D(\reg_array[7][0] ), .S0(n174), .S1(n172), .Y(n7) );
  AND2X1 U67 ( .A(N160), .B(n6), .Y(reg_read_data_1[8]) );
  MX2X1 U68 ( .A(n25), .B(n23), .S0(n176), .Y(N160) );
  MX4X1 U69 ( .A(\reg_array[0][8] ), .B(\reg_array[1][8] ), .C(
        \reg_array[2][8] ), .D(\reg_array[3][8] ), .S0(n175), .S1(n173), .Y(
        n25) );
  MX4X1 U70 ( .A(\reg_array[4][8] ), .B(\reg_array[5][8] ), .C(
        \reg_array[6][8] ), .D(\reg_array[7][8] ), .S0(n175), .S1(n173), .Y(
        n23) );
  AND2X1 U71 ( .A(N159), .B(n6), .Y(reg_read_data_1[9]) );
  MX2X1 U72 ( .A(n30), .B(n26), .S0(n176), .Y(N159) );
  MX4X1 U73 ( .A(\reg_array[0][9] ), .B(\reg_array[1][9] ), .C(
        \reg_array[2][9] ), .D(\reg_array[3][9] ), .S0(n175), .S1(n173), .Y(
        n30) );
  MX4X1 U74 ( .A(\reg_array[4][9] ), .B(\reg_array[5][9] ), .C(
        \reg_array[6][9] ), .D(\reg_array[7][9] ), .S0(n175), .S1(n173), .Y(
        n26) );
  AND2X1 U75 ( .A(N156), .B(n6), .Y(reg_read_data_1[12]) );
  MX2X1 U76 ( .A(n164), .B(n163), .S0(n176), .Y(N156) );
  MX4X1 U77 ( .A(\reg_array[0][12] ), .B(\reg_array[1][12] ), .C(
        \reg_array[2][12] ), .D(\reg_array[3][12] ), .S0(n175), .S1(n173), .Y(
        n164) );
  MX4X1 U78 ( .A(\reg_array[4][12] ), .B(\reg_array[5][12] ), .C(
        \reg_array[6][12] ), .D(\reg_array[7][12] ), .S0(n174), .S1(n172), .Y(
        n163) );
  AND2X1 U79 ( .A(N155), .B(n6), .Y(reg_read_data_1[13]) );
  MX2X1 U80 ( .A(n166), .B(n165), .S0(n176), .Y(N155) );
  MX4X1 U81 ( .A(\reg_array[0][13] ), .B(\reg_array[1][13] ), .C(
        \reg_array[2][13] ), .D(\reg_array[3][13] ), .S0(n174), .S1(n172), .Y(
        n166) );
  MX4X1 U82 ( .A(\reg_array[4][13] ), .B(\reg_array[5][13] ), .C(
        \reg_array[6][13] ), .D(\reg_array[7][13] ), .S0(n174), .S1(n172), .Y(
        n165) );
  AND2X2 U83 ( .A(N184), .B(n5), .Y(reg_read_data_2[0]) );
  MX2X1 U84 ( .A(n178), .B(n177), .S0(n215), .Y(N184) );
  MX4X1 U85 ( .A(\reg_array[0][0] ), .B(\reg_array[1][0] ), .C(
        \reg_array[2][0] ), .D(\reg_array[3][0] ), .S0(n212), .S1(n210), .Y(
        n178) );
  MX4X1 U86 ( .A(\reg_array[4][0] ), .B(\reg_array[5][0] ), .C(
        \reg_array[6][0] ), .D(\reg_array[7][0] ), .S0(n212), .S1(n210), .Y(
        n177) );
  AND2X2 U87 ( .A(N183), .B(n5), .Y(reg_read_data_2[1]) );
  MX2X1 U88 ( .A(n180), .B(n179), .S0(n215), .Y(N183) );
  MX4X1 U89 ( .A(\reg_array[0][1] ), .B(\reg_array[1][1] ), .C(
        \reg_array[2][1] ), .D(\reg_array[3][1] ), .S0(n212), .S1(n210), .Y(
        n180) );
  MX4X1 U90 ( .A(\reg_array[4][1] ), .B(\reg_array[5][1] ), .C(
        \reg_array[6][1] ), .D(\reg_array[7][1] ), .S0(n212), .S1(n210), .Y(
        n179) );
  AND2X2 U91 ( .A(N182), .B(n5), .Y(reg_read_data_2[2]) );
  MX2X1 U92 ( .A(n182), .B(n181), .S0(n215), .Y(N182) );
  MX4X1 U93 ( .A(\reg_array[0][2] ), .B(\reg_array[1][2] ), .C(
        \reg_array[2][2] ), .D(\reg_array[3][2] ), .S0(n212), .S1(n210), .Y(
        n182) );
  MX4X1 U94 ( .A(\reg_array[4][2] ), .B(\reg_array[5][2] ), .C(
        \reg_array[6][2] ), .D(\reg_array[7][2] ), .S0(n212), .S1(n210), .Y(
        n181) );
  AND2X2 U95 ( .A(N181), .B(n5), .Y(reg_read_data_2[3]) );
  MX2X1 U96 ( .A(n184), .B(n183), .S0(n215), .Y(N181) );
  MX4X1 U97 ( .A(\reg_array[0][3] ), .B(\reg_array[1][3] ), .C(
        \reg_array[2][3] ), .D(\reg_array[3][3] ), .S0(n212), .S1(n210), .Y(
        n184) );
  MX4X1 U98 ( .A(\reg_array[4][3] ), .B(\reg_array[5][3] ), .C(
        \reg_array[6][3] ), .D(\reg_array[7][3] ), .S0(n212), .S1(n210), .Y(
        n183) );
  INVX1 U99 ( .A(N18), .Y(n244) );
  AND2X1 U100 ( .A(N161), .B(n6), .Y(reg_read_data_1[7]) );
  MX2X1 U101 ( .A(n22), .B(n21), .S0(n176), .Y(N161) );
  MX4X1 U102 ( .A(\reg_array[0][7] ), .B(\reg_array[1][7] ), .C(
        \reg_array[2][7] ), .D(\reg_array[3][7] ), .S0(n175), .S1(n173), .Y(
        n22) );
  MX4X1 U103 ( .A(\reg_array[4][7] ), .B(\reg_array[5][7] ), .C(
        \reg_array[6][7] ), .D(\reg_array[7][7] ), .S0(n175), .S1(n173), .Y(
        n21) );
  AND2X1 U104 ( .A(N158), .B(n6), .Y(reg_read_data_1[10]) );
  MX2X1 U105 ( .A(n160), .B(n31), .S0(n176), .Y(N158) );
  MX4X1 U106 ( .A(\reg_array[0][10] ), .B(\reg_array[1][10] ), .C(
        \reg_array[2][10] ), .D(\reg_array[3][10] ), .S0(n175), .S1(n173), .Y(
        n160) );
  MX4X1 U107 ( .A(\reg_array[4][10] ), .B(\reg_array[5][10] ), .C(
        \reg_array[6][10] ), .D(\reg_array[7][10] ), .S0(n174), .S1(n172), .Y(
        n31) );
  AND2X1 U108 ( .A(N163), .B(n6), .Y(reg_read_data_1[5]) );
  MX2X1 U109 ( .A(n18), .B(n17), .S0(n176), .Y(N163) );
  MX4X1 U110 ( .A(\reg_array[0][5] ), .B(\reg_array[1][5] ), .C(
        \reg_array[2][5] ), .D(\reg_array[3][5] ), .S0(n175), .S1(n173), .Y(
        n18) );
  MX4X1 U111 ( .A(\reg_array[4][5] ), .B(\reg_array[5][5] ), .C(
        \reg_array[6][5] ), .D(\reg_array[7][5] ), .S0(n175), .S1(n173), .Y(
        n17) );
  BUFX3 U112 ( .A(N20), .Y(n176) );
  AND2X2 U113 ( .A(N179), .B(n5), .Y(reg_read_data_2[5]) );
  MX2X1 U114 ( .A(n188), .B(n187), .S0(n215), .Y(N179) );
  MX4X1 U115 ( .A(\reg_array[0][5] ), .B(\reg_array[1][5] ), .C(
        \reg_array[2][5] ), .D(\reg_array[3][5] ), .S0(n213), .S1(n211), .Y(
        n188) );
  MX4X1 U116 ( .A(\reg_array[4][5] ), .B(\reg_array[5][5] ), .C(
        \reg_array[6][5] ), .D(\reg_array[7][5] ), .S0(n213), .S1(n211), .Y(
        n187) );
  AND2X2 U117 ( .A(N178), .B(n5), .Y(reg_read_data_2[6]) );
  MX2X1 U118 ( .A(n190), .B(n189), .S0(n215), .Y(N178) );
  MX4X1 U119 ( .A(\reg_array[0][6] ), .B(\reg_array[1][6] ), .C(
        \reg_array[2][6] ), .D(\reg_array[3][6] ), .S0(n213), .S1(n211), .Y(
        n190) );
  MX4X1 U120 ( .A(\reg_array[4][6] ), .B(\reg_array[5][6] ), .C(
        \reg_array[6][6] ), .D(\reg_array[7][6] ), .S0(n213), .S1(n211), .Y(
        n189) );
  AND2X2 U121 ( .A(N177), .B(n5), .Y(reg_read_data_2[7]) );
  MX2X1 U122 ( .A(n192), .B(n191), .S0(n215), .Y(N177) );
  MX4X1 U123 ( .A(\reg_array[0][7] ), .B(\reg_array[1][7] ), .C(
        \reg_array[2][7] ), .D(\reg_array[3][7] ), .S0(n213), .S1(n211), .Y(
        n192) );
  MX4X1 U124 ( .A(\reg_array[4][7] ), .B(\reg_array[5][7] ), .C(
        \reg_array[6][7] ), .D(\reg_array[7][7] ), .S0(n213), .S1(n211), .Y(
        n191) );
  AND2X2 U125 ( .A(N176), .B(n5), .Y(reg_read_data_2[8]) );
  MX2X1 U126 ( .A(n194), .B(n193), .S0(n215), .Y(N176) );
  MX4X1 U127 ( .A(\reg_array[0][8] ), .B(\reg_array[1][8] ), .C(
        \reg_array[2][8] ), .D(\reg_array[3][8] ), .S0(n213), .S1(n211), .Y(
        n194) );
  MX4X1 U128 ( .A(\reg_array[4][8] ), .B(\reg_array[5][8] ), .C(
        \reg_array[6][8] ), .D(\reg_array[7][8] ), .S0(n213), .S1(n211), .Y(
        n193) );
  AND2X2 U129 ( .A(N175), .B(n5), .Y(reg_read_data_2[9]) );
  MX2X1 U130 ( .A(n196), .B(n195), .S0(n215), .Y(N175) );
  MX4X1 U131 ( .A(\reg_array[0][9] ), .B(\reg_array[1][9] ), .C(
        \reg_array[2][9] ), .D(\reg_array[3][9] ), .S0(n213), .S1(n211), .Y(
        n196) );
  MX4X1 U132 ( .A(\reg_array[4][9] ), .B(\reg_array[5][9] ), .C(
        \reg_array[6][9] ), .D(\reg_array[7][9] ), .S0(n213), .S1(n211), .Y(
        n195) );
  MX2X1 U133 ( .A(n10), .B(n9), .S0(n176), .Y(N167) );
  MX4X1 U134 ( .A(\reg_array[4][1] ), .B(\reg_array[5][1] ), .C(
        \reg_array[6][1] ), .D(\reg_array[7][1] ), .S0(n174), .S1(n172), .Y(n9) );
  MX4X1 U135 ( .A(\reg_array[0][1] ), .B(\reg_array[1][1] ), .C(
        \reg_array[2][1] ), .D(\reg_array[3][1] ), .S0(n174), .S1(n172), .Y(
        n10) );
  MX2X1 U136 ( .A(n12), .B(n11), .S0(n176), .Y(N166) );
  MX4X1 U137 ( .A(\reg_array[4][2] ), .B(\reg_array[5][2] ), .C(
        \reg_array[6][2] ), .D(\reg_array[7][2] ), .S0(n174), .S1(n172), .Y(
        n11) );
  MX4X1 U138 ( .A(\reg_array[0][2] ), .B(\reg_array[1][2] ), .C(
        \reg_array[2][2] ), .D(\reg_array[3][2] ), .S0(n174), .S1(n172), .Y(
        n12) );
  MX2X1 U139 ( .A(n14), .B(n13), .S0(n176), .Y(N165) );
  MX4X1 U140 ( .A(\reg_array[0][3] ), .B(\reg_array[1][3] ), .C(
        \reg_array[2][3] ), .D(\reg_array[3][3] ), .S0(n174), .S1(n172), .Y(
        n14) );
  MX4X1 U141 ( .A(\reg_array[4][3] ), .B(\reg_array[5][3] ), .C(
        \reg_array[6][3] ), .D(\reg_array[7][3] ), .S0(n174), .S1(n172), .Y(
        n13) );
  MX2X1 U142 ( .A(n16), .B(n15), .S0(n176), .Y(N164) );
  MX4X1 U143 ( .A(\reg_array[0][4] ), .B(\reg_array[1][4] ), .C(
        \reg_array[2][4] ), .D(\reg_array[3][4] ), .S0(n175), .S1(n173), .Y(
        n16) );
  MX4X1 U144 ( .A(\reg_array[4][4] ), .B(\reg_array[5][4] ), .C(
        \reg_array[6][4] ), .D(\reg_array[7][4] ), .S0(n175), .S1(n173), .Y(
        n15) );
  MX2X1 U145 ( .A(n20), .B(n19), .S0(n176), .Y(N162) );
  MX4X1 U146 ( .A(\reg_array[0][6] ), .B(\reg_array[1][6] ), .C(
        \reg_array[2][6] ), .D(\reg_array[3][6] ), .S0(n175), .S1(n173), .Y(
        n20) );
  MX4X1 U147 ( .A(\reg_array[4][6] ), .B(\reg_array[5][6] ), .C(
        \reg_array[6][6] ), .D(\reg_array[7][6] ), .S0(n175), .S1(n173), .Y(
        n19) );
  AND2X2 U148 ( .A(N157), .B(n6), .Y(reg_read_data_1[11]) );
  MX2X1 U149 ( .A(n162), .B(n161), .S0(n176), .Y(N157) );
  MX4X1 U150 ( .A(\reg_array[0][11] ), .B(\reg_array[1][11] ), .C(
        \reg_array[2][11] ), .D(\reg_array[3][11] ), .S0(N18), .S1(n172), .Y(
        n162) );
  MX4X1 U151 ( .A(\reg_array[4][11] ), .B(\reg_array[5][11] ), .C(
        \reg_array[6][11] ), .D(\reg_array[7][11] ), .S0(N18), .S1(n173), .Y(
        n161) );
  MX2X1 U152 ( .A(n170), .B(n169), .S0(n176), .Y(N153) );
  MX4X1 U153 ( .A(\reg_array[4][15] ), .B(\reg_array[5][15] ), .C(
        \reg_array[6][15] ), .D(\reg_array[7][15] ), .S0(N18), .S1(N19), .Y(
        n169) );
  MX4X1 U154 ( .A(\reg_array[0][15] ), .B(\reg_array[1][15] ), .C(
        \reg_array[2][15] ), .D(\reg_array[3][15] ), .S0(n175), .S1(n173), .Y(
        n170) );
  AND2X2 U155 ( .A(N174), .B(n5), .Y(reg_read_data_2[10]) );
  MX2X1 U156 ( .A(n198), .B(n197), .S0(n215), .Y(N174) );
  MX4X1 U157 ( .A(\reg_array[0][10] ), .B(\reg_array[1][10] ), .C(
        \reg_array[2][10] ), .D(\reg_array[3][10] ), .S0(n212), .S1(n210), .Y(
        n198) );
  MX4X1 U158 ( .A(\reg_array[4][10] ), .B(\reg_array[5][10] ), .C(
        \reg_array[6][10] ), .D(\reg_array[7][10] ), .S0(n212), .S1(n210), .Y(
        n197) );
  AND2X2 U159 ( .A(N173), .B(n5), .Y(reg_read_data_2[11]) );
  MX2X1 U160 ( .A(n200), .B(n199), .S0(n215), .Y(N173) );
  MX4X1 U161 ( .A(\reg_array[0][11] ), .B(\reg_array[1][11] ), .C(
        \reg_array[2][11] ), .D(\reg_array[3][11] ), .S0(n213), .S1(n210), .Y(
        n200) );
  MX4X1 U162 ( .A(\reg_array[4][11] ), .B(\reg_array[5][11] ), .C(
        \reg_array[6][11] ), .D(\reg_array[7][11] ), .S0(n212), .S1(n211), .Y(
        n199) );
  AND2X2 U163 ( .A(N172), .B(n5), .Y(reg_read_data_2[12]) );
  MX2X1 U164 ( .A(n202), .B(n201), .S0(n215), .Y(N172) );
  MX4X1 U165 ( .A(\reg_array[0][12] ), .B(\reg_array[1][12] ), .C(
        \reg_array[2][12] ), .D(\reg_array[3][12] ), .S0(n212), .S1(n210), .Y(
        n202) );
  MX4X1 U166 ( .A(\reg_array[4][12] ), .B(\reg_array[5][12] ), .C(
        \reg_array[6][12] ), .D(\reg_array[7][12] ), .S0(n212), .S1(n210), .Y(
        n201) );
  AND2X2 U167 ( .A(N171), .B(n5), .Y(reg_read_data_2[13]) );
  MX2X1 U168 ( .A(n204), .B(n203), .S0(n215), .Y(N171) );
  MX4X1 U169 ( .A(\reg_array[0][13] ), .B(\reg_array[1][13] ), .C(
        \reg_array[2][13] ), .D(\reg_array[3][13] ), .S0(n213), .S1(n210), .Y(
        n204) );
  MX4X1 U170 ( .A(\reg_array[4][13] ), .B(\reg_array[5][13] ), .C(
        \reg_array[6][13] ), .D(\reg_array[7][13] ), .S0(n212), .S1(n211), .Y(
        n203) );
  AND2X2 U171 ( .A(N170), .B(n5), .Y(reg_read_data_2[14]) );
  MX2X1 U172 ( .A(n206), .B(n205), .S0(n215), .Y(N170) );
  MX4X1 U173 ( .A(\reg_array[0][14] ), .B(\reg_array[1][14] ), .C(
        \reg_array[2][14] ), .D(\reg_array[3][14] ), .S0(n213), .S1(n210), .Y(
        n206) );
  MX4X1 U174 ( .A(\reg_array[4][14] ), .B(\reg_array[5][14] ), .C(
        \reg_array[6][14] ), .D(\reg_array[7][14] ), .S0(n212), .S1(N22), .Y(
        n205) );
  AND2X2 U175 ( .A(N169), .B(n5), .Y(reg_read_data_2[15]) );
  MX2X1 U176 ( .A(n208), .B(n207), .S0(n215), .Y(N169) );
  MX4X1 U177 ( .A(\reg_array[0][15] ), .B(\reg_array[1][15] ), .C(
        \reg_array[2][15] ), .D(\reg_array[3][15] ), .S0(N21), .S1(N22), .Y(
        n208) );
  MX4X1 U178 ( .A(\reg_array[4][15] ), .B(\reg_array[5][15] ), .C(
        \reg_array[6][15] ), .D(\reg_array[7][15] ), .S0(N21), .S1(N22), .Y(
        n207) );
  CLKINVX3 U179 ( .A(reg_write_data[0]), .Y(n260) );
  CLKINVX3 U180 ( .A(reg_write_data[1]), .Y(n259) );
  CLKINVX3 U181 ( .A(reg_write_data[2]), .Y(n258) );
  CLKINVX3 U182 ( .A(reg_write_data[3]), .Y(n257) );
  CLKINVX3 U183 ( .A(reg_write_data[4]), .Y(n256) );
  INVX1 U184 ( .A(reg_write_dest[2]), .Y(n261) );
  INVX1 U185 ( .A(reg_write_dest[1]), .Y(n262) );
  INVX1 U186 ( .A(reg_write_dest[0]), .Y(n263) );
  NAND4X1 U187 ( .A(reg_write_en), .B(n263), .C(n262), .D(n261), .Y(n24) );
  NAND4X1 U188 ( .A(reg_write_dest[2]), .B(reg_write_en), .C(n263), .D(n262), 
        .Y(n28) );
  NAND4X1 U189 ( .A(reg_write_dest[2]), .B(reg_write_dest[0]), .C(reg_write_en), .D(n262), .Y(n29) );
  CLKINVX3 U190 ( .A(reg_write_data[5]), .Y(n255) );
  CLKINVX3 U191 ( .A(reg_write_data[6]), .Y(n254) );
  CLKINVX3 U192 ( .A(reg_write_data[7]), .Y(n253) );
  CLKINVX3 U193 ( .A(reg_write_data[8]), .Y(n252) );
  CLKINVX3 U194 ( .A(reg_write_data[9]), .Y(n251) );
  CLKINVX3 U195 ( .A(reg_write_data[10]), .Y(n250) );
  CLKINVX3 U196 ( .A(reg_write_data[11]), .Y(n249) );
  CLKINVX3 U197 ( .A(reg_write_data[12]), .Y(n248) );
  CLKINVX3 U198 ( .A(reg_write_data[13]), .Y(n247) );
  CLKINVX3 U199 ( .A(reg_write_data[14]), .Y(n246) );
  CLKINVX3 U200 ( .A(reg_write_data[15]), .Y(n245) );
  OAI2BB2X1 U201 ( .B0(n241), .B1(n260), .A0N(\reg_array[0][0] ), .A1N(n242), 
        .Y(n32) );
  OAI2BB2X1 U202 ( .B0(n241), .B1(n259), .A0N(\reg_array[0][1] ), .A1N(n242), 
        .Y(n33) );
  OAI2BB2X1 U203 ( .B0(n241), .B1(n258), .A0N(\reg_array[0][2] ), .A1N(n242), 
        .Y(n34) );
  OAI2BB2X1 U204 ( .B0(n241), .B1(n257), .A0N(\reg_array[0][3] ), .A1N(n242), 
        .Y(n35) );
  OAI2BB2X1 U205 ( .B0(n241), .B1(n256), .A0N(\reg_array[0][4] ), .A1N(n241), 
        .Y(n36) );
  OAI2BB2X1 U206 ( .B0(n24), .B1(n255), .A0N(\reg_array[0][5] ), .A1N(n241), 
        .Y(n37) );
  OAI2BB2X1 U207 ( .B0(n24), .B1(n254), .A0N(\reg_array[0][6] ), .A1N(n241), 
        .Y(n38) );
  OAI2BB2X1 U208 ( .B0(n24), .B1(n253), .A0N(\reg_array[0][7] ), .A1N(n241), 
        .Y(n39) );
  OAI2BB2X1 U209 ( .B0(n24), .B1(n252), .A0N(\reg_array[0][8] ), .A1N(n241), 
        .Y(n40) );
  OAI2BB2X1 U210 ( .B0(n24), .B1(n251), .A0N(\reg_array[0][9] ), .A1N(n241), 
        .Y(n41) );
  OAI2BB2X1 U211 ( .B0(n241), .B1(n250), .A0N(\reg_array[0][10] ), .A1N(n241), 
        .Y(n42) );
  OAI2BB2X1 U212 ( .B0(n242), .B1(n249), .A0N(\reg_array[0][11] ), .A1N(n241), 
        .Y(n43) );
  OAI2BB2X1 U213 ( .B0(n241), .B1(n248), .A0N(\reg_array[0][12] ), .A1N(n241), 
        .Y(n44) );
  OAI2BB2X1 U214 ( .B0(n241), .B1(n247), .A0N(\reg_array[0][13] ), .A1N(n241), 
        .Y(n45) );
  OAI2BB2X1 U215 ( .B0(n241), .B1(n246), .A0N(\reg_array[0][14] ), .A1N(n242), 
        .Y(n46) );
  OAI2BB2X1 U216 ( .B0(n241), .B1(n245), .A0N(\reg_array[0][15] ), .A1N(n242), 
        .Y(n47) );
  OAI2BB2X1 U217 ( .B0(n260), .B1(n239), .A0N(\reg_array[1][0] ), .A1N(n240), 
        .Y(n48) );
  OAI2BB2X1 U218 ( .B0(n259), .B1(n239), .A0N(\reg_array[1][1] ), .A1N(n239), 
        .Y(n49) );
  OAI2BB2X1 U219 ( .B0(n258), .B1(n239), .A0N(\reg_array[1][2] ), .A1N(n240), 
        .Y(n50) );
  OAI2BB2X1 U220 ( .B0(n257), .B1(n239), .A0N(\reg_array[1][3] ), .A1N(n239), 
        .Y(n51) );
  OAI2BB2X1 U221 ( .B0(n256), .B1(n239), .A0N(\reg_array[1][4] ), .A1N(n240), 
        .Y(n52) );
  OAI2BB2X1 U222 ( .B0(n255), .B1(n239), .A0N(\reg_array[1][5] ), .A1N(n240), 
        .Y(n53) );
  OAI2BB2X1 U223 ( .B0(n254), .B1(n239), .A0N(\reg_array[1][6] ), .A1N(n240), 
        .Y(n54) );
  OAI2BB2X1 U224 ( .B0(n253), .B1(n239), .A0N(\reg_array[1][7] ), .A1N(n240), 
        .Y(n55) );
  OAI2BB2X1 U225 ( .B0(n252), .B1(n239), .A0N(\reg_array[1][8] ), .A1N(n240), 
        .Y(n56) );
  OAI2BB2X1 U226 ( .B0(n251), .B1(n239), .A0N(\reg_array[1][9] ), .A1N(n240), 
        .Y(n57) );
  OAI2BB2X1 U227 ( .B0(n250), .B1(n239), .A0N(\reg_array[1][10] ), .A1N(n240), 
        .Y(n58) );
  OAI2BB2X1 U228 ( .B0(n249), .B1(n239), .A0N(\reg_array[1][11] ), .A1N(n240), 
        .Y(n59) );
  OAI2BB2X1 U229 ( .B0(n248), .B1(n240), .A0N(\reg_array[1][12] ), .A1N(n240), 
        .Y(n60) );
  OAI2BB2X1 U230 ( .B0(n247), .B1(n240), .A0N(\reg_array[1][13] ), .A1N(n240), 
        .Y(n61) );
  OAI2BB2X1 U231 ( .B0(n246), .B1(n240), .A0N(\reg_array[1][14] ), .A1N(n239), 
        .Y(n62) );
  OAI2BB2X1 U232 ( .B0(n245), .B1(n240), .A0N(\reg_array[1][15] ), .A1N(n239), 
        .Y(n63) );
  OAI2BB2X1 U233 ( .B0(n260), .B1(n237), .A0N(\reg_array[2][0] ), .A1N(n238), 
        .Y(n64) );
  OAI2BB2X1 U234 ( .B0(n259), .B1(n237), .A0N(\reg_array[2][1] ), .A1N(n237), 
        .Y(n65) );
  OAI2BB2X1 U235 ( .B0(n258), .B1(n237), .A0N(\reg_array[2][2] ), .A1N(n238), 
        .Y(n66) );
  OAI2BB2X1 U236 ( .B0(n257), .B1(n237), .A0N(\reg_array[2][3] ), .A1N(n237), 
        .Y(n67) );
  OAI2BB2X1 U237 ( .B0(n256), .B1(n237), .A0N(\reg_array[2][4] ), .A1N(n238), 
        .Y(n68) );
  OAI2BB2X1 U238 ( .B0(n255), .B1(n237), .A0N(\reg_array[2][5] ), .A1N(n238), 
        .Y(n69) );
  OAI2BB2X1 U239 ( .B0(n254), .B1(n237), .A0N(\reg_array[2][6] ), .A1N(n238), 
        .Y(n70) );
  OAI2BB2X1 U240 ( .B0(n253), .B1(n237), .A0N(\reg_array[2][7] ), .A1N(n238), 
        .Y(n71) );
  OAI2BB2X1 U241 ( .B0(n252), .B1(n237), .A0N(\reg_array[2][8] ), .A1N(n238), 
        .Y(n72) );
  OAI2BB2X1 U242 ( .B0(n251), .B1(n237), .A0N(\reg_array[2][9] ), .A1N(n238), 
        .Y(n73) );
  OAI2BB2X1 U243 ( .B0(n250), .B1(n237), .A0N(\reg_array[2][10] ), .A1N(n238), 
        .Y(n74) );
  OAI2BB2X1 U244 ( .B0(n249), .B1(n237), .A0N(\reg_array[2][11] ), .A1N(n238), 
        .Y(n75) );
  OAI2BB2X1 U245 ( .B0(n248), .B1(n238), .A0N(\reg_array[2][12] ), .A1N(n238), 
        .Y(n76) );
  OAI2BB2X1 U246 ( .B0(n247), .B1(n238), .A0N(\reg_array[2][13] ), .A1N(n238), 
        .Y(n77) );
  OAI2BB2X1 U247 ( .B0(n246), .B1(n238), .A0N(\reg_array[2][14] ), .A1N(n237), 
        .Y(n78) );
  OAI2BB2X1 U248 ( .B0(n245), .B1(n238), .A0N(\reg_array[2][15] ), .A1N(n237), 
        .Y(n79) );
  OAI2BB2X1 U249 ( .B0(n260), .B1(n234), .A0N(\reg_array[3][0] ), .A1N(n235), 
        .Y(n80) );
  OAI2BB2X1 U250 ( .B0(n259), .B1(n234), .A0N(\reg_array[3][1] ), .A1N(n235), 
        .Y(n81) );
  OAI2BB2X1 U251 ( .B0(n258), .B1(n234), .A0N(\reg_array[3][2] ), .A1N(n235), 
        .Y(n82) );
  OAI2BB2X1 U252 ( .B0(n257), .B1(n234), .A0N(\reg_array[3][3] ), .A1N(n235), 
        .Y(n83) );
  OAI2BB2X1 U253 ( .B0(n256), .B1(n234), .A0N(\reg_array[3][4] ), .A1N(n234), 
        .Y(n84) );
  OAI2BB2X1 U254 ( .B0(n255), .B1(n234), .A0N(\reg_array[3][5] ), .A1N(n234), 
        .Y(n85) );
  OAI2BB2X1 U255 ( .B0(n254), .B1(n27), .A0N(\reg_array[3][6] ), .A1N(n234), 
        .Y(n86) );
  OAI2BB2X1 U256 ( .B0(n253), .B1(n27), .A0N(\reg_array[3][7] ), .A1N(n234), 
        .Y(n87) );
  OAI2BB2X1 U257 ( .B0(n252), .B1(n235), .A0N(\reg_array[3][8] ), .A1N(n234), 
        .Y(n88) );
  OAI2BB2X1 U258 ( .B0(n251), .B1(n234), .A0N(\reg_array[3][9] ), .A1N(n234), 
        .Y(n89) );
  OAI2BB2X1 U259 ( .B0(n250), .B1(n27), .A0N(\reg_array[3][10] ), .A1N(n234), 
        .Y(n90) );
  OAI2BB2X1 U260 ( .B0(n249), .B1(n27), .A0N(\reg_array[3][11] ), .A1N(n234), 
        .Y(n91) );
  OAI2BB2X1 U261 ( .B0(n248), .B1(n234), .A0N(\reg_array[3][12] ), .A1N(n234), 
        .Y(n92) );
  OAI2BB2X1 U262 ( .B0(n247), .B1(n234), .A0N(\reg_array[3][13] ), .A1N(n234), 
        .Y(n93) );
  OAI2BB2X1 U263 ( .B0(n246), .B1(n234), .A0N(\reg_array[3][14] ), .A1N(n235), 
        .Y(n94) );
  OAI2BB2X1 U264 ( .B0(n245), .B1(n234), .A0N(\reg_array[3][15] ), .A1N(n235), 
        .Y(n95) );
  OAI2BB2X1 U265 ( .B0(n260), .B1(n231), .A0N(\reg_array[4][0] ), .A1N(n232), 
        .Y(n96) );
  OAI2BB2X1 U266 ( .B0(n259), .B1(n231), .A0N(\reg_array[4][1] ), .A1N(n232), 
        .Y(n97) );
  OAI2BB2X1 U267 ( .B0(n258), .B1(n231), .A0N(\reg_array[4][2] ), .A1N(n232), 
        .Y(n98) );
  OAI2BB2X1 U268 ( .B0(n257), .B1(n231), .A0N(\reg_array[4][3] ), .A1N(n232), 
        .Y(n99) );
  OAI2BB2X1 U269 ( .B0(n256), .B1(n28), .A0N(\reg_array[4][4] ), .A1N(n231), 
        .Y(n100) );
  OAI2BB2X1 U270 ( .B0(n255), .B1(n28), .A0N(\reg_array[4][5] ), .A1N(n231), 
        .Y(n101) );
  OAI2BB2X1 U271 ( .B0(n254), .B1(n28), .A0N(\reg_array[4][6] ), .A1N(n231), 
        .Y(n102) );
  OAI2BB2X1 U272 ( .B0(n253), .B1(n28), .A0N(\reg_array[4][7] ), .A1N(n231), 
        .Y(n103) );
  OAI2BB2X1 U273 ( .B0(n252), .B1(n28), .A0N(\reg_array[4][8] ), .A1N(n231), 
        .Y(n104) );
  OAI2BB2X1 U274 ( .B0(n251), .B1(n28), .A0N(\reg_array[4][9] ), .A1N(n231), 
        .Y(n105) );
  OAI2BB2X1 U275 ( .B0(n250), .B1(n231), .A0N(\reg_array[4][10] ), .A1N(n231), 
        .Y(n106) );
  OAI2BB2X1 U276 ( .B0(n249), .B1(n231), .A0N(\reg_array[4][11] ), .A1N(n231), 
        .Y(n107) );
  OAI2BB2X1 U277 ( .B0(n248), .B1(n231), .A0N(\reg_array[4][12] ), .A1N(n231), 
        .Y(n108) );
  OAI2BB2X1 U278 ( .B0(n247), .B1(n231), .A0N(\reg_array[4][13] ), .A1N(n231), 
        .Y(n109) );
  OAI2BB2X1 U279 ( .B0(n246), .B1(n231), .A0N(\reg_array[4][14] ), .A1N(n232), 
        .Y(n110) );
  OAI2BB2X1 U280 ( .B0(n245), .B1(n231), .A0N(\reg_array[4][15] ), .A1N(n232), 
        .Y(n111) );
  OAI2BB2X1 U281 ( .B0(n260), .B1(n228), .A0N(\reg_array[5][0] ), .A1N(n229), 
        .Y(n112) );
  OAI2BB2X1 U282 ( .B0(n259), .B1(n228), .A0N(\reg_array[5][1] ), .A1N(n229), 
        .Y(n113) );
  OAI2BB2X1 U283 ( .B0(n258), .B1(n228), .A0N(\reg_array[5][2] ), .A1N(n229), 
        .Y(n114) );
  OAI2BB2X1 U284 ( .B0(n257), .B1(n228), .A0N(\reg_array[5][3] ), .A1N(n229), 
        .Y(n115) );
  OAI2BB2X1 U285 ( .B0(n256), .B1(n29), .A0N(\reg_array[5][4] ), .A1N(n228), 
        .Y(n116) );
  OAI2BB2X1 U286 ( .B0(n255), .B1(n29), .A0N(\reg_array[5][5] ), .A1N(n228), 
        .Y(n117) );
  OAI2BB2X1 U287 ( .B0(n254), .B1(n29), .A0N(\reg_array[5][6] ), .A1N(n228), 
        .Y(n118) );
  OAI2BB2X1 U288 ( .B0(n253), .B1(n29), .A0N(\reg_array[5][7] ), .A1N(n228), 
        .Y(n119) );
  OAI2BB2X1 U289 ( .B0(n252), .B1(n29), .A0N(\reg_array[5][8] ), .A1N(n228), 
        .Y(n120) );
  OAI2BB2X1 U290 ( .B0(n251), .B1(n29), .A0N(\reg_array[5][9] ), .A1N(n228), 
        .Y(n121) );
  OAI2BB2X1 U291 ( .B0(n250), .B1(n228), .A0N(\reg_array[5][10] ), .A1N(n228), 
        .Y(n122) );
  OAI2BB2X1 U292 ( .B0(n249), .B1(n228), .A0N(\reg_array[5][11] ), .A1N(n228), 
        .Y(n123) );
  OAI2BB2X1 U293 ( .B0(n248), .B1(n228), .A0N(\reg_array[5][12] ), .A1N(n228), 
        .Y(n124) );
  OAI2BB2X1 U294 ( .B0(n247), .B1(n228), .A0N(\reg_array[5][13] ), .A1N(n228), 
        .Y(n125) );
  OAI2BB2X1 U295 ( .B0(n246), .B1(n228), .A0N(\reg_array[5][14] ), .A1N(n229), 
        .Y(n126) );
  OAI2BB2X1 U296 ( .B0(n245), .B1(n228), .A0N(\reg_array[5][15] ), .A1N(n229), 
        .Y(n127) );
  OAI2BB2X1 U297 ( .B0(n260), .B1(n226), .A0N(\reg_array[6][0] ), .A1N(n227), 
        .Y(n128) );
  OAI2BB2X1 U298 ( .B0(n259), .B1(n226), .A0N(\reg_array[6][1] ), .A1N(n226), 
        .Y(n129) );
  OAI2BB2X1 U299 ( .B0(n258), .B1(n226), .A0N(\reg_array[6][2] ), .A1N(n227), 
        .Y(n130) );
  OAI2BB2X1 U300 ( .B0(n257), .B1(n226), .A0N(\reg_array[6][3] ), .A1N(n226), 
        .Y(n131) );
  OAI2BB2X1 U301 ( .B0(n256), .B1(n226), .A0N(\reg_array[6][4] ), .A1N(n227), 
        .Y(n132) );
  OAI2BB2X1 U302 ( .B0(n255), .B1(n226), .A0N(\reg_array[6][5] ), .A1N(n227), 
        .Y(n133) );
  OAI2BB2X1 U303 ( .B0(n254), .B1(n226), .A0N(\reg_array[6][6] ), .A1N(n227), 
        .Y(n134) );
  OAI2BB2X1 U304 ( .B0(n253), .B1(n226), .A0N(\reg_array[6][7] ), .A1N(n227), 
        .Y(n135) );
  OAI2BB2X1 U305 ( .B0(n252), .B1(n226), .A0N(\reg_array[6][8] ), .A1N(n227), 
        .Y(n136) );
  OAI2BB2X1 U306 ( .B0(n251), .B1(n226), .A0N(\reg_array[6][9] ), .A1N(n227), 
        .Y(n137) );
  OAI2BB2X1 U307 ( .B0(n250), .B1(n226), .A0N(\reg_array[6][10] ), .A1N(n227), 
        .Y(n138) );
  OAI2BB2X1 U308 ( .B0(n249), .B1(n226), .A0N(\reg_array[6][11] ), .A1N(n227), 
        .Y(n139) );
  OAI2BB2X1 U309 ( .B0(n248), .B1(n227), .A0N(\reg_array[6][12] ), .A1N(n227), 
        .Y(n140) );
  OAI2BB2X1 U310 ( .B0(n247), .B1(n227), .A0N(\reg_array[6][13] ), .A1N(n227), 
        .Y(n141) );
  OAI2BB2X1 U311 ( .B0(n246), .B1(n227), .A0N(\reg_array[6][14] ), .A1N(n226), 
        .Y(n142) );
  OAI2BB2X1 U312 ( .B0(n245), .B1(n227), .A0N(\reg_array[6][15] ), .A1N(n226), 
        .Y(n143) );
  OAI2BB2X1 U313 ( .B0(n260), .B1(n224), .A0N(\reg_array[7][0] ), .A1N(n224), 
        .Y(n144) );
  OAI2BB2X1 U314 ( .B0(n259), .B1(n224), .A0N(\reg_array[7][1] ), .A1N(n225), 
        .Y(n145) );
  OAI2BB2X1 U315 ( .B0(n258), .B1(n224), .A0N(\reg_array[7][2] ), .A1N(n224), 
        .Y(n146) );
  OAI2BB2X1 U316 ( .B0(n257), .B1(n224), .A0N(\reg_array[7][3] ), .A1N(n225), 
        .Y(n147) );
  OAI2BB2X1 U317 ( .B0(n256), .B1(n224), .A0N(\reg_array[7][4] ), .A1N(n225), 
        .Y(n148) );
  OAI2BB2X1 U318 ( .B0(n255), .B1(n224), .A0N(\reg_array[7][5] ), .A1N(n225), 
        .Y(n149) );
  OAI2BB2X1 U319 ( .B0(n254), .B1(n224), .A0N(\reg_array[7][6] ), .A1N(n225), 
        .Y(n150) );
  OAI2BB2X1 U320 ( .B0(n253), .B1(n224), .A0N(\reg_array[7][7] ), .A1N(n225), 
        .Y(n151) );
  OAI2BB2X1 U321 ( .B0(n252), .B1(n224), .A0N(\reg_array[7][8] ), .A1N(n225), 
        .Y(n152) );
  OAI2BB2X1 U322 ( .B0(n251), .B1(n224), .A0N(\reg_array[7][9] ), .A1N(n225), 
        .Y(n153) );
  OAI2BB2X1 U323 ( .B0(n250), .B1(n224), .A0N(\reg_array[7][10] ), .A1N(n225), 
        .Y(n154) );
  OAI2BB2X1 U324 ( .B0(n249), .B1(n224), .A0N(\reg_array[7][11] ), .A1N(n225), 
        .Y(n155) );
  OAI2BB2X1 U325 ( .B0(n248), .B1(n225), .A0N(\reg_array[7][12] ), .A1N(n225), 
        .Y(n156) );
  OAI2BB2X1 U326 ( .B0(n247), .B1(n225), .A0N(\reg_array[7][13] ), .A1N(n225), 
        .Y(n157) );
  OAI2BB2X1 U327 ( .B0(n246), .B1(n225), .A0N(\reg_array[7][14] ), .A1N(n224), 
        .Y(n158) );
  OAI2BB2X1 U328 ( .B0(n245), .B1(n225), .A0N(\reg_array[7][15] ), .A1N(n224), 
        .Y(n159) );
endmodule


module hazard_detection_unit ( decoding_op_src1, decoding_op_src2, ex_op_dest, 
        mem_op_dest, wb_op_dest, pipeline_stall_n );
  input [2:0] decoding_op_src1;
  input [2:0] decoding_op_src2;
  input [2:0] ex_op_dest;
  input [2:0] mem_op_dest;
  input [2:0] wb_op_dest;
  output pipeline_stall_n;
  wire   n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n1, n2, n3, n4, n5,
         n6, n7;

  INVX1 U2 ( .A(decoding_op_src2[1]), .Y(n5) );
  INVX1 U3 ( .A(decoding_op_src2[2]), .Y(n6) );
  INVX1 U4 ( .A(decoding_op_src2[0]), .Y(n4) );
  NOR2X1 U5 ( .A(n20), .B(n21), .Y(pipeline_stall_n) );
  AOI31X1 U6 ( .A0(n3), .A1(n7), .A2(n1), .B0(n33), .Y(n20) );
  AOI31X1 U7 ( .A0(n5), .A1(n6), .A2(n4), .B0(n22), .Y(n21) );
  AOI31X1 U8 ( .A0(n23), .A1(n24), .A2(n25), .B0(n26), .Y(n22) );
  XNOR2X1 U9 ( .A(ex_op_dest[1]), .B(decoding_op_src2[1]), .Y(n25) );
  XNOR2X1 U10 ( .A(ex_op_dest[0]), .B(decoding_op_src2[0]), .Y(n24) );
  XNOR2X1 U11 ( .A(wb_op_dest[1]), .B(n5), .Y(n30) );
  XNOR2X1 U12 ( .A(wb_op_dest[0]), .B(n4), .Y(n31) );
  XNOR2X1 U13 ( .A(wb_op_dest[2]), .B(n6), .Y(n32) );
  OAI33X1 U14 ( .A0(n27), .A1(n28), .A2(n29), .B0(n30), .B1(n31), .B2(n32), 
        .Y(n26) );
  XNOR2X1 U15 ( .A(mem_op_dest[1]), .B(n5), .Y(n27) );
  XNOR2X1 U16 ( .A(mem_op_dest[0]), .B(n4), .Y(n28) );
  XNOR2X1 U17 ( .A(mem_op_dest[2]), .B(n6), .Y(n29) );
  AOI31X1 U18 ( .A0(n34), .A1(n35), .A2(n36), .B0(n37), .Y(n33) );
  XNOR2X1 U19 ( .A(ex_op_dest[2]), .B(decoding_op_src1[2]), .Y(n34) );
  XNOR2X1 U20 ( .A(ex_op_dest[0]), .B(decoding_op_src1[0]), .Y(n35) );
  XNOR2X1 U21 ( .A(ex_op_dest[1]), .B(n2), .Y(n36) );
  XNOR2X1 U22 ( .A(ex_op_dest[2]), .B(decoding_op_src2[2]), .Y(n23) );
  XNOR2X1 U23 ( .A(wb_op_dest[1]), .B(n3), .Y(n41) );
  XNOR2X1 U24 ( .A(wb_op_dest[0]), .B(n1), .Y(n42) );
  OAI33X1 U25 ( .A0(n38), .A1(n39), .A2(n40), .B0(n41), .B1(n42), .B2(n43), 
        .Y(n37) );
  XNOR2X1 U26 ( .A(mem_op_dest[2]), .B(n7), .Y(n40) );
  XNOR2X1 U27 ( .A(wb_op_dest[2]), .B(n7), .Y(n43) );
  XNOR2X1 U28 ( .A(mem_op_dest[1]), .B(n3), .Y(n38) );
  XNOR2X1 U29 ( .A(mem_op_dest[0]), .B(n1), .Y(n39) );
  INVX1 U30 ( .A(n3), .Y(n2) );
  INVX1 U31 ( .A(decoding_op_src1[1]), .Y(n3) );
  INVX1 U32 ( .A(decoding_op_src1[0]), .Y(n1) );
  INVX1 U33 ( .A(decoding_op_src1[2]), .Y(n7) );
endmodule


module mips_16_core_top ( clk, rst, pc );
  output [7:0] pc;
  input clk, rst;
  wire   pipeline_stall_n, branch_taken, reg_write_en, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [5:0] branch_offset_imm;
  wire   [56:0] ID_pipeline_reg_out;
  wire   [2:0] reg_read_addr_1;
  wire   [2:0] reg_read_addr_2;
  wire   [15:0] reg_read_data_1;
  wire   [15:0] reg_read_data_2;
  wire   [2:0] decoding_op_src1;
  wire   [2:0] decoding_op_src2;
  wire   [37:0] EX_pipeline_reg_out;
  wire   [2:0] ex_op_dest;
  wire   [36:0] MEM_pipeline_reg_out;
  wire   [2:0] mem_op_dest;
  wire   [2:0] reg_write_dest;
  wire   [15:0] reg_write_data;
  wire   [2:0] wb_op_dest;
  wire   SYNOPSYS_UNCONNECTED__0;

  IF_stage IF_stage_inst ( .clk(clk), .rst(rst), .instruction_fetch_en(n12), 
        .branch_offset_imm(branch_offset_imm), .branch_taken(branch_taken), 
        .pc(pc) );
  ID_stage ID_stage_inst ( .clk(clk), .rst(rst), .instruction_decode_en(n12), 
        .pipeline_reg_out(ID_pipeline_reg_out), .instruction({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .branch_offset_imm(branch_offset_imm), .branch_taken(
        branch_taken), .reg_read_addr_1({reg_read_addr_1[2:1], 
        SYNOPSYS_UNCONNECTED__0}), .reg_read_addr_2(reg_read_addr_2), 
        .reg_read_data_1(reg_read_data_1), .reg_read_data_2(reg_read_data_2), 
        .decoding_op_src1(decoding_op_src1), .decoding_op_src2(
        decoding_op_src2) );
  EX_stage EX_stage_inst ( .clk(clk), .rst(rst), .pipeline_reg_in(
        ID_pipeline_reg_out), .pipeline_reg_out(EX_pipeline_reg_out), 
        .ex_op_dest(ex_op_dest) );
  MEM_stage MEM_stage_inst ( .clk(clk), .rst(rst), .pipeline_reg_in({
        EX_pipeline_reg_out[37:27], n8, EX_pipeline_reg_out[25], n6, 
        EX_pipeline_reg_out[23], n4, n2, EX_pipeline_reg_out[20:0]}), 
        .pipeline_reg_out(MEM_pipeline_reg_out), .mem_op_dest(mem_op_dest) );
  WB_stage WB_stage_inst ( .pipeline_reg_in(MEM_pipeline_reg_out), 
        .reg_write_en(reg_write_en), .reg_write_dest(reg_write_dest), 
        .reg_write_data(reg_write_data), .wb_op_dest(wb_op_dest) );
  register_file register_file_inst ( .clk(clk), .rst(rst), .reg_write_en(
        reg_write_en), .reg_write_dest(reg_write_dest), .reg_write_data(
        reg_write_data), .reg_read_addr_1({reg_read_addr_1[2:1], n10}), 
        .reg_read_data_1(reg_read_data_1), .reg_read_addr_2(reg_read_addr_2), 
        .reg_read_data_2(reg_read_data_2) );
  hazard_detection_unit hazard_detection_unit_inst ( .decoding_op_src1({
        decoding_op_src1[2:1], n10}), .decoding_op_src2(decoding_op_src2), 
        .ex_op_dest(ex_op_dest), .mem_op_dest(mem_op_dest), .wb_op_dest(
        wb_op_dest), .pipeline_stall_n(pipeline_stall_n) );
  INVX1 U1 ( .A(n13), .Y(n12) );
  INVX1 U2 ( .A(pipeline_stall_n), .Y(n13) );
  INVX1 U3 ( .A(n11), .Y(n10) );
  INVX1 U4 ( .A(decoding_op_src1[0]), .Y(n11) );
  INVX1 U5 ( .A(n5), .Y(n4) );
  INVX1 U6 ( .A(EX_pipeline_reg_out[22]), .Y(n5) );
  INVX1 U7 ( .A(n7), .Y(n6) );
  INVX1 U8 ( .A(EX_pipeline_reg_out[24]), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n8) );
  INVX1 U10 ( .A(EX_pipeline_reg_out[26]), .Y(n9) );
  INVX1 U11 ( .A(n3), .Y(n2) );
  INVX1 U12 ( .A(EX_pipeline_reg_out[21]), .Y(n3) );
endmodule

